`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2020.3"
`protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
KC09Q2uxRQFYMyPg9w0O/oUjuUJ/wfEpxLzgay5G0565nXgcBv/GCmO/9uuvGoRh8dASOeJ++hl1
GBzOXuSvPg==

`protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
MoN3Cu5MMf8A/D/Et/jS1pM62FH4GTOH30Bsum+lprhTHqgFzvwRm6gr6mY+izobO5blI9kGhJMO
Grdqnls3mZTMmqWycxTxDURQP/65d8KHbWeB1RgwRbsB3miEadtBDEMNTIjKEtnfZ8v1riAc4vlG
DoVoeTdtF3igVH4l/Uc=

`protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
REiFE6BGwfX/9Gy2SKwpRz1NTgODK5Yts5rCD69n0dA05mbCCYRiw76TurtT3kAKdIvzdcqPpqd8
wgyGUNpbTTbGhm9SytleuiORBfePI6xgVawHLFMf8g6g5NwDX9dYyKrOijD+liv2DnpVNfAPbDcg
Tovnf18xgGuroMIOh3wthqvzfzbN4bb/FIBPg9SehYYXSJwGO0frVebWlhyuTkzHyjiK0wPN/R2E
SErGyAlDb2cD6A0ZzLj0oVVW8VZad7h8ThDxOJXVhhwIIBoH3FXQRfzQaSMd5YR/Hut90ybIgFgf
TyHrDYMePv9K+VaDOyItm5MP6UN78adAZXRp4A==

`protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
fZTybnin8+K/iw4ct+7PwD44stx+HRvxwFbe39HRK2NIoYaVZiaMM1Ud0zJFXexLIIyFAuasVUx1
kWED9JDYoxTWt0Z/FvaSb+RIOSL+bMtg0TFVH8H90AY4sCxmUhZjykzvkyIkFXrLjvKhUyeR+CAw
TS134Gwk5op5tpAJtg6m7pvHfzr7ghmu+55LvyV+uD/42IZw7AzwtxveCJETQxamX6KxppePGGK7
smfzq4t50140dFkm37l4Wt4hjFvn08ib8ymlKlVj3Dy+6YpeYfj4CluHuerBwVQcBonMtJgnbG+k
04Po5NiqXyd74+iUWuP3KRBJzA0383L9Xv8XuA==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VELOCE-RSA", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
avyxM2bpCK2VST8XK5nnZwPEs00648rgcUf9caYtcUEasP+ZGsvazauK5FRLCmZ6VNbhtSaiIdjf
frWVZ0PkFUo8/u4/nnCy4behMKZXYobEEECWmMhKBeUh3287wUJLx8CsNPU0ElMyVk2pDcZpyEyl
4J5ULzRXHbLhN5xC7sQ=

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
rrqVXk74zV2OFXif/fSF5FhEqRUT6iPT3Plhh+Ez25qHP9NCgU+vYdawDHCOk52dTIsbIfLu1GxV
d0Oh6UHKAyIWsBzsZXhDhU8I5Sb6oJ34QZG+2E9xbSoANvowVtdJCdSJHSYW5CX2oX4SNtrGXW1+
XtCileVcxriZEyobLxpv7bNxUZ55/V9md63zztlUAxDDySA307otDPK8PhkLApHWyUvdrniJfwAu
9Tgl+K2kv8LmYES0yz9OpBDw/ju2wFi7QirTBCPNsltPnckEHBqB9kBG48yTrdWvXrzUUKnS8Gxc
YO7yLVWQUhh5ytfUl+ffpqPbfBayDuTRtk0rXg==

`protect key_keyowner = "Real Intent", key_keyname = "RI-RSA-KEY-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
evewr6wVU+ZUQdhDf2PdACzpJMMgwHMfd3Euk4XZDXDyLZKyweFOmdH8GCnP9+9q10ka5rAayi4b
lSTXUun6Z/8Gm8wdVIM1JoRv2PWXknoixvwBo0R9hhvfRkDUFJ4EOuatsS3PKhL8saa7a2B96Gfp
CwgL6MmSfDS2oxGu3xYnqQd1i1z72sk+JTSl77t50ZUupsg7c4Ff0R9IPZwGkM3K2SQinKz2zPxf
ORlS45obnAA1YseY/4B1T0c+SgEOTDY8OOUqXjZLLSoY17bDgD/8b5Pht72jf2GkL1XnX0lsYMmF
N+gfW+MvS2F3DoqJc/DXcwn63nlZbjlD3VWhug==

`protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2020_08", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
XFNsTf6fx2/lQ1mBnmw+PGjdutQeGcJ+mDglE2tNwySDOmT2JdsKRN1ypmspciHnol8nD7z7mu48
QAjdHWExFVd7i+KL63tSwXG3QROI1hqgz+M662N+5YUJ8ZXi/UILO3mEnOvMqf8i/dLebaw4CdUE
LpEVFTcCCL0dDkFXhkTsV33K6IMQX29BbnCavXk9j/p6o80cO4oHMCoOc/QiIqpvyOzRTVrB5cCF
fTtveWkIEEz5usrMTPzFkx5OJjn5s/JIRcux2Ya4C8AtM3a61FeMbHv5TxtXHFn/mA/d08G2Vg2O
7SqGynU+RscmAGyO8nFy5SrxOC2tJWLXfnGffw==

`protect key_keyowner = "Metrics Technologies Inc.", key_keyname = "DSim", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
jbJDUJzh8myGUkoIbnMxQ+bf41SJ20FeDS1hH5f4F293JE6+XD5WLgUyZrA6Y5PfnfaK5enU3NhJ
smhzigHCS3Cb8WL9hS7CYvqwuXGI5yQEaApRiQWD4Gna27/TspJZc/rUna2nyg+wExCnPlF/lPZB
ZoUVeNbw+FveMRI0mzSBc+BaCoudszfaTloA+NvIgDdVYgD/+Ux2ml0reagSxUf7MWyB64SZSLBx
R2tSWewH5A+BP/WP2HCTqJ18hlDaAy9XTEDwuljV6FS58hhNSBmzYY5LbzwBcrnRmbDMIC9jyQ1D
wu7X4jhWkR3SmgtG1UtK++Ctz/DtJU+9PQ2OtQ==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 135744)
`protect data_block
NkH2UZL2rLc9s6ga3a/FCXEN0qlQus9m9NlW/pH5lAMyYnpQx6FV1qq2N0G2du1t757V4opF4JIn
xPgYhfHmqN2HTRQM2Y1jIfsUh8f2ZfRJbVAh3H5N4AxA3KOxM5KucF3IhszG4Ypaw/hy+faa3zhX
V2S+qrHCcwpU1oglUo9shY5dJzL5X1/ClKXOvkrP3R2aNhEAczq8bbwO95zmRAQqLIA3PPd5XJaG
LRvpcWC8g9AzNMSMG7F4niv7E573P7bJSbs1+4MhTMxNdxEFRtgWFdYELApZt9mnr6SBnXKUj5is
k2qSIxh/c9ezXmxHg/zE+F7f9QVcCB2LDsdwrYf4YoHDLQrshQd4bpY8jY3GkrnLj7RYoD/RUVkN
otYZARQYSEXpma5f3JwbHGhClrpsT9IoEdpu/IDd8RrNkKA+VCU2gIIxDGSNFb3x8UoG31g+QB4g
jHAV936ax10YKE8+D4F0WnKVE/L25NmKvw1lZSkpmprrOagAWsqpmTWnQYSMj3eXxr25i/K1Vqv0
Z8m/+WQo3cFGtahiZTeQmgIWAWg6ko7480/TkcEpgvLUL9We1TgRLxJYmWl93/F++1wWCWpnRNiw
C+tFMA25fY8mWXRr7il65GTl0a/QJ1XK6sFzTeKT8YJN/9cFbpQLH/4WunS2mFx9gNUNyKLIhoEk
Wje8vdiwW7EI8a+yFTPoy+9kZZMhwIKKKHP2sgCimbaa+BMvHR3GKQLrJ2DmrWMiRTs3EeXbux39
dpNBLlsTWzajvHMV1KYauvJzoXXVLXoYhWwOZ63Itljox7hyb+Pa25W24xxIJdf2tye4BYEDosbn
vFkVo6wyYAk7T9jpwSoumxe1YKDpwVmwdvLVLr9hjM69FTmnvGRriv8pOGwWNkySOR4yqd5WR6Hu
0v2BEV0nwXYEfI1n/pMXFAhbrFVw+mNy1bsqZW2m8TLCqS+WSjKrOHS8tgXeTx+1G549kc91vHMo
MYIXFGzJluhCIlI/NUBq9IHC5D3xiMrjOqdsMREZgm4XQ2m9X69fVBbSYUJp3ntC1OI5e1Oi7YJT
FP/aPp4WNMhp2e6jApj/AOntKMrSbK6iBzdbT50w5nYjbxvUgR1uDv8W9ojDrww09rGukfHwZf3t
N03HlojQa+bcc7lW15DjPPTw9KgHuo5LUkXka/ETRir7czCTKIB2II6JR5/GDKLoJ/Mf5Xw7g7Ow
CXKVnQs4xQda6E4OMz3PlS4m+yn18SuZHfOPo+Il5E8cWJVa1HGAFmf0kqMeoxJS7Gd97jHPqEMF
cZYQrqT1U+oRh4eUnjXc6/lr80YxmyU+u1GfCJyQrXZGv2ljRdsPZryHxQx+bJeII4NqSq/1oGO7
1kNLytb5+1Kn2c3XYWmi1s4EaMY63QocgZlH/28kQZhbjWWfn7KNjljiHjNJ6SKWdJoamWfv+vYq
22uM/2Tl8kt4I0jF/9CHjEnt0wKp8E5tOKY24w/U2Whfxd8B9QOE9w2C4M2ZXc0w5w+1CpYzcLGj
L5Co5JAFHJEk2SyKDc1qo/VpmQiXE255fgzwNkbzu8aiWPXWgy7E4BHNgEwjLkCiuV3yDNjH0U4M
LsjvbHizzMvkHyRaKPAcasZW71HYQ+nTI3jXyCMyneMH5uAQLyIqljtCsNz3lEhM6uKWxT1dGVyy
LG1Tk2Pf0JQ134MB6nUnwCPaxHMT38/IurVv27XmCH9lyknHbzmr+pdLA5KlH/Vp5YCZPf6d2rCs
pMeHtyWgTOs6bez7ATNvN8PukW+c7mnLE5mRI/46lGZoQfa6kXfmQWzZTDNNA57LA5JNY95nfSuz
/ryOcIRs6urKUczVpXmIpJHKs2ekW9aPpewp5WKRbbBF67Z9j57QtcL/M2DaqXDoC3GwjSQzvXMM
OSJehDUjjrMiDAwECCVsCwK3kNhpan1P8cVW7GyWaw10ntHzweiNeudlrw6uG3BWdNQPIeFvZB6m
crytQTcZB8sDMLBYm1lz7yOpQ+KzC+0bjdxPDfIYotewNm92nmKSBgdIxl2MP5Vqm0FBcNks8vYY
/ELAuwPnTmVZS6zRG02hb3nzIQn0euDokFrBJUU07FYEsrNVOtLui6FxazyFiF6myAFpKmmLFIoK
W5Ulc4CxgkD5Y0MSOJpHdOfIGcb3WDGt8lpQjJJ3heppL30PnvWpE2L8la7vO5iVhTaiIrofO/rR
p9pZ08a/22sGmkWFjtEfQvGMkWPBX2gh2AhFfiuQGLD9qtVw0KHXyGP1CHv3YCrwlDjjcrrj8gQq
7X5a7/5IF05/Ant2GMFKLI3+5wBzGINx+JuM2fOMlJN1/OFwFqks7sYe86q6dUP+skDXbIjKjxKA
Z1MyvyLQViLwCRGbvPfTGOT4zGnWk+8xtMcseSIyHowYH2C+XWu8glSiOw+tHU9WewjwsbySO3K9
az/SE2IudmkhxXU0v8qFxUN7H231z3z838RR4PF3jiVrfRZGMVSkFpYgaKWVdAN4AXozZLPMRNS2
ycwN+j9iIdQAOwzvZ8Vny/uk4vDgsrwX/DBMJdYXhFQvGG2FE4+LLjX6XCF4AnflL3A66U0/BLtG
38yGgTkKi124d0qoX6KdWzqa+v/C0Y8XG6C3zqyI8M/JqUat6BmYdWeRnXg2QoyHb2oHY7bLSCkp
GKrvYBhnGza+L/mlzJOhTpdijQT76usaGxfMw8RwHerCCaTmH/0cmfnlBJe9uOjW5gtYCjSrtEqi
4rfciD+fwYc45mF/G16HL/+Og8JQmRLpKuV20ozE39tPa+MI7KtVdj0KFzeAItCjp+lGAIA/0ql/
bnpBuDKLrT6s5v+xPkFr5prI9al0wg2qNE2DAj0V6Rfyn/d81DbA9WfP6SOLrfSsf48p4Oc24P/S
sqbszQ9JVSHAJRCguCCci2gq2DCTWyWAqn5AQSyLSaR6WGG/eiMlqCOOOM8LJKCBckNbdD2t633k
sVCsjD9dlxkhqclfmalYB0BMVrJgMuYzqkOxlB6SzKa/NtXMivrLe1DqM44AOpemCRjXTJquE1/G
Ri7Ewy4dRfcFESXmlW8FkOsUhakDSdgIhk8rftI65KY3rARou9VG8oDcuSXH+TN8eMV+OYOuQQCx
Au4rd1B2O9XjaO5Q6qJtVEqLKunjJa9P75UCxzhISdBqcdHP3xcfEMhUza96C7fT4zdZlLdsyVXl
QKphlFPXjwulQxSg4fOdLe2rjcrnm2OjnokMBUIowJGwkFqckd1LvtCx2KqAHHlTMyFPXeKxu+Td
/pRJ43yMA/8Ub8FuHt++iU5XU+E1A7RhWzXrl8WvJGGGyCO4v3gWvyJnpd1iWLAkbwZtw7Gp8DhI
zLlayjGI22dLsnpkUupbh9aMbyuZAXTMyxBaff08tLnEnpPZPSXplatzowhgTVnjbYuBabHc5A/4
KV2bgoHoPyb0DLE2tbAgzg5N6pf9I6fg8Ef1MKd/6ZMcSGdaFkIXooOvSUtW6mw7Su7fxnnzB4ot
8MsG3/LQP7GRunyBO8A9ezMarTybTbUi/e66+ISCoxKFT+SWiqZuvHgHqTyb6aIYOWOx3BHbpMOt
sQz3drKpbUM19MzjmBT5/glIUGSGSdflULdyzOEMcdgXJNzXFuMAGGISrZ5utqi+T2MIcCwU9/zO
PwBJP6botWd58MHr7ob95YcCBhVuq9YeF8PuQO3xPn3lxxHa1bsZISZoZw9NbSTOfq0BLLnRSRJe
JeA5j9szpklTvc3d3GW1ESUEZAeXfkUA4KXAiMokcBwZuzBeNrUnlhYSozZDv5As6R8TFpzgV2mw
hYIcjUxCptVEhuFMVeLb6LcvkzAJfD0kLUmb1xXebG/YrINOJkgJkiJ/PTt65+gFE4/Tlx93nFQE
BEjvEuxll3B7DRiQ3+bGX4orN6Msa/OKhERVzu+q5Jv9nwtf8FvLCawYa/47sZ3Mgcn+sJljWNhm
QopKvDwas3A0Do3HKs/CIATzuHtBEc3p49wRBu93M70F3yneBAO7cuMDJ24OI62SPk7LZm64lia3
Nf1H3OQxVnkCFUhG0RzjOTolH8NKz5a+Lq/1ce8rtAZfMYIVFZxrnwQHU4DIU7zYf7sx1gth/lA0
YAcybpZ07XL8Xq2Yxvi2TtgSHTojxSPWTLM4STFtsvyOa3u+9I0rQvZvl3AzXra8t+wlZ6wx3uV8
EcWd+TMCKSZTMl9Vd7gq7wfGgOZ106kCcHs53fT/FBvdMtlhju2kGlbYSQ1gp6bpUci3vPaEVdJ7
d/7R4+NEDhpgR5EkFEkEivbcxBwCdpKZUyd1E0UmAz0URHp2WEp0TAYIpKE+eTCIWXlaEeN/knEB
1FanMzoEdG+BRsgZg0cijI6lu/inv4PrU1uiFuiIPk4e3Gl2YvvujZOc1OpcZTark/XWuZrXD8Kr
/ypd6N8PPgv6mmsSSe2t3/XU5P0cMwyamZPy2htEByvpGsyxGudgVjoiz0NDZZPOS8W5repJoV4C
3mgD7kMb57yMP9SPgcFwJzQ604p2GPVlRXgUWheSmcQV4fc7Uaj4X67Qh8Rb1qqXxJ4gM8z9XkCw
U1g5fdFgRNwf+JxbbVfur6H0n2msPW1ePdz10YovHtITl0t5lCq1bymJsHZcwzaNjFwzJUjn3QHA
8+/z48uxsBUTdQDYYcmmdf6QNUZsYyasEGBf/7IsScX4i8bMBYnF6hZ4Enx4wSRg4qDyilOtQtHN
n6enT+9jwa4SmYonIRMMXfr4eaBDeXFYpdNEW0ywQE3Ust5DY9+MjPCJhlJ/nfFGdDVYJ0Dzay6a
iYjCEeCqMWvjukaJuP858qHb2hDJCY0/zZVYph+jMyCDtpAWvI3V1DhKEt7XLZGbu2JWW9bypylx
9dkuZx2eXfdNkAvS4gNrcs7WSYt90NSIbtUZ2nnpmWGQCYBY81MPZsKY+OxXpKjRAUqFQPAKUMLN
ORQVTyXtJ4AqwobeMAyeSgKsD6ecxAOvhjU2Aw63+ADChvfT8razZNWFBYd8L3gXKDBcRB5vJ5pR
+UicfeD+WpU6D8aHTKaTRuT890acHyJMKgVj2Lv9mu1Kfht91jg5GBVHu19iTD3/nrmxTDTWD1vP
RD/vQ5XAk8WDgqnV+UjCxClZ0s9zb1ug7csvUooG+qZC8E7F9z/WIRq1pdbTt6thQfaKpWgQglmC
bpV2I1hpbhWjAB1NpF6IYMTcOnyqvQw+hC6eXZfoHLhWAU7r37psnuTc9jnBHAh2GR0KEfIUZl4A
w7OlGi2f7vJnsmas/rplemfb9vWWfp7H5Y3qHVrUL0SZFB5+BcotrocWOKiSelWY8bOldtsCxCeb
4m6CBQWQK1/rZAXX5OPfxIkx5aYtg3WPMQ0l3rw2Ib4hUSTj90dvGUhguR3OzxVpICACpCVb4+TK
k0egK3GSsIfqDpF9anxM6Wa53y6FjoYaikV1FnV45CzcLmF2zaYe7ApBV/YnDP//MtnWOhBQQkEd
Vn+Pkakn+rvvS3RDel1KLvU0cr1dQbIG+GR3oMy88zDvFExxzB1xMupl04zIC9ujmCnEVunAhVLK
Vj1sSX1ts8BI3h1HFoMw0unw9Zb62NsyIot6M8ZXk3BDEqx0htMXFEHG+LrQyLzrbFyDJl8pfTSK
NW3XlY+HFdVLl/R5o9t7NXu+l+VYQfitEc9vD2X28JOF0CAe8E5KLvYwb9hvMTPAUE16vdc9XQBP
2glzBy2WKuz0qKQ5GKE32Y46Q4u5A7VSKFhox0A4unrEBLuh3XJBI0cHhzMOhi5+BQVx2YvD/zZ3
LEaLlurW6H6/pTRjsU6NMPWeoxpeyy7+zxycztktDx08pZRnrixobLyWOunH7HhxEV9/PL/36+ZH
SeJGIWqr5g6AuTKvzB9v4Q4UMmNf4dKkM71wA1mVtzAPX7VYJWdBTShzOMGFWVcKW4KQWvHc8WsC
IfBXt3Dj2XSo+PV/DgK5JD36SRJd4yDMzxJjdBU7HhrhFXeGTOhs1U6HEGL4zHduSPTNOM57kdOf
ksOgTv6QMqCxygOZmIQo0Vn/C9sp2EGMKWaIaCWMRcMrXEW72W2lBH6T/nCy0IF4mzIdZYjb/Rde
3IT83sT+yjER9TdirDReQk+TZP5X4ihR9Mgm2zm3ypldgnX0SHtXSffmRpJv+xv5FhXHvgQurv94
upeQihszNo1367Psgc+rQa4oDu8NRUQSH7HF+m1stBUFym3uuAmQOzHHEOOp06c/8KgYLFeSoTCi
iLPnAlxxsOe82Jz3hwwtnrhhuA72FcuchGy1rqxbl3TIo/rikmUJM3N7LLjOPwStwT3Rpfq4Ceql
OKyszO8SzF8J67WK6AkPhe0vyWWzumzXMx/BhsH0U3QUBYp9n1K3Vs8oz09gqYMfGDy2Vuo9Y5/K
Qoggm3fDC5zamSXc2CwDPpyLFJ1wywxWsnSuTgEesbEN8rv2nAPiLctrkOeDelH7TvP2dJTiwdS1
Ggrd201COTC+hI2mPvTAMa1wHVuNfCoNlzPHfNloa55yLvP5ljOv3v9dfB4A6ZtzbTmsy7vg9kQc
aDzqnbeUwv6hQCMm9ZQtM8RkV/1VfjOX8+Tke2YQoIQYWgWIIdBf+Yj71wrHyhLwJTj/H9W6pVqy
zD94gd1zrFCSCWoG1MxFXVB0jNv4nQ+k9cWpXJ7YjtBvhyDOYlsJKD+cs/IOpEH/t+UzZRlJDH7M
54EpK8vxbAoa2YpcNSufpVV0UTXiGgHaGuas08JGnLwqdg0ydkShH/bnIbpwKmzMgsY+mr038E+v
DL+MxMVTLALCnE6qxcGSNRwwFN+hrDPjhNeTFIsFVGt+Rxxp8UcvtcbatYpoCg/b29pxCCgKAyZB
oohF4H4PVyql2KuwZam7SdlJjHquZUiXOHXD63wKyuTPjqOZR5smcqduWZSeN1AuDMf4A+YA2sHj
OTdDmNBpgmATNndCeYuHSq4ifyypeYV2WcoQXCnIzqj/gCoNEq8bepxox00WW5ex0KQnOD0c6SxJ
S5quay7ORJY8zOq7hcC5M2mu7MHJ6is5hIA/gJ20WOzoywenM2R7q8dPOWvs2B9yA5MOe9bPufEO
izPkDhySMWGEFBRZarejRvTaAfciM07RhhOcLvbLEYGVBQCpW83UravCSrzbnPhzfpB4Np5V+wCS
JUZgbhv+gk7nfgYC2rJlP1ci/FpxqNIA4PjHaLVhajxitkY3KIl5JzIyG1teeCjU6KrfMRQQn9od
HRIGFhfXn/TxyJGIcntX7J2QvpPc4COPY23iag0w68KGeCOkNOhT9VWYVAxd6O1aoDbHZn3Fz6G1
R8jP3h1P8QiNuL+Chd8SL76JC+W8kqKSLJImKpMRQb1CY21H0PpmW4h2HFqBSG91VyZnylM1hT1G
CwwqBMMhLVFLLGQLyqxgwOB4kvy97wgjvA6TMGKq9Rh/o1SpwQc7P7r3jTbMdvftOlnsUGoay2+E
ttwicvAaIFTzglpLoNNcRUStHwj5Wggl6Iwl0xgUAsbj5O7x8Vuyg7IH1JOJL1n+j1bHxAmxWkv7
LrmokbKGVOyFv95gxWgpgFEHVpPZeBHdYGShk24KwHm0aq7GXs/Qw0uFdlbHJQsJeS7S+DHX2ZMB
eEDdOhYZUU6IF6bDGP/eAx6JMYVGPQdtlUyHsJ5hD60GZHFmuh5bZGKmVFmxwaoxbrriUwRb/4vj
7oEk4qbtM/wGqCkQmCWZ7M7BNh/REJtybuFYcY7KBaLO9RVg7BpDSwW21sJHY3qHbHWXWT6r/gMj
xr7OAqQHwWjVw93hDXYI+Kx/mDY/C3fhWibOAcC0DiE0NiIRk1NRech2lnaSGcGkCkaUDiCXVuO0
kcNFvEZE+ztzvj6WsSH8G0srd2MMeQ82tKTTedHeUt4sdt/CmQMBTK2jY7UiHPSdRpRApnjZj0nr
dzsizsfZ3B3pB8WC45iOkffRF/CP2PGJLRM8ACwE4mOvU2ZeXLPt8O3mzKuYZFxLXI1JOwfY+ivl
vSyNPVxsR5B7pnB2DBmI2uTVVHwAgfg2OQ7WjXsoXb18WqRQg7rwxXk0ha0zUsVbQJWEHrdwbV73
0++oED08nNI6ga2CYOSeKQX8buJstHrsrdf8lIT73mL789ivcyTi92x3JRR2tecAa8TbhIaPgWrC
HZmW5mPApBhBzdDMqyF6NuJYWlNbHFZzTbf+EICG8AczmpkJ/ZWSURuo0Vj3u3Jv5P4jc3EoS2Zv
TXZJSQsSoTvL3T5k7aRlHUI3UwlmwJJLUD5LxbopyO1jns36MSlSOR9/lOTZCxY32D2wZIW8Waos
F4zKoTVTmIleWThpDMyMXAhrxXNsbUjIb16vbJOer6nCVksWZ7zB19RN5GL/r/BLHRWdKLhoUusC
ejm5H9CGyEah+B6Y8NqnCsm8sXWWAJvZdrz0pMcbJL82irr8Zr9apoYP8mGxczF46Ln0vMkwhE86
FWCG72mFgi3AnnA3N7n6jU8HdBSR5T6eQHclK9RwrTu1EwwJH92A+S+uquxQ9Pb/r22IATN4cPtc
oqbnbMV0SBeIg63ymVEBGepx4an4pARbm2dju3tZVqWXtClTUENTt9vLhtFgtnEHxMt5cFMH54vO
bZO/6Vwu7fmLrmxG12CsUWWklI8rM5TJstpCR0AmQdiEbOj8qVhRiFqFoyjunm3KTBS79naNU9Dv
EvDmKPup9eX1DqZIDXBcI15grh7tYYaa2pVo4BQTnivLRz5lWfee/ZluMVe/QuVZCcqT9dZGlGQD
0nu2MD7lxt7q0LCWd4buwz5i/bLT/geV8Fd8kNZVkVcABtI3AhlZ9FOWsoNcKi7YlOwUnfSZz1eM
E9o8sJ0qEsCCRgs1stCc8Nd3exdsIU7RiNDGRPCGqF+2ZwpO1j8mTzq/DvA7TiqALp+tl1iHF122
RN7lSHDnOCoZN8qIupKlhbS1FSThzxzBPGPJe7yR2Y6lM0cKZjYAU88hHOUHr5Z+adPXtjMoi9Jf
127yS2Q71KFeX7fDKgYZBO/ZG3xocUxrFxTnzY8SYDPGoE2qbOIb17Hw00bAZ3XbAXg1+3mOo428
l4im8V2hPKYS7h/rNvydJ7kSsArB+sZ+XMzkcd1AIqcFR/aOh3BxhypehbwmkBIiMm0giMsJOupG
/8cxvgBoCHdfA4jMbtkWfCpfyWdf7BbST9ZFTkSAxy//+/Gs1oswbjvO558iVO0rC/e//bRdFWtx
E+GluW6k4Kb4I4QHZdLPtWRw+SvN2eMfCSSPWlLI2FkGUF2Ba5jR9k9oolJdW9W+HqcVtkAXnw6p
/c2vslB/QLWftfzR1yEGo83rVyehtDXd/8qJFBg4adb1YTXp0vlibdI8EDOdJ0EAz8PsfraFmmvF
uD/Myvd48VdyWdJJBfCaBC8FUO5Gwz6gDzV6JIVYi+DFxqpt80Nphtmipc3xFOSPMUUKHBG+bMwP
LIQ4RME6bPmZ/xJ5EpRsVwHthrb+Mrpg2HaPPzynTowJ/3LOdscytABl+hwZaAbo4tI8eFhRk40C
lvapgdGNR87oKg2dfC5w3aT7yrYynxg11wBgsoReCZt7Sle8ZaW40eQT1/4Jo4+/yMZV87Hf8DC6
X/SmzcRsMshCCml0dbg7Bi5wzT5tYKLW9qmZIUFVNxK5DHcGs/B2kkXGIoT8mHTH+8LFzqX6WeSK
DypUWSwz01dQ+zmgAB3tj7WG9iJNz+9RTMusXaXTTv22pIhhKCTpGyMklWe1HpmCDtrxQAGXmwv2
MKuGIrGhF+RLqcoQrqeXDJFKYdyMVBwy8TCrww0mM593lgUGN+Ux+6Kl92WR9LKp9V31IPmW4Grb
XhWw6CFCIAwPHmigs2buRwUqc3lHfL4lqGH6G4GhZTDvH3eXLcBjQ5/A5Iqp6f84jc9wGL+u3HUd
EhPeP67kG4aKtb3y0pf5wmmfShWOzpPku/sr7/2HzbZRi5cLNCO7bukQoxgEZev3oHjYxVLZtjIc
ofpIxGKxnkcRt2cMcG6c3jQS2DRH1EP3+0jxtj+9urUwyxVnc6SbsEEiGOYUu50U3qtyNDTZjnt1
dsanbyCCApHZryXNAyMTaTnO9lQdJXeKApxZo30sSBSr5Fcidsvy+qHGBZR/hLSRxyfBfWPjkFmP
hQOaw3HuZ7aYC3zxh7yt6v1fk/ekfgc/oUamPCJXmgyAeTl8lVSNd71oudPrgGUyKsksN+hCs8rO
cE1WsJsWMU6sxz7M/gga+1xrBObAj5+iUMg1AaqSTkc5PUB0DlUzf8tAUjvLa2yPbZPmTuT6Ylps
LmxxuTbqfg3dZ76Mh0IXmxFaVcdVfttnrKNWM0TudVhIq48m7TLIdkD1MNpGC9Ehs/TEBSf7/9wM
3V+hHn8S6uIf1XoF60Qs9UCJz0hqo1H8LeMlDw9H+dwztSvFO1oRJrxR2gR/NDVRmBYWzzwDphND
6gDX7pDjr3JWphnVB3J72uGeM1NBU9EPegxvztEf6TTP9boY1B1wkhRDQEfQ9M0wexPQJ/JWoRp5
AxkK9X3ArgCR20m3zClNUxili1UOYw5WxcvNg0/ktJbOLL04m1IIyBuM/7d6wYZzc7H9/s0hKjqH
P5mLKTqZeUjLZab1EGgTtCB7Z8Okx7YX/Ws5vMz7s0+bGnZoy2HDHPXCkhdxHSQzsQkGoinTW+5X
n9ikdiAzmWE++urdMrA1/Af5CotsV0KmSBdgqPQOMA6j92+Z46FQKqx6xtRtkDYzZ2OjNJAYZWZp
F1/nq9z4p8TQD/4YEtL4ecqcbih3ia6cBwXCeTt6RQEk7t/ue+sQxsZdePirZB3gQgnOk4HDIeXz
f2QbXOBa/ijpJSgkfK4E1m/ekYU9OA4BDfz/Qz2HV6UfMT2ylk6A6z67isyJLiWoF8yU51IyiwrE
S9gyuPSfQobAfTAzqzw59qc88rgbTaogtzd/0XeTtopN27XLrOdKFKVCKHIR9Nd25G+MWQGcf4lO
m223cHG8+Xi58hIxqcQACSk/XeVGHZGQBd5/5AHdacYsthgf6SyFG3QOMptunyhsPuFkhI+NmbWS
o2n/tsoJF4fqUNo7Y3KW5oGeO0lk14k5+OIMeYtfAktu8uUCgt7CpAOugECpRZFNo2KpdtkJLHCM
i3vU6tlluFnL1rvVysls0gekrvq+doxWLxy/sL2D0aDIu4CX2Xqqn+JCgzgPVGr2gYXANat0sxY2
VC3YgsbbGt8jCuAG4969pNoMsPLOENEhH3b5OND59j+EOsbHmzcPKZGErUGMm6QtBaIGr4oFd4Ys
2BDbQ0li3n1WoJOfWnT/2+cwtWHz0xPsggk1gvGvyPWWIY/5Bm4AUVcXtTJ9vS01cWgAqUVfi34F
1zDw4qOitHyQO2rxwdGzudN0w5Oy49TQzj/bO7ed8xWcsXiph2gSEPBruOGvUVLd9KaIzigI3UUL
OKdYik1RkxEuh4C5wztg9bKjsyjuAfg026cuqcrNWG31kjyRMq+b2n0EBR3iOFaiPJkSdu3ARa8F
ExDLMXFbnKXR0iZ2kYynaVtlGFHZv9i+ZliocvW8+OykUG9q0fgIDq5k9gmSoFuNag1E2A81uuSE
eo5i864PafWtwZlJSxccKZlFVrY9bHq9FYy1OEWdFoT1KFne7XvW3SHgFNuQOBx4ll+YAYNM620k
Wq/BNwR7lVrwumT7NK+rhF5UalIK/GihU8Dxviw4XhBg3I04NEuqDOHk9bkM1BV59PKrgiBp878b
IESiW2r2WpE3xvonwr6L5WVrVT9MWNjecc5k1OFjV4KksaT7bSMVhFhZdg3RFHQZ5HZzMlVYu8a2
SUlWwtGmYwkyPUpzq1vYLnw0scl7ahTbf792lp2ZGZiF9EWfQbIL3qen9iNDVgLVYhaCCMDOK/5r
gev+Gyz29VG/V1/z0aLWgeGUq7Rs9nZOdK822fmT//nGczs+VChP9Mzqe107SzlyCz7dqUYIu6ma
Nbf4R9G9ZV9ZysL2YgaQ0SwQrUvEMMzrDjcmChpQQMfEpCFzxoKx8/kYSdTTCT0DahgeHO04lZqK
8XfOQCuh4hyC3DfBUgzoRs4E6kd9Fld02m+DaoNLHeMpc96BaMB6f4UnZRBt4ChDG6R6VkHEoss6
ekLerTMX/z3IV+QsByvgf6P1a/FXpW3S2v0fn0RsroBNqqQq64M1G+bznK8L7OEii3CwuSTJCC9V
gfgyBtLX8ktwbqQ82zX9vnqlMdgRVQ47fTT7dFo+92l7KSpR+v1Ve+Nz6/77CNqhrM1ZGScd/mjf
H04WFyOGBLnZFsHI2Le1HQnumSaPhmO5jEz9cVLD6OZUuVa07ystRi0Ef5AMc4g9v49EJLppTkUR
lBmHXjfA6zMUgnPpRiIIoltZV1d6RTdPb4JwUoIfwlWUST8jKo3g/uirCGLyNWDGgLPi2IHhbn5h
TP6+OsAv/Px9JqDXqJiPE0c8BLW/MN2uOgzJyhbJa/sIPqLL2hGSxG97xkZfUlKlQ2Q/qPaG2cur
nScFnsl2CFGY3Dr+k6Gb6R7wujlRHELktxISnH5P12TlxCij8iAu2mYgkDrz5ec4RAUVC8hVQU0q
YUE7NojUADPrNeIyHO3ciXh0TtTbt11XCy2nJJvuYbTb3+Q0kQ9KEykuakqcRnQGfobUJPcZilGZ
a4VbpTY/wpsEI6hdPkHS2/y/U2Yj8a083H1/0KY9ZVTv7FGZfOgQWSIps8yyo02u+T0yi0mRsQJt
omRbgcxynFg5ATZQpic22s07f3wMywYTBjZtu64IT3KfAxBSnwOKUgAKQKk/WVdqkeETlr20afzV
p/n2OIJ5eHaToIej3FMMdb9ctHlQKiA1E10CaKYXhvvTXXcG2SoB3hlY+3R0NZ+X6Dd9gafBx52v
XMRb9Km7a7WYDrRCaVZdwWBEC5am0XPdfpuw5HWNbBXzM1BxbmJg5MS+yPgPCXtoJsAmS7//7XQA
keWTWA1B8hH7Kg3gk2IgPNreZOD3hW8CnuIzz3noej3nNhldKZnJV2T3HJNumoWjHe60uEJlOIcX
GPLySFXncAX5MpgeEFr4nHx/2GAId4CpOSYU2Gby5H7LmhNXJ9sMkVeLD+Va3XG/kjWI0w+nOtRj
/K6yIWJxrVWnf9x/uhy2168XbnWn+urw8xMGeVHGtw2+0OGdyzaWfvSinfzc8IIVuUhEoHQnWbs/
B4ZCTXHPTX1IM+LDXkK9ZYvCZzAUOvKcTSWc5fk5HPZ7VW5oNW2j1cuT4ZjJFoNdVG0vyHoBsJxg
3pydT4pU2olMFI8unS6+JXzwIyE8ArOzv4WdHmlhe/Ih60vNYaKsrLW0ehXkVkT1100etTV94pdm
j6qyTqiml1TrJ/VynOWVHUHKRPEenjLnZ8RA51e/9hufbJjt6V0vl5LTickE9TqCQNKInQ9phn2M
vr5TNbjjJJCt1rDleen3NGjE3NyQfwr47+7fMyqlYYr6KINHqyIUOawcp8e+D1wjH6hVFp3njbc0
kfcLjGCu5UXsI1Yi+i39+x1PTssAclXFniBIuRO7FURh9Kxd++nDqnYmFL07+UewumJjzsNi5fI/
7IqM8EYF/PXHDyH9A5T3HDcAvPINIagsHNSdNhrAMPmVl6t7+Uut8MPKApZ2Csw5sZeJXnqPt8Ju
+e1nKVMfHo16M8LBEufs5pyvEITadrznSGfV5tgpluWs8tyAtBzOGf5QKiL/9jX+f0yTlBWMi4We
OY77SEo4nZZRjSkOlz4q0fbUgeXgeYp8WU9DwWL0xZbPKOb6nkvEAZmc674rYgretLUVZT6axaQd
uaOKBlJrVHwQnoyi3qaVLqvE0MY1Y7FqMvH4KSvb801V9Lta2OwmCB/42U/IlePnia9nQS59DE6y
bNCywu7sObyLTBp6etMZuXfRGDgylnOjjCNe6zGVupIE2oZypdSqejm36i1zSlPtGsC5rYYrGou1
xon9sf0lmeA4jnrt9Bq1Jb2W4tzxiJwBZDkAVBiETbSFKNo+9SAKrUi+UZ+Y8cO9SUZYK6Hw57/n
nhCVWAnhIe0OSuSH1BSYpIhr6xKmmskFuUmdBnWtG4s83Jo0NjzMkg5yzKp1oAI5kBX8fCD8v4Go
M0LvLoT9eb+TfOUdyxNoIXLBzMzurAzDHdlfTnuQUR9h2pP5zTkiT2NLjSWGPpS6DOExMvrXyswO
BWyksWWyVG3WjidW0rD6bRPpwRQVLFen1wVYZr2kdlT8uQVlsXOg8KLvBNvTGCHGRLu5SLQ9yDlR
/ue6ihBTxEdRngUhZqrqVVr4LkDonSyn3HQMb0cqZrcgcBCHivabC4VkvZ+kuVphC4LW7X4CNXbW
fvO38zlrYMwSuv4H/Xl3AP50/KWpBO8KOzPK9clz/9AuekIe/PEKyJdFNV9mSsoPRIAJAgw610i8
g8u4Z88LyCgtQPGSd7lYvFUJg/iSe/+SF7wgJyQWHvmtVFQiPc91MMBa4fPXHNE0phjyScJ1PXr8
DFcLaDbUwZjdYxMPncQmFuqMTzjAKNb+zA5YAUuWfv3wVrC2c3oxZbX3cg53V91SJk2eAy5lEOSe
1fqFvmVUrfbyuxPx102TWGodKlO7SyFmpWHVUMadseo8D/YwD2SVIXm/OzEulUobfTtf02DsavHb
TOYsE3Weps14TcL3YSCcqAYzVisF3Zb1pdPRP5syxd2ISEGtRKr6Fp7g1Eodhr/U3bI7l6NemnZX
ZQKpIPiYhkc6xtVMnf2Frf070nX7NHADHLZx3QeNC5a7FCW+xd9VENI9ulalV6avl6oMh2SACTqP
RIqdCO+uy/RNg7Ahay9wHjv7z6wDQA06FNpGsWnU/c+/kSWYP1yL145yRBPAkDAL41AX2XGFenih
OJTsD9zijX90mBCcKFFibjZneiPHpHGkW3Fglo5B1n4qys9u+oWRs6aCjdBLIEXm70B1n3z9aEL8
qXENJzFW0S6TGas/dHBRHWTp7PTu9UoXwcJU+tiz8Ar30SKRj5HGcAiO0VCCESjMf+oHNpfTrlTC
BKFq8tkw51EYn5M5d07sDab5UTXpKUJYO+TbAm74S/bGsPVGfOrYf8IqMyscfboooUdiYVz3x60v
zSMXAViydHoGdq6xiiU+rtD0yQTDGmFHV/YJqdx/L+pcb6QrLMfYbXvGF2fUYlCHD2uS5x/ljK2w
z8T9Yfb5KKYAMs2z7YapeZrunVhmlwkIo3/l1dsWMLn3NoQoKWD5gjcTSjhmKBJOvhvyrpSpvwMc
7S+medWu9kfwG5lSTt9co5ajqJzdrU/3WXS2K0Ff82Pq2mVhUldDSgMpKqkpcl7DIBcIc9QZWTk9
Q+9Vcj4EOg4aY7cEJWJy5prAzlqCA9Hlh4DTzg0u1hmX+3dN8gYa0Op/zCBcYjUNvSsjoo+bftS/
DgNFOPrtr8ZthkubZR9OC0xc8zNUY56Dyeqzxa5OAArcSh/hoQ64jUIHiJjxORO990EPMUqJu6Gn
XxkojbqK+bbJGzaiqeELdwTDwHSWzpxuPqeL7DR6KtyGe7H0AjHTJT6vLrkUZJ65yyDWh7QGc90k
FOYYbnRmVMSm82s0fJQ+b16AyT7SKXG4YYgotIXHF5u+giaoBGYi6KJ/nXaCjWykLTD1m7Yp4x/c
xq2V9Jc+gR/O2dQwS5xl8/IfPaPL9vh8jc6/41tkCZ/d2ZCR+z/Mp8X9Jb01xeH2pNwpZjsvWBem
711SnG/p3oVOyYz8gIMEFVrRJXiI90ukJgC0ibb00hwkI2eiT8lP5NOXnsMPBABEVnaTAY2/8QWk
Pqa/yps69cdZgiH23Bc7a9ePfRcVoRSWNFuKsPJf+exlyFjfpiu34X844pmanvBHLGBuaoo6CY0C
8FpPM/qzPnZ7uc5vCQRshRbxUVlv5AovfdAq6V7B9D26ryu0rtY2Eg91vHWsBZo8nyFohh2w1szA
58cVzh6pI59GBOdSaCI+cUD54fFm9JkgFNEaq2DixAitSIgyJl4uJUBeHoaIHW4mG6hDAPc+hECQ
0kP1wBgFliQGTJ0ViNYxw+yN5X965RhYzZ/c0Vp3RwxXuqngkMTO+ppAy4qJtzuQQZYfsOmkOdvY
krEQwsmtP+Z3OIWgkPP4WOs0BbTr+zJNKHfwIskTsRHA7dotb6uoO0ENcy4cCmebUkGFOM1nxlAz
j/VCpw5sn2l7IfsMUrIQsCiyGjOMJW3VGzfcW7hgZDGgP2QFG7SLkn9zSI8wDhFBQ/gn6igMVMYj
8Mp2k2CtHKecCH6mMK75EUF8wJvhRWaQsKH9xWztWz6cbYbJoun58zDWvfP/J4m+GB3b255E8jDk
WdVmywG/GY2ZscjsVv652Xa+z7bpGckt2Sl74sGmD9fk+Pb8n7Cjx+YkmLpYBte4yDbBj/duoOZo
ntfZtlhshIt50qaTtqL02ehnOb0Y5dhs4koMAJzw3C/GC3JxXRLqogSQbPTg7zaN32Bm4gZnXLuC
DgI6EeqqmDKhu+T+3AMLsUuNTXr2wBxVXMKv1DrqIR8D+yBRWsU7iq2ijRBge9l4NAljH5Ea5J4O
2OGPGnXZFJsAZ5wE2aBULMKlWHUfZuXXAlH8oNMmr9wOxl4qWDa+sFjxSk5SWRPBaVI65S8N8vse
UB6yXKRLZzpyYbmPs4eCfLI8Z3agDvbrcpHyQiswg4DsJYQUYedVGovnGSixDzj6qguMh9hMliYe
dCITADdknApxvoxkQ9JYYYQhadFO/gn/9/R1CPFF7/3TclYsOI1YiFCVaJcMw5Zm7qvzrX6nAROr
l4WTmGlqZTn6xQ1AWDK1M85w6pJF5Deh/IAALzZh1DZbdMJV8NHuxe1AfRitdRrYhzt72LYPtdg4
xNVdzORgPaL0xDOIrERls9CnZkoVNFd+uMAHC8xLD/OjWDPWbCd7CUKTlfCU4ui5OeCZ7BT8KnHp
tYCJPwj7mFspsXAYSE6q/EXjGbH/HNdAy8wdE+eACjR5Qtt4Wgd2Xk42JVVB8jDkrtP/QOSynsaH
Jt5w9Qxt1e4+f+1uqv/Atf7spPh4AWUbM1I32hDx1nBmssRz2p9qt3uUCI6iNs3zvycmGF+hQxzr
i21kr/gqzr1nMT1ws8jwMaEIcN9HXfexKQlGIHoWF79M1lCHQ2lYJVXgK+5gL5U9nitk7LW8ZO8K
Sb9n8w4zcuRUTgZLeYNVG7IzBbpOCArpmfGA8NwnRmsJguUv/HT7fYIm2wuUK8DhV/YiWOMO5YGQ
1kiSxv7d6WBTqJmDGM2fWrnKd8MzmCS1c6/OxYtAfiwd51SEC9W5eQ9M34xwnp63RNk5pTvOlC57
HSWU5bNZDHtvr4GOmseRt7X0taaT+oaKkgO6AIP/1csjKAIL9cMqxYAzenaLniWMIdMzEra8mdTR
zJVUQ+htbSf9qfOWHfl1Pw9VxhZlNhTZSlwMpmn04U4vYo/USW+6jbvmd16THQyWC1mvUpo71GOq
xnZ78ewcHbo0fpDDl+DnktPT3tt1cBz9WvpX3WZ/cKJSMF+MkZlLhnNqQXGzH5W5u7XOxCnm6pCA
LZqeHjsmHQTO7ZxU74dp6UhCCVuDg9ZPzeMDW9CYu1Spcy8rQ7rg0rJW0L+vHK5n1MF6I6TBvzdS
oPp+IMOSr7pXaHsrerWsRco6aGgOxjjGK3lMCe/YXK8sESYs/2d1HpMxTHA3NeiPUStA8yJfCFmy
lhw5GeV40klfPtPALz7bAEcJn5EhdJ0TOwM+GVSTfidPMDPnwlyIXg/heBXL1Kr+Sp9fgDAL9lIe
stXwoHHS1+IogiMdfb2/VX86CnEfv8S2FDTaCrBsK9Tvb41Ah9NY9nEit8/+IamROOvFC8EkqZQy
dWIaM3tMBnoaYbotxSvavb8NMOnjReRDCmPQyfw6MlCQcQhV4PsWR4rl58f88vd/qmYpuI5k+No4
4qFK47w8A/5EeOb6Q/9SBKY8P//dn2FBugnRCWOquCKhgHA7NEsfbe+PMINIAv4alDUt/GeXhpbQ
0n8aIlATezfPzhTYlmx8TWmIziEoTnx6C8FAnVPzLT2gsH9D+pWL+5rGCaYgy3PUqpPdFFWCzhzG
9H8o7Ta9daJySFebS7NvOAZGPVmmUGNzfFG9lSsiYlQuR/yzizUAO/vML+XbAFQRlyHslj2UdlgI
NornE1qDGHhhVAhmIqLsdOCvHcIgcwmonCa17PMBQe/YkCeqsIWQwS+pyZbEgcdOV5O41VKKPjdp
jqxDKtkoQXHKROUYrxBug4d7f2JxYlApTjJhPDsg7EDZ7r8ritqPE0V5wO1s/HGgLTZ5hJ6NvETg
QAUU488Bo8fJBFuQtHSKMVrhNiB9SQIG/4cT8E1Nu/Wh6BOV92QLnCr22LV+gS0TnnFZnywnucwl
SRBakg0rJRGh44CZBySZlIE0/5aKw94xiRFNAiEdfS6JMd87DOFxjYU15uNPKw1vqmEWilAgeqMH
tljC9hjMVzxeoujNiKfMIIJu0lkyMOEvA/1Dze7YIBn8ZNA7OFkIeVTiUr69Jhz69eTt4kg7KALn
E3qmQ7B2mFXWKe1kxbANAXNEx7hs1b3+LjGjC6MIJkO/hT0duUOiXRwx+1oY7YSZw6Ku46PlvmAl
P6W92Q+WgawY3bkBcftqPCNhx4rWkz1knjgqipaL83x7aUKAJAAQZqZqu7qA9V/Y8CLdg27ZzHDc
7rJG1+8pLmOqRslUuRR0MZaE6AVfBbGYxlF8ZXaQTPMSZNhHXfIl7imS5rDnUYu7GMfAsE7Bx8Yj
iGqcKTOGvEujmy8ovi5uZdNttogeXaV+pCFGPkmZUlumO9M4n/6LvcZu5KrFkEoOmX27JwsCuOZV
3ijbtJkuiQNpiRyA67JDBGUZU/BEMxQ+4kZPXBLDxL/Ht1PC2en+yWAIzDf95P61tU9wiX3YQbc4
+p/QA0loFdHCcEFzcXzJ4pqVP7dGAGDnid/cdj/GShlt1peyrBINS4WcTl23Db7hJ9hw7oDCgXfw
3izXdsSO3dAYdS1RmCZKhqIo6y3LnfDXaYOY5QKn5jjMrkoEFIeMfhHASefwdC3XrwUlm6Gxy3UK
Pj1EsRHtFjUjaitaUpTo9J7VqAOs9AcjP5ycq40DEZg20Zy4QoOCiiOptNIplwQA+IqQnzvsiDC2
DiGT9lBgezooXB7E0U8jK7KWeRXg4HeQg3Ffrt3vRoS5+WOOQJ2KF1R6JFGz3Pam1lNj2xmaKG5W
WgHm+4DOqBxb3JRPY+29PAqlCrstuXkJL+Jvi8myYqqmq8j5xXZJE08YhgPBB66VZlSVkeVCJXAJ
2raKCWLB66LOEsqV80sxZrXhXa9EXx7RDjFd75miOHY0tbiy2Vtr7GBTHj8TIVv79iaKx0+HtDFi
byJuiAyyJOYRDZRhyQqIssRmPREDNMfi18+e8wvoUbuc5AucboDIvb2bpduFIgzO8CXWIaH9OTYZ
W6iYG0RACiViEgCI+9m9zsayffVOvezT6HiO6Q53b93ZN2uo55oT7IFXNILPzYTX3sNUH1ocNHC8
oWfUW8aDiBZhz4eKsTjWMSlyMT2M584oXv2UFsf5YxIy0j27CbAkRjKVZlj/Zxl1doDiQTXZEOFJ
1ID0Yg96CneQ0AEPEh70m2q0uWVt8uCYSITIssf4CPRL1gdBuFlhCiWj+D63d9Sv+0JlUuQxXZ+i
2GQ2wxA4doFOcVL+8gfY1nN1KVD7ohB/4OZMsqPdn/uJksQCRNiTxNB828gEF3r5xOCzza11DPIW
GSBFFDRCOuQLOUrWTRoOI5WVajOYCLZcKi1QPGu9blLWjZA+70YyANFFvtPLLHt3pYO3+oRjby94
s1aplt0pev/uspBUiH+f/M7QKN0jZ4vdT7/nEyTlzi1+BvojKF/DnebuOeE6GDJVfgMtvbMGouyA
lg5MIndxGg71QKuhhbHcJrqYz/nqbGibIKsgfY8Rw2IaBfphBCvVy4OTDAuXMwDornBJeKAINsEi
JWUaN9rTGPD4lEU3qdoTvGxxkKbcStytmW0tqoCUh5eN2oYlt6UomkdeZ4jXZ1nMaWs64VBUqGml
AF/h9SvfLnLUmqle6Wj6vf7PifObXpSAfcwnxgVEQ7Xa9Y8s+RKLLHj/jRU5ciwKzw3kzjQwSJCW
BbjBUa0r38cO9hH3YaEN1Tx3HQFKWMg9tj3najBQJv6nDku/PJF5bdPZbpNcqNDMUgU0rlCUOvh3
29WeEZh70hXyUTP8TwDxRboeI22yQreXRK2tEdiAL5MvinLXR46v9WjVe4VhfJScbVnUnN761Gf1
8BFnkCmBo5TwkoBJXHjqCgouZuRUibsd/oVaGaoyLxGUUh7BaNAN4CNiblm6VgQf1SkHIc5GLybD
fLLVa+IqTx6zs7OW3W4OXxmF2W92yG/jqBG5bi5YEwtv6/C9eSXU54v7MltAAzHLWpuLRt1+/KKD
nL8IuKr2gP7RYh/ZqB8UmNJU5l8q8k+/TDhsnlTeVyE4x1sk7RHE1/oLzu+KDMnsmJ6rq48Tlrvd
FH8KL1W3JEyf0O/xNJSAQJ4v15zNSxF9qH9Y3oYc/ZY6RUDTZEGsjF4Q/vCFs7iJEzwKUWraJ4+M
6E7optP9cT3R9Y0OXHH9caCD4WRUnbR1GkJEpK6AXdQ3+sbg9+0d374/ifsJgVuU6Y67P9595y1A
VW/Dg8BBvFTC9S+0UOAHGL8yn+2xe6SH6fz9ySy5mEACbsF2NhAXsbd8KyNl4DdV3ZCNkeqKjb2B
1imbG54RA1Cr812QMng7lIX0wlPTHervSnGvPj/+nc1teiKiKFPEUleA7iZdsxy/pPI+AS3PSdSL
vxe3sa3y1ZqXs6FdC/Zb3w4PMbKzZZRAjIWZXo7jYdcwEhUaHy1KBEEYDawv4gkp9uKe56PoEq/X
Q6vht7NHQYYtGm8/eVfyeBW4QZVTdxQdI9s3ftI8ggQbPOY3vlL1j7mIOuRZFnCr3MqMcRBhUozC
u6d4RO0IjH+Q70/ZEqDSgNZBiN4kb03JtCMoxUwpZbzu3yx21cML/oSRdv05/N7HzcaK6NwxqTj6
3j+Fe2JZb2On8OiCgXBGy10WGETebDwxk9f1sJUU6nbY9n0lsPROEUm45/3jx8BN/H18SyAMRSyV
GWhXIonnDI6W63l75BSfuLevovFjKcFDyKzKzwJrJyab2t2uhn429qPHfYa7Od03MLvrWMRtIe7x
H8EYggbtFpDpFstHhylDtOeeKqjdwGpRLDno7nJig/90VqPnXEhdJ71HRJ5SfPNxdL6CjkZWwUR4
lo5c/GI4KGdXGqtvm59h88aubNK6O9jsojY3yycvHvjsXa/TJAJD9BaSJryhpE/FnV8pEInCC71K
xlbhvbwZhFksWiEA6C1AVtCFH6R3FIIVEiNmfp5mh1GZXweoQbNaidwUrb+I7zsMWNvnxP37i1Mz
6057bZ+oDrsIZpI/encThXY41Ghnv5SQlcYw0Yu3vUDbZg4NWoq3kRNP/SIFvKSOSLFAUvHPc13W
siFgTVvrOUBP38Qx5rLZRRkUglOkhzKLRH7S909+5PENN6l2e2Rlo0YrKvT7U1lhbuZ0WRoohGwU
H/jcACiIyRocIZgjrSm1XUVEdFlMIOtPj7tx/SBPphJiV+c0rGD+fQjHopyNLNCVshl0Pj+wSKdT
d70jRTnWrizywlh4fsaD1jthRncn0v1O4PWNS1hhCUj/hmiWquFBveB2G/2AmO10ZJYEIjjWOBaa
5RBVQjiYVOSvvD523SJ0lnVjMbw3z24ksBbFsm9dYq17DfaJvt3oo85ciX4D2u47qqIN78cF5CWX
TTASTSYghC8rUziedji1U0cRYMXG7uzFTM66D+Q/3Sx4HTYxrRyNfhNddUgtBVjnZEn0Rsw/rebO
SNXGVQ5LgF+QakEbx5HKjlro73X/33kNAFXMIHiJZ+6AfzMBFhcr7ph+3hQkVVhApfMbKnHtCNuw
loHnWiS7LMra9cwBoIlhLRFHpaMtaPDPh0kdO/Ln/TP8+RKYxxNxF+XX9ekIiP4O5uQbaTKDFq6l
gIy4Ji0h9mIcei1W4RBwji71LtCk+vusLYNd6GpnilqRCR6LFgn7t7KdD4oAa5fEEvte+ij+G1IP
muj6N++1sgMgvMEMK2PQu1wk/RdYl+5kJGPVNKlmkC70mD+zrPzOAHKJD3C7DF8NCvYn8f8YG6XB
bXlKlJKEwMRP9xWDunuILubZQE6+qaKdzQdv5S4qfk+qhUhosz0UFfut3/mkDKIxvafE66JNHKw+
gOySpZSzXMojOKY2CIuPrdkBfyHyFBv80kywGmOe0xCSWXVe6GMc17ocdo90FqDANPYwzyb6bLSH
pGQ8OSc+dIZO4WWicLoGT/xiCft+pGNpJa/Jx7s5uqZ7uzNwBVPLW1J0r60z22j0Bo5rH8hkyePo
sq0T/WUv6chSxfKtek/bGrnVpn5n7TqiLUsAFTYMyzK9CGB4K6oXC6aFPn3cRgxhUg2r1/sFMr69
3eDCpl5B26xa6po5kFPmCgHLNnP92Vj+2IaL0O0h+VlvlaK9CYAbk3jTQ1ovel/V98fldn+PXPqK
m+YzIIZ4SMfdeRXqN3toC9sGdav3bltUsFKbyPRnfvjGN2+a7Sf74jpNJLcKaQ98LU0JcE/sjAK4
82hEKnBbQ1sEV6ACq2b4e9Q5v1aBkg3oOPIUyX+eExm1oM+Dmq/q9wVPtaOJIloijkayPiUd7s2T
hGLR/XQ8uNYstKdE57HHz44/NYFmaYJAqT5CUwIbXJkvr2IIu6hUAeV0GF/On8vfB7RBCQod2Lgi
tzafF1vUw8KzD7LyY5KNmJ5g7hDZKVPpSIZWh35U/WAEJF5cvfb+PK+WfumdrByNfx0OEmwsRcu2
+PPX3kntSxm7BAqjyuVxiioNAigQCOpJExj2kSdQT4pcBmZVoOxuCzO1qM0OuWR/Jn07KG9bN+EA
y8W+NiIixYXC7azs1RBEFTqvmf/1OgcY/WVt8FEOYt3jjk+EVyGJTYF/EXMZiYt/QRO8mV88q4I/
Oyg8cfTK4U3F55e7Z88MxU+TnOZ/+W+wK/DkxAcH3EgHvPNqMDtmIx5i1G5sT2Wl+xdInkDMPrkj
CF/WGo7k+CLgoaqdvMTs0JTZ/EabMOQqjGFkL0QHMWRcdN3XjyV0iVkb6c14FjToweXkk3dTa/JA
vnaB1YcDnWPgmNSse+PsjNTNBy9QlJqWw04qK3uAQG1BbT3OXjme2APOOngp2Ui9QzRYCJhfOm6q
39ywCVUgtqXMi5k1cafVm/mpJgOjchR7Fd8svfzclpHZXDYy//ZwvIJxx7L/Z4cdlQoCylJ+4DKX
i23eHrhB3PItEXpnoNhZ8CghVuV/4QJ0SsPEVZoBBL27+pN1awXzFWRKCG0HRGSvenHdJFYkSi/X
jUZNbl7+Ioiwg1FY+3nM4mzIF2D+HOceIWac823Ql5pFz5ZGEuDcs1vR+ai2rpMtGZc8AJ0DiA5X
rhEfXGHglZFa7zFfuMdThFH1QJsC3GxWSfZLcIUG7siNbS3MCy+Qe4KC9p9RV/nbLLNxj2vvSoIg
o03PSnX/UJcUE1tfgxbv3z4wHSIw/wkikTHyjrLs7KMP8d3ZrMnU/rUodpo26YRIuHY9kMpPDOp+
AFMfmn92hDA/r8uUtGikbKXsrIPLVXpinBLa6sY+5j1pINasz0W8a9ea/I+LBy1Zw9trwO4wEy8I
0ACi4i3I9sr7fMZXRaY9XzoEz5YAf6k7KzGwLYB7E0ShWOH+M3WRWlyLRQtahJdD6C8wJCPfoAlF
mk8oEy/n4WQIaJeSNzmKvsGPMttJIyxCkgO+SyrRhSIfrPOFdyEuJWiwYrFdv7KGpEZ03L2IcSJe
4Gjthyz3xqNd1quHtfylzDrcQE5IERjGSIJLTeGNrcy6DrdWJJsYCU5gbYrOadQYUyqDEdxxDrBE
3uE30zxGu/YUSeE+WwBGUZ3J+9snJ2nhS/Ep1od0siKIZWLtEhjlYTpMHzn2wfqiHh0kTuVU6Ru3
h0TRHK3bbGxuhEGHzk5B77g37NfM+TC1m1+idFnsI1Nb7jpM/7CdfYc/e1QcSYqBVWUcJuxCm+Gl
XqBfg73ucQKpti9gRR9iydb+25gOa9zdfP/MIJCjPth91ZHJ1CH5qDslvArKW5nr6STdAsUeFWaw
uwwVs/cuvK8iyHBHCKT/LAoR5M6TrNTbokq8o99N1hhTxosBShVLIOEm9dwY/eLWze5bS56yMl1z
OyJ3Ixlx2NLtfwx2ZrCDoa+muo/S1AzC0UJj7XNLxZcxwEGFX9ddXVO+YdiZvBi6cRh8nSlBerxd
MNiDlBnuFtGx4AMZjYFGom3YMCVVwW4teqimrR8iOnCNV+2unl+WKg8mlTnnO9H2HqRvFMeFMaiH
5L2Uoz3K68MCjWeL8aSbMH4dVFiMkgDCRkmK26R2NYFM+HquOVbJKJ7Vzk7Yj6/06+JlKrHZOHIp
T6C4HDZPI04Gm4ez2Ik9MkOsiJDgxGUOy1knHYyQgDGVOIHiYBGqLqPQToabeo8ucFjbB9DqeuaU
12GTPtxU9dUICe7TZBQZ8n3izuiGwkIzOvlUTQQd2YuHW96fVJIpP9M1CNNKhXIqJ0yDtNeTCxBb
isisBf+LOgFIqTcKDtWF8AXR1F64Worql9iCv02hmQ0jcQFsqXsLLybCM1rQBaLlc0HbBkmHdvkN
2sukXt/Z0W4BOKvQI9CKha2iclOgwK9ZbW4ymUM6Uyz13+1ZHB7JZUwTdCU56MGsLNRj8WJb22N9
YfF5DePKoj8qvZtAbn3I0PTlV51l8UFIAu/d1CbvE0yklAZ5Cskb6JJ9G5ewSAU4GC4NIkb7ZrDm
02WzxyRSb59TJTMTaWLFvbszun+WwVFYnZ3gfSBKqcl/6lmElpzrC/1UN4/QA/ReYWbAHoQ6zLb0
SMoMiWtB7xWTy9FQvwwO9DJxm/4amT6tOrlBoiNAmovgbMNvYDVlw+Hx+XKqQglRsYvKfhTqyo55
HGX8D6km9evk0spXNA71W0m3OblBI+2rfwCAVPd1t4591mXAyOtqdVaOlhzwIaMfJrVP8/MTDMSw
6KGXIWgaw0YX6xKaEfcagjjD2MQwqqNEhQvWZErqELoobesTJ/R+GLQpi3oEixR7tn5cTBr1KtVv
dNSYnNdFBf7p23Vtgm9OL6nIcgbtLa766sIBf/B0hb/sNNPiR+OcNUi/7KxcxujbJsDbxOaxOgLi
5PGOxcVbKWuM22FoR5p+sIGzzfxr1/Q1A371h5zaEuPWExPVUupLqgeGQVqrc/AV+0uGTL8LthJw
6n+mQLGLDyQ30vyrc4lFNKo7Xt7WwFAI9ZIgIMRMK9rualNv4WlQhzwRCYs75fe9zgW3WY5xf+mc
7r5hAfe7cIC2x00aPSJpPWDSuu08/Krm6GiAJf1zcx49TFEJotcwdfIpcl8VmBjStLua90umihZM
S5TeJnreI5phRgMTG89Lne1mrDXd6Lk6v/th0FZLCGmm3RuOTmnC46uag/r5chpM89GoNuoZZ3LF
5vc0KseFpBcOOqz/sJTXigPfd3l9PiMvlFcFLjmtfqyt1cqKKxrw7z+Gu/ym756t80RLB8GOUzvs
8YX3xUELo7xJ49fsLeJK0F/aSYGQYoiRUCAlKeq8qLyn/+vZgyp0UY1SYuJPEGyf2HeWD30y7YVl
yIa1jT0bc3LgP7e32nSn9hxNk/FvZwyb1IFF81cvJ/UoO6/FAjuXMIYFtQ8zf6R15YFRzgbMK3Ai
/AP0qvHlhSltaVyvR/XuPo5u21SHfWxwKKsFTx2r1T+A/v7lnrF2jhNotb21VuqE1/mfvaTglZ5q
Z/RijFEAWmerqlcupJgPAdoz8KW348i4iOAC7kES/N3Ar7KiQktgH/jdH0h9bupIeLuLk6vSZPdD
VR6TdP54NI+1Jip530aw9HUA4pF8VDQhdUpk5U4liHiFmUxxaPV3gPqVQ4/faZbr+EI7cxxS+0PK
aGKG9CTempdEkuYeIEwtE0JIWDlHVZySsUdlSAT0Wit3MOTWJdRkkIe6rB5zKJ/rDzUD7FzSNYIt
0Gb6XLvcx+zpaSP6HCVtLk82mCBZCH7IUcHBeq22SOldqDEnpShTacr4/aqtZ+J96CclFbJJ+Cdl
6+MAQe5AeFLd4YD9PqdqzznBlEcUUpg44gqV1XSNj74GPqaS+hMspeyrZG/UIKco7zSdNlNmGKRe
F3/RqQQSCCg1xWf2P1C6RkYWR/lr2aHsA+BvNbtNd3IhPcuQKdMahWzXnMfK4kILZxBNd6Yv6XgM
lbUkbA52m8gNM0xSGf0frKiYYSyMz0g6wZnDww3F2zJokyg8v0qPA7c8yM781biT5UtG21U2K9ca
OW223j+sJpbi2YVXouHKuV2P5ZD0ZTS4nynZj7CqRmtfu6HGeDxfIJgLKjH8U1ZI17Gh/SjkzUSb
WQVm6tLCFav9grsx40Icqp6BSPrSAofuu/bxKMYCP5Pm2f6eAItTMcw1mWLDBtAf9JZwVvLYTcye
x9BdCb3Vw9Rhl7i23PsWIIpRUiL1mq7xb0tI5AM+C7pB8ABZbm+1clVcJY5/+D+zHYuIv5v6CYOA
RqAHpDHhl0sl/roynG06D+MHah1o6iJ4aZEVWFiAm9zwwHd/wL2e6qaqXjy/3TjJdgX5Zoa7DLSb
3esU3xywBPiQ+9/5QFH/ra0iV+kRiJtJWbGCgdgQ/OvLDa8afaA9R0DpyDb84QVRXcNMQRcu14jH
XHrDvTbOSCcqAaCXicuvFz30bUKXW6p1sBADsMvmO3SgxGvboSpMaeM6MWzYPPlKi17+jVNWWMz3
0qbA4AFz11detV3xX2Qv9RRDFnPRRXGJkS8Ob1NTdsutrwdzPPBw0bwkpZB1wtfvxeQgzTq2e78C
NrRYfFR5aty54IitBC2Ga4tA437gBrFiVkNXvPw6HQBWSAEguKvOOsm1y9RSeiHzTKol1oah+30I
qeECKDdbbPGKtgrD8ruqQQuc0/VKf20hsTu1laTxsqf/HpozPmUi3q/1aNCMl7Ha5ntaRjeTAwjD
iht5Vn8pTxLvfVawXm6R/hrcaAvYCjl03Rj1+4i10LwZycYTGn9q1b5TyUi5GJ1ZUIrBwufTTTMQ
7Qmzd3E9SZtCxEZnzlTFFgHQXsQZUMZdxsYGhK/w66j/50vxUb3sfVNOQiTu7jyb0S6hMy+j9ao1
9U92FxoZ9GMfNmnAGHoZnNJkemEKq9SbV9omMuBcO1QG8aGiYEyhmdSoInFa+M0pZcPBDP3LzaIV
lDXg07BcgKwN+pLeeZcn1NsI77hmnbprU23u4pTCHDmy6wE9wKMLeUkrSlOGB1m9c7/5oEDhUBFG
QlHzuzetDk+bmKc9WfsFy3AiUOBllJekhuJgDF5X+f7vbHpkahlEvn98Xz+811xBaeLXimbb3zdI
roXi7fS6/jR2R4TuSUQYeEfGcT22Bcxp/qxFwzXCLP6UYrulXEMFLDhYn6CydsgVWJffOxT89P0S
S/ehDFyGbDwuNEQjQEgDXxFtDH/0gZG3ZYzneFlDSiXDb+aYyCP3PROWvOv5v1Loc3fAp535PKnR
rHApkyaUd1gtbV/VQNrHU7RLGG03/UMRJNgcug3z1z6VmnObbTWgBiVllW7LsA9qtsfHz24Jjxab
pw38NwbGYU+1t/Wdby80/V7wzvROJwNt6uWyW9yXCt/SefA8pCGzWz4OxsSDxKPJOLlx2BtQI3Xj
r1aV4zb/UMKtJ57bBEtR6miwPL2kzg7oUD+LD2Gn1SBCNX7jOIed4q7JjmxNqxaZer60nAnZjiSh
cGlcfyrrQQBfn4ZF7Vgt+ln/cchU7LwwU5z4rGfX80J/rfIcyj2ts0RZ/LvU9DwtRoHvmOmmtPEq
eZjTwrRUb6B+fZPOMQIrP7uTUo33aQ48ZaIYqln27FxaDo0iCHZrKiWIC5AruwvEbFt8Pcy4+ElN
ne1wVOyq9bLEqGFmgaTCIE0IZWTExp4DhhL45d1dziNFWFZWFLPLQy1xAZQElppDT+NzQxtXro8G
4ES93TaStoVzfMO4uTr+I5LW/tCYzXmNBwO7RLLA2Ybel2v98YvXNuYfaabhJ6Fdnl46UORC/lQ4
Wi1XSR7gaBNZC6qOdexAc94mqtvRNC2gRE/+D1uTzBcRSH4qAXw6gJB2tkqeqjID2pJxJGlXjhJ3
E4qwHIMIz6xxMMmb9CqFRnGTGzpGAb7kALsS719YLqdwlLjlDh3N59rJkD+ePZEk/K1vdpUPwWKO
YFHOrVi6b/xpWstwstZ7fgaEnq/MYmpmtIEn7yUMBC1DotAqVzb+Y1hUX3qS1kBPvefzy14QWRZ4
GLOA2/CYF5bvu6vVIWlP4MURkxXZV0TKx1bzthDMblgqOReqPFIwj181xHOJ9i5a7iXQLb+Sm99p
+FSw8GOE1EK94inHurDP5JnmWmv/qrPMqwZFUScRthIo1qNZHmtlhdVBXvLVPPHcep4Q2a9MkJAc
yZrNzsTFu3z4+5nBgbVp2x59pMwhjCFgwgbwOaQpVIGx7m8+nszyallhQLP7xekKQeHYj50NhHTf
geJ8NKal+WiwG+f2y7QnbRAGo4HAqA4gieX20xfG/P7ogJyhVtx5A90nwL4PClwU6ZiAEjgsKcyA
sVIhAy5xF+EObDVGAfNfVHd/13EfnPb8zOdI9kNktampLOXMZH5UlOoE555cbWQZ+6jmHwc2G4e6
g5Yb/ANUqFlk9x4+8KwxF/kvO/NBJ10pMmyNsNSxMuziHf0Hc5aQDnIeFX3Wt1GufH24qiJkvkp+
PhrZSobUWmYjcBVLrMH83TH67zZfYZ47JBX2Oz4m5ceDqansya7txJc7PVSOA0sLDrO/jbfX11ky
wOvoBneNHtEt+pZjIunqmXJTBcWM/SzYjv7ASvaBVd7a8l6RB2xIGvbZQ58SMsK5avA/3zZBoiR1
RbquBNH6+b1IESgJm5FBo2vV5J454ADmAj/BYqbf10YQbCMRrHP1ryjcaLiEZEwQA+LhOAMikU00
HTWd4mt4bDlta5bEj9Lf0m5kxfRrWNSkWMLehmZCSOjs78gSJQh6doKDuUIfowzDRAqEU6vIs6lb
jkNLonp9DhlEYjSwOFQeSLHBlbx6xwrGGEX1Y75D+7P/+1Y6EfWa37GmkC0ZCNxZ3Ni85jRnRPAV
TmwI5yiJI9W2jFvf6i95bzcAmi2GfXso3SpmtFj9AhIbAlYDfHwyqXEpCYwrtS1T4jQ08PPsF6sT
/rpNLdjJM79qccep/SkUnrg+HROrCB5cLVy/VEEVU6DqAaD4fNBLaAweA2F0JRMsGihlNynn/2aA
R82BEum3NP+RZh5dJf6q/4v2b4YaGIAInHSZ95Xnn+8ceDoi1bUMTV6RpaIcnNtfRh6sL9YhVKqy
WDTI2hHRF9DdVNMjaOfw56fm5rSoSDiGrM1bkb9t73gnkoXGtZ7QTTdvNjFvSHJdm5iIEzkeI6fb
O4Euj+7oO4VeH3D1fPeeOUWMwZ5HS2qf5AEUTAkbdfVztBwOhdeX0JSyOQ5zhQ1oykyq9H5+Y5D4
sLu0UAzeQFHK+yebDuBFG6drO6SvxoWIqmDK+P0niKWSkXSSRf5HFItT4piT1Z7Zv5lMsK14/MH1
5fVW5sk61Fy6mnxNSS1WiOXjTWKKDWXwJiVS0WMgue9/48RROveAt61kbnd8AT6KkV1YhSCi2aJf
jLQv1vvHl/mL3sjySY72GpwWQ8mSOdUfcJ6pGA31sYvYH4zsoajc/jpznIHgjuBIdvMRR/GlJiIL
dOXtfeP8Zm7IAFXgtdJaH+j5nwVG829gvtM1korHhM77JVVZh9kmbZqATNqE4piq3QheyiJPPg5h
lRhLib1NFwwT/T435IifhNk+PQNgHz/DFT0qVT41J5KmAbf6kYtX68ONTclPAwQ8vPAuCzdYtcjW
iEzGZk+KvYCYR05CPzI4zsvn8JTsGAHusAhmIhZZPbNt29GN+TCDvlX6+Mn33V3H+J8Zt3t7w0XJ
f+wHTkrYGXue0MZxeWGCMeBjg8LhsYp5cr9rfeNHm7vW575YG5As+LKM7ePFpS2yBXd4QjvYIxtZ
sFHsyj1DDitIiS5rUHwRM9eGR0WV1/ZY3no/ovo0N4+oZD7jxYaRPG6Crc8U9nxVFUIbtcpGjQ0G
luhsDNntGWTlKbaQgJTMDDgEJ/V7CmWDPYbE6wodg5G3lkU7R3F5GaERTmihrJh6fonlRvc7I7eb
kmiF77GVoLfQR7EXTfJTO7fNDXxMSsyOMK27tuRujNbly3huimWUq6L4YWulMDQUjcTyhtz0Ijw+
ciYFTiuoN/pBVEBCX8B7L+eqHgflmZpLnB98CNKJX4kh6mWgonkb7uGJIhouHtuAkpK8tLmgUgdi
S+CNahcpswnvZbkodwUUEnsEt3X3c57zwDdBysQK9CaDKs9eknR/hpP1gqs65uAK0OjrEdyO9bEq
RKyvqw9brvUHvqQDsci3JaL6M29E96yPErw2GjSwR9zwR5tBOmY0dTkj5T8eTOf9su7YzKiKT3Mo
YPhJjHvf4vwKszOyOeabExDRjdFayBjdRKNkcyZI8lnE6RC0670lR+v0FU7Uel0FEHxa7H3Us4n3
qqTGyn3Ksob0tqiPo1SoOX262nqMSne4UoGOODTamSX4bX4wfBgeGbbNo3kMLMqJ1FHBkLazZs2m
NLkjY0EwP0ylpoXo1aPvuoASQ2wD3JjVaD3WCDubaQmLtW5ORpkU+oN/DLLxP3GfhV/Z58lsz/3q
ikWO8/TbvG7JfA90SZ7Kbbpu8FTx3zbQ3Mn81cUL9Np3QdcfnyI1J9Jjo+1reeubKE2MtkuxiIFH
+QFlowRRvr3ReLydypZHMRM7hI6n/T13p6XIOdZzVDC/mO1mo+HgYuRGGMlh8ZMZKqaRtJfiFFed
W+2n8l5MJb4DbWfcRGRvjxQPpcxic7/GXS7qr1w12wx2NsyLd2e/JEJ61FN9Nog3NgkzkfVluXUO
hLhexoXxibBMN6vul8WBgkPvxO0JlQPknw7uFpK18ygzEABoFwDGldVuQ1vI5ujIhR2HI1VjQB7o
8OT6+XZjuoA4I9VKNGfEz76Gw6sWfuJ4dJYLyYyTZzZ9qwlGZoTQQ71ELjKTEEmTnG+WAmtMjVeK
y93uqmr9PGb1A6aYuNi0ITlkCnLEdd9sVUcARZA9pT+MIHEeRKVZ/ii41/PUFKie2/v0WMRgTo2O
T9blP2JwCmH5NcbT4EkffllYxk+Ti7jUZCt4zpzJq/2TzQnUzVlsw0Z1XjHSyabdKGkONQjmIZ7u
sx05WgZqa6ht2i+xKmIPilHOM18/4zu1U0k7Cio6mWo3EFN+PUq2FywN2jRsNkFXDwr1gn4Zsdeq
4+/WGZwCZ5mOZQuXZpAekKU+VfKxVImsDWkJbIy5Jw3/gpM/tj2sr7LzB4m4yEJpj7ExD/boBS18
bCdtUOKKq6dDZcmx/SL01/c7zdnzXrtiY6OnielRuh1JyhmaMA19XFA63UANJkqMs76N0OMhjL/H
4/PiHzSAyX1qc88Jc5skuv61b1aXTaMAFazdUCGwnHdEGl7jZI3Ta4C9JMDKNfVjaUAlihPujnuo
6ecIK1CKNhtHAH845jdSLFmJ9AkjWARxNXsXKcI28M0bBd2JyHPjVWgZmKTp5ncWgHwd3SQ6YeBj
1IN2k13SZMtklIre2v0+ImppU6I2v9IniINkRYB6fT9OjkG5PFqY/PR49G1AJuWXqRruZvv7Sme2
OWv2c/EkdV3FJhta5vP55jN2RCvE6PMojMqrMbAaYA03+Qzy09w/nu2ZNu9XFHpl12TsvIE0zAxJ
5QEc2FA/iHk++EDfKP1FH/8ar3ZU51a/Y0o1Bxy7OGFq29UwuZnJJfNetZfe7QqtTCyJWswu3UZr
tQjDX7AOBCN8ThJbLmCbDrvqtbqls56peCubRY3VlMfVtuzAeEjKkTywOOKZJOHuqYEZk8EGrhRB
fnOggwiLStNm1pjaKFHJgGJfgR3NCLK5aQ5trT8KbApkDTVCs5Rm7Lf4v+QJKcRW5Sv1Y+CV5Zh6
bdUgp4s1e/W0liBBkKoV4NOr6JKcog29qVjQVygy8zE+qL5Z2uMqpFw8ncN0go/A3wooy34IANDq
twEPu2J6XNkkEFZh8uMXNZWSRC8ZeJ8KvpBHEIAQQLf442EzPBH4veyegvrXTyHw+DTOr9/qg12e
Nvhqud3TkbUSe7MXfSbAYQW+sEUvtpubf9VRpnIR9EMf+e7Roa6MktLV1fKAFEwZ9DmzZlzBsdAH
S1FgICisrALPSQCNV6uKYZpyWQDMx0hNJhMYpgWzCNm4Zs+BJSlZdAzGyl6cR/PYQuXefS8AKPK8
RI+onjGWe96wXNPRmQ4qRVwVfStizXavnJ1zSmPpsKN7xSsRAby6KrwDleFXb5PG/Woc880Suz15
uYUDjHA3hmMcZZHWFsbO4Avt0nPqFMPOol02hCniQ5HhWZya1mdHOpXXcDzUAhpTdEkYFHpVgAsZ
UAMrExmGgnIslnV+kG4vWu6acJ2iEUvWtsLH/WVp1kjiXmwnwZU/kGuFDOA+JbelJ8w21xE9KdXy
IeEnQI7z1UXo4AY52K4SABbzKvKivxf2l5ymqNTcgjd2jUFTUeHm/QplUJBXKnxm1FEtO8V2VqtN
ETL9KdsLlyFhF14TOlMo3aq9BQpyYC4YBzQzXFdt7eXzWSTWpXk5kEWIuAlU0aK8NZkZ6L/KRcsl
9jlmsGDjK+upaTgP8q/ab/ZX6R+nMXEorputgaBQWo1b9XPVuuwpMhWTjymTo7/qZ+A0SZbZ0FFy
OSjWkwd9AlDBTwzoWJmrdxcjbHNJVQUu+IANjz/LOsHYdYlP/2Bbho92u5KWwzFTX2p321JTzdVa
B8MkrM/qcDkCCya3fRt0eBFkQM/Q46WEjJBIqPZZwljOhlLBTnKcd0cEU2VVy0anl2cLNuCxUJKd
c0JSr12p72DHM/eKA3eajY0ELDA1EysqNAtxoGRWBGk62aIz9QVXMFbpPkAROQUe5mUQXRVIr6O/
u1AGhyWTfikhDqVcHr+zJHySrOsNsXzRYwzGWaDhbKoFiNtmzONAgk+VGhVvuhBKbKQmJnf4Q11J
lQ5FMB2eBfeyyEnk0qjaT6lgjoTAomaII44SkzxmuTL0rBDoM4uKfX8/PtPpeIODKoTpMH8euR4f
IEut/uyhdkLhJKpJEjm5q4jh8AycG146ckJS0bSCJQHXqCkgSXd0R4EkoHnRguzIRt+6F5AwW3IP
knqUpprOmQ+48obub7eqyI6B0FqQbyf8DWR1a9xj7VYih0mbCwxLZ+uYaiVLj1rBxhwJ5iyBLFvk
/e4ulpfzbisDlRHaYU2kpWDbUjh54QqtEn3wwretquLB4PTcyV4PzSLH/36mpTQzpeUr3+G0Wgvp
e/STTKLAKuNBr/zgyV2QdSDoGS1KebPcj7a62xJcRxZoqyDWXeO8GSCDWvsxwNSQobdNMuX8gwFp
oLagXU9+4B9Dslz34Si5JRq37WUD+9lUZVE6+cTnf45Z3P7MiRUzBM95eLxbUjrFXPvsNvU0z7JM
Xzo+Oer2O0wYeoT4VOk+Ji6UmSq/bRalPP0W4Wt0CBs62+1G/p+CXJSzDYjJWLJm+GnxRTDgqe8E
6IL5aIoeIiGkvYBDPIjRZvywqzzEKuI0gHCYKBua5Q1j8jgONWugFJXLSqAP9E81sl4D+EPDqOGi
2XkzL9IJfdzj359GWeKDjc/8NmQrYN7P5Loc3sX8k1nGfAunHT9dOnrOlFXUQiqPqiV4CtXAJePU
akhwmEuA+jyNeuORu7EW5XRU0Yj2w3GaMen0eTJvwHH0fIVK8wQr0ilf8SXHQTdWWkQxFFCVA83l
rkDErC3ApNHZu0vmiZce+r1KTP7AqUorcVt509pjDSJ0dp7NqPtLS20LGsrFXSuTi8rA3V+65gAH
x0RwygLTXz38OPkKvvE0fO7mnfN6XWl3Trl8eD2fUvE8mEUQQzoLPWVHBUA7OqVZiAkrn0bfWQ1B
gHAxpd3E7uEQCMhMDlmjSjmp08RXWCXu/RukA0e6EJ1UoupAKiiwJNxHyJyq6xvSKwYjogkgbn3r
EuvsNjwCJGjCisGL1HD0Ih6CVaiBFnEeur1YTb+4xVz46mnvm0/9QaLxnQqVU1ieCnWuvxTk6tgY
a8BelZfMLF8vxBy/ILMHVQK00QlBPyqvlzZKTxwb+/4bgUd6J41jiJx1yS0bapRKNlPUaSRtb0Do
dG+W6esBcZGtfLLX+ivghc/IzNjj+xTkt2Sk3kvxuMWFg9A0oyVhT/3RHBprYVwaciD/ctZoENYI
4xNUlkuk+cdiR8aDcHFeBwtXng4DwSoIREHxHGMUXLS5P83DWG33CfdTYD7poVtsE418oKtuNk8M
hVyWnbjfO7KpDzDFupNiGyy8SyFSyPvd/0ToKLFGbhFKmOTZzMoqUZlmIgNkIv8DpHPKgbqrNtRt
l7kGY3BcOwuk7BxIzlM5DgniVOANOgRJFegbJqAkVBvSSyDpLGjfGqFqePqbbnqL0mCPipC0LoPt
9i3SVFhn1XykkPy/acJ3kbIQTtTGav6SrmiTz1SirjTc60G1repl+db8qltaz3YUMu0UsH4f55CJ
dziOGYVPqUj4CcZvu91j3J8EtQnMZMJP5Y792jA68DMPKZfu6uk2AxIL+JDp/frP4uykhtNcsT2z
3TabGW5ggvbeFLvLezVebJRR/YnUW1bYW53B39JQ/N9XcqSUOchQDBr6OymtBa1DINkniQNnb+do
4Zb15tP+wNcevnKbaWkH4BsWAFJTiS5t/YkwtBAUhLLVHI7mOb6vx6N2pp+pTPurUjZt2lrvjY0d
25QhEXo4L3Y0Zihi/6oNB6hFEn2bexG17KR8HNlcHA8XZov+9pQnwcKGf61KN2tzBBIdJjOCnZPp
KWh2WnOVIjexeBebD37Usuye/bLO4hqPuGiUxxOFMiU8T/KYBc+/S2kQlyVNXrhd80vXs2l+D28a
vSQq/28FkrpT3ovvNc8nHlXD8OfdXhIj3zyVL9E1uHsazUR4r1WWJReJGlaSOHNj0KGyjpVGU86E
c06sK3N01K7E4pljV49qGTJmXxGH2/UB2EMfPh+6v9BtBfLyUgv4gBZXtE/Sy534ppEv3khvMa3v
UNbp5WZqu3DJSdCFYblq4JuYP3eU6FMyWVjE7r4Gw/ZO8FudYUeETFXkY5lasuM5ofj+cy2QSr81
FErQuJCJljvzBXfPP6ccGdV8lU9LQ8jJ23eL1XUhduPiw03UWshgxCMJUoeazBjv3e+YYvAiuLGu
jyAQEnszgQqu9WScdZhfiSQrr5rMW2kvC3EYUiz1BxuNcWDUyx7hsiCRNSL9Dy9POb4dUvMGbpkl
ru1OMd7islQJ2VIFxDCU9kVzyKb7pt5XsZS68iPRmhFc3CdmFBhHZ00D9EG2N1cFN+qVCM0T52qL
HkjALkqGPxdMjiWDDjbs+C/GuYgNzDSK7asFQQ+pNOTsN012OeiZXPFwI4s3twxxjjnz+YNDrign
vQoQwAJLMaRUKFAcg7kglurHF/uBVdON6EZCmLZasnapatDpMbsPq7L3oGQ7JRwCpKfw9obTHkpq
v/oqm5zOCGv49c2ht85Oc5WbzwL0I3X3XGpRSb7leCKltgCzWAuPL660lENkf7uy8zzLmTbF7q3K
REWGUPJC4txgw4uKPq9gHZk5l+U3/vyLL9kFwk9xWULZNJ3nx7sgWCVHUft7Wt7ZGw3vaeUHEVcF
moxSypZP44f8QGRolm8Zs/HaoVFDUnTwgO+Tu8BkGcvSlli34xc0nnu08LcPu5uZK+RAzgtOS3BX
K/YrVTruMVzkMKEcfSwA4cUU3NepnV1TMqXczTjl8hlo7/vmIh7yr+zN926B23dw5RAr3wFXEHGn
NZnM4p13/n0ocpjVPXwWg7ZxgPTxoJcMsg2pSN8FdbK4HpSkv3t3vZnLpfkuMoZqRJax+KTWi81o
/iGnFrradFsxgvq9z+yOzwaAzroDQgeEbhR1eBqBhW01SXoUr9rohMSNSTTPkXmZzAl0euFiVlpk
Fz35jnVktZiDJuZT5kXjLPaRIHuq5oyp8+VWYX/Ew3QKV7Y5i9BEmWHwwaupLceUqYEh5vOc/SlZ
1Nx673AjnngCTtbVg45+NyrDlqlVzPpU9x91gxWSeFuo8jKVKevDPbs1NcNKMNaoPx3Xv/m105/o
CxVaJJH4ZYIu6mBi27otf0ilIgsRkqOEHZ+16pQ7bstdmPVysXU71LTed3TfLvGhNeDSuH+mO+lM
x/8rvL5T8Gw163SEHORmhgXYDM+Hz5Qh3aQu/xwDQjE5HCK0pdhVXcoFTPhbgsjQB5iElMOkjgDc
VILQUBtxv2SjhQvjdvsa8ts8iBhqZHQoJNh+M93qtQrBTMmZog9RmGSEAqNheq/em5xA5vRNnzxb
zJeKdrrgXlvxyFFtvhQME57tQE0K4NP0dAOSEXZRnT53ForG8qqwVMEa7jO1csergl+DmQM3/5Hp
/gN1B/1T3XNd+ejc5QV+n4+Q4VKL0PvLwmCpEKED/B5Z8b+r/ipJbZAzL+46YHx6YKdsWE0Peh69
1eaKriw976OrvVKaiESlVh8amjj5ZdhvTDceaFSkgFI3lkibFoKpR49PDzaYArbqA3mAi5eh5XnG
hpjDvV2zx3Na1Kt8wQ2ayjk3jiGF+aLJyozsRbwNyZeK5Q3x0wyI44qohbBTsPVQ8FcILMLwupzk
dFc8BzvJc59QEJc+FVe454PtbjH9si++YJwuf0/xaYlLxOt+ZRJGeFynpdxUuzMvkcTWRzRMEZyF
jCSdzBjbqSA3JD8uFQ9HQUjA48jFHtuckNWFApNlhT+b/NAqeMlio0YirySAJz20v3qLevGSx88t
xcQ58j39xQFaPROdbN9jFRVRgH42c985EYikaDvwOPZVDuIxoiBhrFlTQI47eUHkippg9NDD3cLn
IGm1i0g6GUHRiothMo9UrupMsjWdQz5y3hc/KsGXFR1o/YcvjlYoWKP3MqoY9/12XB8mxpL5o9nQ
5oOqrfrY+EyPzsRvjaD/gZcfVK535twPztIV6W66fCaOJNZjudBBKM8woanAKHIamyEJGUFOgO1w
9s67XnEhkBOxBY7Lpq61ANh5Fvo7EX3jf/Ec13bJtTz6ru/kn8gPiZtPJEVN7y3qZ1orPeQgn18h
pvEjUOLiCpi90SmRR4MH1dhPmFMxrPy+8Xyi5taJzW0fUYSMCOcinl8pO7/Gpoa7+EErWSauQjBL
glx+aQrGvRpjC6U4MccUVcAm9KjqXB4lOFkoXreZeM5TU84MPpBQfqjATLT4qn9tPlAfYZfFXaLT
N/K9D3P3cCFWBvM+pUIhNoFZnvAkYHzTM2eAiy3lfBcioQ+XM2j/R6ern0jtFmim4Mnm90ce58ly
EPFuFIEMlVmOXLqEd/6YsHKcR6ezb3SZBILNEA2rFeByzZdtuOAUYnk5vKXpFEZdh8+M6nqmVYNF
VJMRjKdACdzsTOr8A/3NUs4A8cvs1eUFBkxSar9i1G6Sq/lkvmv7qM+pfID6ZTXsdUGq0xjEElCN
ghh5zUnPr2fdA0YCchfDLzyjwfQTDooMSj9nqeXRtv5KXTn7tp9FjgXlP21VN6DX9wBC9csm6GKN
EUBJ9htcHdYsBQpXR/tymzcf/Rz7KXyaCgCQpCh1cvl1h//W5DQp9zmDx7HVUh7zum6/6u8YvPTt
S4FGuRmGwu728Zsy0mzW2h43TV9S1dLVSg4jwEskJ2w5q8MhoROM242+YX4pDt2B4WUHM7x5ppA8
ysEhW8+ZkBx+K4HhTozVIXNLRFvqazIAAUjmMQrb1RDmHFl2Wu21EAd8jH+vFuI1Q18G8lIZa0H7
uhaduP2u72DWl9RHay6X8IqarKjJzqTZaqPjaxdhfGrfzkvu3v1v4djVzhz9hZ9wf2oz/s++3TWH
Wsr2kSikB0uepD+QFbV+mpvcJR+gf0S4CIZFrxVDRENHkuvCsUSa1YBxmVD7m80Rq4gKriCcpYRQ
yIb/rkCgqvXs4Hlek739IMnhnHc0mwagThQw0xvYuHDatgl7or24o9sp3XCb0W7IoKUljzAuTfdv
nxLk5W9xegAFvKC/JzMP4bscbuYIQY5s+R+gU1jRNlok6TNyk01OhKqZpBn8rm1K45MZrtmtH3i7
4s0KpuGiRMV4NS0TG7U+aQPkTIp3nPO76eXsixNqCe3bdD/ng0sVWXeEkKwFYuy9f2K19StenO1S
xrGYYtzf6pJLVHlU98oHjpB35D2WWmUqs53ajSIw48UcuQo2cSbWlxWoDPTXR540ZM7zdtOs8PGA
sUBZtW16o1f6+35HMKDP3XOHIDpx8NYvTrUBLvc+myyRTH9kuq4lxuv9eRrdRHq822LZlowj4pzf
A5XxEM+0QYHotgWnmFoTDReA9PpM7SboSGcL7VfvpAPOHGlT+VITO/C2IXE/0VAq6vPnf+n4SD9M
GiNiZ8yVULkSuCaJIajw+gjnWSwiOuC4ZIl4oSjLYgnowChyQYCd9yymmm5qYxSrA2rPEGu7klS/
CvvkCTO7AnMFFdtqk4DgUbXjj3isygbHwHcNsKVIxc+3l+5Dgd4/xoiVinvipfD+N/Cfvi5n7kEX
h8VxrbRkxEWs/1SVZOIRTNPWd/ynrii+x9MzTiXG41MHb1PnDttPe5XBmB0K09GyUQ41xDUATH6U
uGzoROwHhsENzpZoAaUSpcD/XcD96CbiiISFucxEMeIoyFLCy6aBH4UF+l5ykrkdWhcInNMmU2dA
ScfiZT1+I2rGmHWThCRz//ME1l0k1aY+Ee0zFmwe+JbVH6TFC4xx5nIlVOr78HL4uORS9Ultfr6G
43u/Yn1jUtE3iDQgg3hgblL0CRzhkp+T8lL9V8Rcet6TFQQPZZKM29sWhM9oBJdPuHndi9GZCP77
DD6RxMdjMkEZiQ5gaePDvzuSizWZku9C/LMe1gyr3dhAV6Mlq8AHuFx6yIkcGsAirFeFa3/UTcj2
LFVU5RSYY3nB1LMiiJ2+T27nL0eqk3QLuBmM+pjwsHiVLPan3/wMS0wc4oFy5iv3++6d9quBwt/6
zJZD5bCfWHLEzEW71scROIM21vueWqD9dbX0r6YOABfpZhlTTCCKwNE8m0LTXBhCcI0J/OVJ3gd2
rMW+nqo6ap9AXTAnxDr+t6Tn4Vvkr2FTwdeUG9d0RB99Ozyl4YOcZUVw0m3ZGfnRdEPPR08BUJzw
h1IJG5ormIf30fy+JwrD9JNAR2NvdflbORx32SE3UZRexZdDqO8FOwPr3GmvWlYOUmiPdu+VCqia
H0dfvfAZRnhInQty/YuSjGbZziInVq6J/lgfLM6dBInNyPwg0nMPLqHXJugE3ps0aZ6gO9rYzTS8
Qez+RdRa+3lNwVYiZ21wpek1uOdpEfMW2KVW0F/0OfcvyQK5PvjKja4oXJVvGeyO3DlC+yCN9kqU
doN/kC3NHoiTfltVXvClOAEKyOorUm5lk/TBpvd3bD6z8y9hExWNMAXsSdj031ZShTi+HZNPNU7w
PDjTNN41XBlT/3ord4yPEr6k5G3U6eIhKXXB3VIDjVAftMVe0oXM21F1MImwqNamvpuMb7kdqH2h
93LmeeKk3ajrD2h9hl9tM5QnSlMMM0b3yndzZHOQh8X5kux8fkaT9K2WsJQ2vpL0LBTql06fJTik
u5Fx4zIiBQ/nqQI2vO/7+o6BuOGvLqAvy8z0mE8HAnPXX+FihlY0lSMtnHSQ+WhYD9QkrNE7CzmB
v2N8TIXxCAl0yO1+zxGD2bJcNnkAYIryL0Pga+OMQXKK5BhVC1spcOIWZRvGo1eYJt0HKQFX+kgV
uB6wwf/ARg9ZaUfx5+1TXmcf5eA6x1N/SRR1lNEAgl9+Nxem5mmxtdgse6l2XV5qDMmmxAT4snwz
zHbiPRIvsC7VT4+07zfhZRZCnDh7NsXGyO1v0PVOow7gqc3ig0sGGTk91mWJYFpfWpriVDD9/CbV
7Dba8+B3CXZX9l5FUA+kyxazwitM6yAVXhuYsj67PDQRgI8tEMSjl76EkoL6SdKz8DU++fy5Y1kF
iqmMKU+fVyD7jO6qCXRgJdm6ktGdhQmyH2WNp6yVC4QrLagAdTVllBEUpTKB01Yxq842y1gxyt6Q
STGZCuAw+PH6Ej/f9Bo+zAGW5mkFk3PrWeZ1v/8+VOb/JC9xYv1IkWBm3O0y4lal0rephURsVSG5
aOIzVvZWuYny7jerNeX22vevvA1Tol695jj/dMpgf9RdFbWg3ES8LUPS0n0eG7rL8k6E0Dl8Wzkq
wQbVkZr89dT3nqenNoC4VVBczdOzcwNodxC/Ti6cwhIDYo3DKv048/B2O+Wtr8RXbck5/2R6KkPl
+u3RxToEeJYoyNbNKu1YDRpQoBBlr1JMT/QmbQ51CO7zM7E+7T4WFwAyJxG0ji2SxaPzdVXGhg/D
rdpaj5BUkPHsT2joHzp+UE4hp0pBiuvZqwMQW7oNVnstlDwomgeL9JcsxjIHX6uqkcSVTe1enuwv
8SxWA98Sdsv8O9V5/5raPZT8HXt/ukgOefLAycY+pgiDSHmBltRHO55E6V5citijRkk7JW0oKO2v
wgquC0Frvbtaz7DJ0Xv2PR5LtA7uQZuBSChbSj7J+vqYzXZeg6uxklaJ93q5U/5X0VvJxn4/9gSH
4tsIP/+zqXSQgLGj4Or9hWPOmEfgZnuArv4JxbE0NiGxd3L2Qu1YCOUCLuFzn6tKFSOq6Qf1+ZmB
DHGata/cq13fwW2xblwdoaSVOxot3dzRJ+QVQfZpu6XIuQdVkc1/t4IsjYHMQyvvYEZ1HcmC50nb
lt/GUr++ds5uFaNsnjOJ2SYvQQUTRNhi832LE3j1zal2JImFvVXS5pykFRH/UbMYfAcgDSlhW20A
ISBEYKtHGRinN162TrnOPcIrmb+mRdXhtPhteFMJU3IOqhBfWqYkTZNE4LPTdhJpNxc/tU0vWKgZ
KR9gUJdKnD3aqII87r2B+WOFJ3enKyG9RCMCkjrZfcM1K9nk89G7sGCQ4BTtoUeYjvlq4tp4sEMR
Q+ZvXgnVXSc5RPyVi8xweFowlatTstU1KKt+RrwBy8x0Tg6pFzX0nLBH5M0FRlay5CKitavuirSl
A2rFJOY8v+LvjpcPhJ2bpbifqXLH+ypGt5X0ZkocTKfUu8bHU0kAX9ayYLAajbXgSzNKzDkb7RAC
6S5ArALeVZvkYbxvPWQW9XVpdXynb7If+N8MNtQwFGtqYTd3Spc977nNzoNv1iaY8bSDsj8f4yIz
dgjdNVFzJ/wQJMXOc/EO5/n9/cQDPF2rDf5YXjVTRXcA5tQFVGzJi+cpP4MUhbXVviQUCdWEAvc+
wIHaNQHdvjpk+b4ObhJZJQpowANZgWCrO3a0QmBq9Seiaf67SF/6Pua42XIQHIkBK2UNikO4E7Ws
KOdrPXoHHsCxJdvykkvWSeXMev7T4RT0CCXmrw5Zfe2WS9Wyjk61cfAJCVTQD3u8oXsMpgGooKyp
vhgwotqgnwb8b7+F+ow+w3VXAV1yn2tW313Wso2rfkrTlAB9xssg7dawRzRUfvZevCJX4zRaM+l1
UZI9VerMMyEYtn6Y6xOVUVeoei/s4f2TOxv8zTXlp8OJ5gatkXoCX3XKdcGVS8x4uqvCOFh3MPqc
JNRszgMnroH36BRA+9BM73EcNF93QsonX82KraUxIA640T11RguGR0+BO/nBdBTiL5tEVpkO6WB0
wSZqVato/LVr5kSgIaNZ+EQsV2EEqlUGYSqpWRjrP60XRud0d9JZcUcs3vPCukKuIdUFhDSzo1ch
1FTg/RucF4yBuMnOm917sys0EXpOT2Y9O0cLUpCSDeypct3QnkpCIhF+YGN10S25izz3JaRwvsn7
ypN5RlrRxVv6hGUsIKul8LApFikhS4t/Ap/nGk7sGVOyqeBrOgdmALrpRf0Yhmsdg0AIje+h7m3z
uFNk1qht8cvh69zI22smBgIqX1Ki5c1SyOPUjMnuOxWGep47vhXgizo+AakxwuVzMdysHgTPjLzC
9XJSuCXeHc+DMNfeugCgFUtIz7ktu7OZXLJSGihJGwxs84wbnTI4UcM8yvTyZcWtfB1i2YU5jkDJ
s4uZF8hArXNf9lS4s2DC+L+tPoR45H5w0VvfmkF+7IRSveahPGEh8V4ccmU1NieQiaJCAVMj/bI3
HJ0SzxL7k/ELZzVr/hGZvKpWwHesFzoqj7TlQtuh1QOjwiKHpTbSfnHm7N6xSIvu94XxFRz2+ezx
KG4pmvswFElzZewcm3jViycVMhaYxrBc0Ywd6ySWIYl/uS+xNY5zjSWy/gD7oINfkNPhRF1UrsgY
1JtqDMLqrAwU81F9RAgtyiu7zMZmfwY63vybq5hdkzGANOmg2pVj1xlqEoRodRoo1zDqfaQuG2f/
j9k50k7kvtWZMUccUogUmHVm3RojYKKdSusU0ai9rJJgy4BVGsTeRQZ09fbJP6be9H9t/4v+9ZyT
YOYpYUDkscLxX60HNJwD2SOqaeNOmlpuajpSdOuRyy+P+ZECWTVL9JMM8PpG9pdoABYXTq14L3CH
DEkrCYJpLGWOIVTEDcUNGC0rW+4/t85zl9vaCIvpZ8jBRXlX1PupaJzugd/HKL37s+3chx1I18W7
vzofAu4MMudGO3BASawBIfXYBDgYJdCxsODZD35KMALHUG+APJHWndOYMT2e8bOdN/I2khBMJQDF
hv9jc/dXEtI9+QQ6O2eNTH1MWu1WSZ7G/jnfRbx16rlFHfNfbhYzZYJs5fmFK/5eJ3AiEc/PEYqq
sVts2hF4qwniqN17/RtlUg9QbA09mOEudMC8Fcvedj8jdbiNS2EaZeMEq25/RgjQIrR1bPQMupX4
wgaqJBUysOw3YaECklH3NTvpAkPw1lq77JmfD/m0d7P9CHYLrRQcTkoA+Hbx2q+HtEbH0TFfzl3L
Ne6R2F7ykeOH38Ij43SCa96UhMrTtotREaF1TTKGfSUi9VgZEpfIg72y0MOQlh13OV6dsEAbCIB9
DZyw78BdYWRLJbG+8TNQD0dBYMbtxMuLMkxC3GZ0c3DdJH8/cqtB0BSUcFkY1yRODm0v0k9yZxzJ
OORH1kGlhvlii2cGXBOH51diKK26eEe5A96Yzcd6Sa+EBEs75eMzXHy0UR8N8MbOFSxbvcHjZtlx
W4lcAuGjpZapbiTaCiFTcvRQpl+swAczLO9nP68tGxQRDbRYyYMs0b5fD465Q5/uaZ4ZB8ai2B6S
4GmheHYGA+kj4k2bSYhhqXpzLI5ewuXgykkuPGaXlIrZcxclUu1sbVBdiNx+VKgMD8VG5Mir1s++
Mel253JOlnU6tC8/H7XYofGnlASVj7yJnmRe6mEEFEegPrL7FOv85K/GwGvMjvGtcOj46awy8D0j
pHmJAswVpAwixCo4AUe9pVzJsHwc0kHa0ayUD7biQcVBFBCubQrvGrPGMAIffetRVzmHB/ioQWLW
W12gU+yvWlTsTFwElvvZQQA0EEw3cdyjJQoMC0kthZQgoDUMbDq46mXY3ivZMikwyk774qKL3E7l
87DViaSz7Jp+JcqrCUmqFbt1wm7JQOYoH29gjliNCbsxMPlncIcxqSohylEtIuDRQaAyoAS/cH1M
mNi8z34fDeBdTE33/eU01/OOocsoQaS5aIBtfqbAM0MBU4AT89HvD/7fbWPAJlCs0eMWW7AoKnRG
pkXXhx/+9BYNjbzMQgzq9r2PCZKkGaBk5RR9cNBITLUZQIBK9PM+wZgUuxpJ19gbghFT8EEks2CP
u9/1YO0X/qbmSZlZ5sq6axHK+ZwxjtKGXuTPGvsy18VAadaqv2HvrgOHewRZOOc7N0ewFaxCqSX6
gBM4zW0UQtGTuOb5F5KhzJQurMw44NOsESPJQGksm3kBKGy2FWPsiULTCInTs/I7VS7YrkPILXjV
69cYifoepV0bLm1nTnCRFg3MROOVMeYtfm+0Ez3XhKkvDFvLPUvhWIgksYDk9m9yYm/bPvkvIb9h
HupeP6468YvMCaQtgyLqYdm86L/rmauX8lGMQ3QefEZYp17JI2QheIUdlBNcOJ9wbUba4Y+vn3+b
BYf+w0J5ZKMtaTeKNfKffJwBvQcbP/hBlda8ZJxfHiIf4LEa6u8eh6wgIq8XPQnQUb6peNeCPb4x
by2WRmzwgUKv6lsvN3C/FmYTueKeIRU2RsB+6qQZSgj0SPXxJpi/VMXoKtBgDao9odacCH7fSaiP
CFIuIhpHa6gks8So0Y9pQxOJlEq7wxI04nm1VhkXEGpEzBgmctfCs8syORM6HsV/h3plDWbwajKA
cz8K+4I5Xmim+tOMjetFAPviI/CfLkQMJAQWTgX0X0Eql5pfpax6WN8UPmi44xcYCmTciR/HK3zh
OPjbT4KMQ4sDlxMMIJf/qOf/5w08LhIU+QN07l5YAkDLiH5qmjGU6OcnImLgIcrbRTx0WQqgWwxG
x5fNkTewzjJpGoHv0ood6Q9dmxYsGdZVNwXSyXxF+KlyQ5ke4Ybl3OchJGazrOG8jxL4dIKwXZqA
TytGbX+SmQyauabO5bmgmvE98UKAUnb2+SWDfg2/WJJ/m4uxxhzlRY7Ebbb2LstJxJfYk0DQEvPI
44K2fTgnxUbmJWWeF29mmms6wiqM3Uzey6XzEoW264tPwBSl77ot8ccYFbOxDhVKqgV0evawUMtU
n1IyeqRU60SbAxTfSc0uhP01ov5i1LMCojyNtGc4pdvqvsW/WUE1xDyi7Ku+Fz5GtM/PDYhcE5hF
MvhAXJ95WnL8tZcMcKMeQx2wXHGN26cPXrUUJf3PBm/bUFRjXQPAMji4y6zy91gPXbQTwgkLUJQQ
erLqcUCqiMr71mx3h5ngHTq2qsEfbea+KYMUITDvQC1caTeJUizEPDAgNrrd6OhW0Vaiuj2V8k4M
P39fh6oQPhLjTrUMzdc8AGm4hHv8Dt6AQn/hlJcOPVuxNdSXmWoi6khMgF+OuBD4A5qZapr/TfCy
69UJzAPDpZ78oxyAHIP4aMLIK972pPIWhGEPGzPSaegZQex+pST2JbcIAEUinidenxZGGKAIrKQN
9D8fvEPc7S9rqpty7BT+dXPjdBw4hr0cIAd4SSV4YeE29WiTcTAKQ6e4vx1fpGrReKC01bIaiXbu
vZVWuFsV6N4N5WEGgdQX6jrkCArqc+77dSgXKvF9gM+xVU5SY8SlgE95wfNZK0N1cdGbD58RNZo0
IrN/v9y+QZ3TuIWxPQotCl7DU7pK5NvO5ZmzON3eZqHaR7c/zawIijYakk+CaxMsZRQXEcsqQgHd
TlH+ykmQ+r2/0Yiy2auxz8jzt/+JkiQtPofqtcSEwQxytV+d6anuTMlqV0/YUa72yiqYft9Mq/9f
zSGf/otIgP99wDBkVT8ew5t5OFnT+RiZOVONRWjg4L07LxCQGUJgzuJbSw3sjhQzk/+JLKuwSZ/b
P/g1t2PvXLIOOAilUy5TriH2zu6NDy9y2Z5NeGD7tspIZ9EKY6Im/Gwruv+Xp9RIb/8zzQDdgp+4
hckR8+vyz89IUacd8STgyFomFyDmpUz2KneHgClU/TGkhDle4t/m3o60z2psUVLWg0wpkbUidmco
DVm7V5v50aIDDpgeEDhIBXDwL6GsWL0Ao8za0T4zujhFNTYJHF2BgrjTr32zEcvMr3XS3NlCOj9r
nYNHCfd/KxqhgEeh5CphmZUXyGFAxSM6Cg/FoEDB1L1mi/ImaiV3qbR1iZZpMh9Q0jVstiEXSPKs
D3WGBfNJNnR2k2/vl0DXx2B67X/1CovTx/ZX5FkpzKblvqSDBAWfOOKBVQNqih5cRxRfvexBoqHW
rc0xP7E9Ph68PtCyNTpxJHbF9H4AYcf/8bkZO4qr+8yFqs89oh0Tos9ouPoFB5iEn/4En2BNYyNH
AZItv2Gdr9rUEDstlURAWPpxPsgExAojtmUZFYU2TBbbsOovml3FGTYlQ8QWQi9+228QLiIxwElT
ibsYNF/aiWd8RDH5mPj3/3Erlmaonk0guwWfPlmL05SwyRgF2M6JdgJ8Apw5cdAO+diYNRf4opbV
NYDWQUKURN+6QWycWRj2OZbpArrWlSH29t0/sybpt3o4jWcvbifXukbKlhOhiJa6hjzOONHs9K3S
DUUgY9ywBsy43Z38vKaCKFFjhEKFJzatnYr7fM9JEae5NzDWtFTOc8/ACPWwIvt0U/xqn4Ivmc1n
M74uOngrGS8Fyj4TPQIHJxL7Y96lr9IL418LUMZvWDlKpXjg1D3gDAQ3bG/YotatvczVQGcZ0gzW
Qa10uTrOMFpcRSYTK8BTlidwliT5A9MgxJgUwP5ddtrH/V8KtTwxBhkJ9teGSZabOig4cpfc3T3o
/OnSZv8MZcBtWOXUTVo1phhIATE5hifyHqcJ9o31j1AR+zA/TRTaLkLVbUdFnTts33kqtxzJrPtl
vHGENUnwkxqq4H38qmT/QdfdR/u/UKbsdB/6aLNjb+nEantFksUG3BkMPTzUKKP2rJVPGx3JkUul
41gqvfWCK0wZVuDgBq+T8Pujx5tAdKL2PbwHDeyqbECBl7ox66ArqvWtUUXVQum2PISApR5j5lTK
TrV1HUDeddj0L8dcM6IxON8f7zc5077002M9x3KEWOqLcmVbRB9IRRunZ3OVNCgmJj6CsTAGPTG4
nrk9DRou5arvme14IZ3CjgMoIvo3EOQNBI666rbdm8XKk8lvLrhAVav34Cryy0M+lpotX/PzeXCn
tiIRDSogK70u+AaX3J1yyTM3eTiEOQugvlhwJAU2DOD67Q7+SukSnVgFK58gfuMssb9JHeUYAmsY
aE1oH2/HEy+un/kwQ9VqQC5wEswHWCrLW1I0d9dnFOVucisUfC66XxqqZ66vSFZ2Ov4zkz1XLreP
yar0Ae8TDol6gJ02GtnsuFXnb23/Oq8P5DXIvGNTAqG34DQwVoMacT65weY9krI9J2Avs4J+gBJU
KeaO4hSpxk9h4d5pvKvjETuz2/EboaWV2LT8jJQxvSQDJnl4UzdX/2Bcv0zTRmtVwWZDKRRLGYA0
o1qrHf4p59zbKeL6qLDGME+qH2ugE11fRiyuYMDhyzjHapwLw4jNfpC29xznKwrPU1AOhR0Q0Mlh
sgMAAwLzwR63dFowsW0AmeLq9h0DtZGQgaOoGMiH5szC9Wt/PKPVyHDzcS3AC9YpOl8/I2eoGz/Y
lBm2BvLOx2UGcO73qxVOgCDRZoJ15Hi49/SqFh29mNoBqzmyPECAdDhxg78kmXVzcRKNqYxGZgRz
9FMbKn3icl2YyGCnCvG5qgay+UxuAMTcJxrQdGtq9MDofIL5RvfLnYDfaJqk1adU6J844vxmUgRb
/BqW+pxvfY6x+KweZYHnGXBa1DorxQKxjnsU9BLJBExtIB5AOmRZxVaZ63KyUGanIQbXMBOsFaXt
HJG3Jx2pRNvM0I2edGvEFs8m6d0ZHoQykpwf94Pjb5vcI4h6JU2Tnn6EPcMfCrtpHMNawFeuf9eY
SxEpqw3PWcUYj2EjM+n3gIegbw0t9vOVVp9LzrMEABH9lf9S7+RV0sueZxY9GuO9ldmHk1olsRzM
s5xRZ+DYtEhmbgtiyf0tqPbGfZrFc3UcVtspT6lxnc7LjXPdt2dSKrwnr3Gwb1HE2+dupOshsY6H
vSUl2P5OMLV7teZTj2b4yG0QUlIYgL70MfnI6bEY98zwhxNDOsQlCFNArKXkdBpeRgWgG+eUYXMs
NFTf8kVYMBmT0GVG4PTiKvvSIxZ4FRodpg/UfWiiSCOB2ahTw3GhSnPbU+5rbvEVZYYth8RJsBSH
EUPtLgs3IfmpnYnaCcoOh4kQ10kHu/udDqB9O/d6XKJTFQ9LI5Uf9aEALGlT2uRN3GmH10FdXJ9a
x3BsoDNStSim+5llssqJM8pP57bsj+hRGwObkLiMZ+YnGOIk41fR5u6oZOLOjTHXqzkYn3YIvarO
+D2EBw8jfhJ0NPc8LQ3DACHeOpO3dawp+OadgChj6l+vKu5Jv4YXgMuoh6YJ/fnyM70byJDDcdXD
QUHvNDfqtR6eEVcJDRaGP0mYhusS+sCJh9FIEmWNebMMQtl4H17HlisrmU+5ZLQNyuNqM8ZoHebd
eqO37yn4Tu7hmg0S1TXRNkaEaKoU7o83DiIyEBCUqHuS1NB35kdpt5syqnsQa9OBVH2iSWBm/oMI
FzRufu5YViYXChyusMT/KhCwPXK51ixfI2EOJVjrBFfiKQoSUcijFhQ5TY9neuMkTpY0k83nB3g7
qHFBUHNLTOPILJwzNynk5HwivrIxtVmqGWU5uSqHkBdmg5bZov/z6hLo57wD/HnGMh803t/nJpnz
qNhRrNbnIQ/4u3GZe3OnLel8HUyNJVu9tgiVoDQlSXi/l5GV/IsK+ApMm6ofxa1wlMUaGw/7TchQ
DfFgP7r4cF+bVdJgxUaUgoWyCgG1DMRK9Nv6W92tTP5Sz0qv2h7oqRVBdj2yFD7opD7yica9GFkl
rFFGfIDG5BJg+IYxDZiMIHktQIJUewGQDxXBEXIUAlQhq3iOyqSH/gT8xzJl8ufFiZdz0OHNqVlP
E/3QyK0aj+vVwxbJ/EMtnzlIU5QuzIYVBlnuIvRP0gYsvtSYEIMVnbwqN1awGZPwhuzlLyfLY+nb
+Up9iWWAIVwQN7nwD0XXptxRdgf61f7Lk9W8IT3bLRNpDZu038QfQ36/FPpkLnvNYhomcgA+f/nX
ic9t5LTk2xdRPah8BXpTu6SI9NY12WmK3qtmzvwWRbs0k8IfyUkrSjMD/qrXqfpjRF848FCtrjhh
31WlP0wNqb2F7WLGKq+B74r81y5bjSMe3yH6dK/c1r/ClqqoThyiPGX1tW+6mfUSdnQp9MofZqsu
1TUwUsd8JuttimDImg2dLu/jI5wTebfR9Y09nfkM28wt7MkyNRarq6XdhYbDvmBO3wQDbO9kLF1n
8xyOmPJZl0Lhe2CtvdmOXnbAReTUS3GcSrMMEo84yD2Gdb40gpEUaF8A57/d54j7q0DhLLuvwjqw
ne6OFzDnUdJoHq/oOlMlSzSWeWwxUjhexkFuDlY6XvF4+xeuEyfQfOT9PXo1LjBi5vpgA/b6enAi
Lu5itPWgyjFOfvq/bRMdmYpR4p7vB1dI69Y+P1qhGVGxbnNiMUIXcL9It0ANIFj/hVickNzL1a4y
TBYYDwRQQl/N4mGRBfCiporSbtUTktuCs6buPjmxsHpHvAmwCYhLPzf7UQLhly2Cl5SCY+Z+hECE
ts1ZJWQ/GAY8AYT30C5cZztTzTC6WBDr5CRXDSjA/PyckZ+M4X0rb8GJjLy5f3aRI95ThnZSb6IA
LwInSzngqdOzI144KPqaNQMEyjoaZvK7nGRhFQU066HUoKvXJeEIPM/mkqNUt9b/C7w4rWnEsKvq
tQi2GhW4WWsAndkka6efkT7YkDs4MDoWC5Te2BQJGjpAFVxk9aV96CHNSJF3CmKCNnSqdTf56GXw
Z4SaCgmE8ZIZJs6gaScNF9nkhcO6F3HoSxmUt1m3/+YvD24mGkCECuTxiYTqzsYDbO2gvND4P5WK
3vZ56uJVZVU3ajEJT7Acvc+BldudopOBGKJjRI4AMrmZEvZNut67QZ1AtnKSXD6005fEvR/NgNzf
7dSMx3So4xsWjXWKSPM6krVhZ182+0KpHFdUT/g+Bssl7nR0fsCua9HewcVAsucZZZKsbBepJXx0
gi4ag0SEBnUT3BZNaJHvRH8AhzZNMQhv0iREMfTlUv0La4mFaVi4aKKfLTOTf68d12yG6e8/zqgN
crn6zqv1vDaVmXAcxTNIeKHU2YbOyXvNHJIEB6gRqn4K5DNxxS7PscW/jQDl+9m7r+vMvX1YQadW
KqHiwURQm8vXlwPfMuCBoAnEY9w+Tt+x+iUnK3JR9CVi6ksZ2GJ3vIiYJilIuZYCiz2n541hHHPA
MAzmOEOwWYVoKcOT9Adqru/GYlu1S61rgW5l/Qp9f8LHaVxWjE29KdbJdh3JGI8dl7MfX+vc4JGp
6FshcoLDoDD2oUTMgohZoBRYopTbcJQILIvKLKeoGDWxYau8/mbhysq0yZtW4aeotvV6cqkfc4uJ
IfUvvP5SxpZl0gqpIdXjgbqrfIw4q8Om2pQ0wmTebIkDEytj0PgCNWgxtRbVrcnn3wqxK9+HqJ8m
MfrREwk1W2pSgNyWXfVGEsJyUFIXvbX8RL4XFCS4PnU1uRWw8F1z/iwIN3wC0QYELFe7Zdy9eQQY
r5WY5frjxMo0UneBnrWu8cDAGY3kTgMcBiMF1KpxItNcbUMjrqfQavb3vcyqavq35YYOAP4I+Jrz
WzCOyeV45rFDApeJ1/rJNXiKyiSKjYqs8XJ6HHuj7etLt+SOMIYQ6lk4Y1QCHZGj6+58lN3uUSGW
iyj55L8/JzgiOQQquOGVo+F6k1zqSZt4k/jlFUFDrtpLOfkbFLEDxT6pr2QS2URM86R/ixeZU/ma
sMY7KDY4ZjwIwKDciHW6A5PMbkNAf9EjU3ukKCicQqBcsR412imhK4B/+ynPSC5qsHukNcrJAxfT
TFwj6VqsHKStKV8ERvDtF41J38kFhybZpgaTMSTSXRWcKHuWGtwy1oyncha8tbD7OKdaTXEsWM+G
0bZpl8SyeFz77T6II9HXGLH4w03fEwZ0eduip76LatCa/8MQEZkdGsmYF8/MvUkYC3aR1SGqHoSi
Ev7dA2VyLhytiTcE/PVh+mCRQ1tfzMOiFW/aBc+vclx6uc0KApWkjzy163tBQzEXi/cnVt2PKquU
azWphyyPU6ij7gnScCtGro8ZRWbl2XoSwHDAjPIPVmXDQ75PR1HT02i/GD3XGQCU8cGMUEegz2us
20c1EqwSMSGbvax9t0vPTBpxRzy0+JFF/sf6hb5ChAZ2kS27RPogdhbmAplaVfFdEYOFNxS4Df4O
9fwTQeQ6Of9e2HQv8WcI65XefucX4MCKytl47ftQC0K/IkQbhtI3IHcsCbriLmZeTeoOCZFkGSgV
/gyqvfTO2OFIzfg6Oh6q3sUuM2xOkoBy8ROkZ992ZYAjWzSKosZNKlFfHGhJhLtgaGGBnsmL/kPu
J25pHF+MHFcwwGOL23jaZckN/CY/8tPYUDFJD9cEGTKIoEmfAtZn9y2NL86cUj8YPE78hqpABkcV
NP4/Gj7JtXNNrXh0nvWZsmk1WtvLgXIwbOCSo8OwZRSEraN4RjNukeGg7J5ZBIRacAW/QBR11HTZ
lRp/9vGGOoeSRzxFk4sqtID+6lsFUcbvlWuVKZpDTmOJVXH7M3bEYmchw+Mbko4C7WLADqXiz/+S
JT3/x8gxyjLwpMUPSspewDplU9XSUpNGR6YTJtApAE6AGsuNY1j2/t0WiVd5w4akuENFiJpfDnr/
Yb+1JsvH02JBXwPrOxCUngdfSq6A9o/SmZRJxK2fQy+eP+986t1OCoCpjRfKJp0/ebqgz+IbdXmG
XJeOKZJlvcZQsNayradzFEEg1PZnp9iZXMfEnqFjc0dTneUN4lPJ+/BVA0z5glGbvZaiO3puukqT
r2i+RI7drEYbOlwL0WPRNLzLIa7ulABtadi8CIB9SXcrjY7HBWAsLrxVTq+VkwXzOQxpXMgR7xiv
PVJhPuHIeHYFMVLWRNIb2LVpS0ECGcYwSEJuC/qXV0yoL+jN5bGylQCppTL3WyCoAT8TUuzzGzQ2
6OrT9jUMQgB1p9YY7CwQf+G4DY5lRGA+rzJ65car2HJ+bYsoql4lWX7+0H7EfxutvdID8c5bC+3n
Eg3jWedWXMyu8tiqSxRNv4Ktmd7SpMHlx0aZ5KqHdiGbzLj0aR3haXn4mG0adyqZEoiftjZP7iaq
swOmHx76x4pjcVyqRw5aw/aoFW16ArTyVxzRqgd7cgTNjTBUiCKyb3U+Nd9+U8Gwx/2LNnPLeq7G
3k7miIKRCQdhGJWq9WSQ9LTIzOQ80Ylmgjh36e5C5DfrH+TwszSIcKQDEPf4ZzLo/2yivGpxujz6
I+qNLJM+vrZnO+neqGqV1QXOHJy1CpstaEtyF23j9bzfKbt3VE3mVnuB1ADfzlZW4jflJ1Vjl/Vx
zRQzz6oAyjyJ1Sprv6TZvJQp0+x4CbJzCKYH8bbtD0yO8ixdf+e7jJ3doCejaLpyPnkfR7WO/Ux/
ORjiyhDpmDLLpFcMDg2NbQ+N3r/uPTRAc7Vc216WoCIQEbNSWZeS80RoN8w/M5bVKNYj9BrFLubY
gvj85RX5vbxz8yK7Sx+qBxCtVNfHkJM4N1zD2IZorJVieNhFOwRGcNz87EnfhlB3+xilopa3rAin
5vvn3J0bdmCua5O7MAu/Z6CsxxRsfSjRxsDFGMLcSZ1+vM5gE1LSKqTtdD6esL+yVHtgi9C1Q0rs
KPBg+z9BOcmlCIYgwmBCixayuT/18Poe8yI6zVvHyRDNLhOSyGhu4PDx0QmgasrTHSFbb5Dpth6q
xhvVWTJ7yEshoT3B63cGYewJPg1ADFe0kzVzzM3+VFApLqj5XApZlfzJdaxnZmg5XKatbOFnjYzY
3vdCYmrLEPJ241wDKnReokBnmC3Eu9szXlZWoJwaPkzCKxao3FAhKoEpJf/mmoc2s8I3oK3MgKw9
kxcr8c86C5lcmMDtcpYp5CkgxbOj0+YJw52e4xNgCEPT0c339E7H6b2ac5CJOHMbSfoRLGlAbtqn
ZnDt/MwV7Qol7EAbVrRDWbL+UXcrqGAlzK9I9spAZz2iIt4B/JRuWjeJ8zfj8SvGIvtWvIP/g1F+
joS6+ypCidOBMDL+d+axIdYNYmdnRZUMqVO7wo21lyc5wlfz2TvhytATmIysKhCdkc2qcB2Eok4r
/Skwpv50IOROPRzrW6XG2EZf+2V68sOPnea7+DjEck0BB1ZpW6cG8DWR65tYGuxwBZv7nDCwWvHd
AmXJ+F5xqGpqfDfn4NdoVpwGJiEiFjKNp/EqpMjADqY/8PCiVeDRhRJCTw4dtZzo6N0I15Yh+Sn9
3DqqbXE1VvoaBPZRlwZwZGcH0qKMmYBQ/wxEoZBeAuCPYmZ1IVGuy/+O7RNzbeGjrJH9qgpZPC1l
Kn8H7/g9yPbvk45ZueHe7RaS9XytwSQn7lYxU4niTx7NvfeV+RWS/vCfQ+tl7GRYSsS5+P5pgEU8
feRTNLJa3LgDozzPgcVr5g6bIGHW+xJKE4VUJxiT1KcYJw2TvXbzrqe12LhCGv7jsf++dsdkMoPU
1JFBv6x2Kvj/4wYwj4hnsVQlcAoarJnBYLMz0479+Lp2uqkZVxfr1CmD+mAH4qHuzPY7ymnkcCV0
0AxlWJiDwxLYkImHskKZNAFrOkjtHi3AZRm6vIA39QwcmcL27zTfPA+5xOaplpXl7/gxwvzKezAj
lICmUOxLjhJOh0Soe4NTnyBff/EoJfBXO0EGfyTh7MUu/G247qMoJu/eiJVAN3DCltaZjET4pqJF
21Shf9teFhzRu5RdQnY0Wry3ZzyDj6wEWTtl3RUB57PW70nLf+BEQJ62AV3u1UJmfP23vrSd/LYg
/6xepMsbnOieaEIVnqIZQVLtfmm1gSh9ElOFeRYRMk/OJcr/RiDkj8ZK48vbNMqN6tyeBM5l+qv6
YQ5qCRcdpVM/LOOJu5Exwvre/Z70FQZzOE8tclavHkihNl/Z+j8lf4dY8n3SI16/5R2mJkssS3KD
vUjSmAxiBZoXPQqdSwvlQEvrcvWNFCmU9CUvx/N5PBSld8Dt1KCWOZFvdPkCtT4lVmxHHe9CcG0d
Wed8wX6j8lSH8VhW70QF0DpQARBgdtfhzZXZhXELnE+1LZ8j57IhnUAyGrWkV2OrD2WQUq+EG0cI
25tn4KyN0uWU64HdltUeabc1omH0kUjPGlNQW+xoD7CduTjoXTI6t4+OVDImWpVnTLklwQDP9V6x
iOJExaiV2+Sf0eUm9VgA3EcqXOvco68JcTxtn9+1oX1Pwhlqom2dlrpFxtcdkIW0yorsmI5fEwVw
I1hybatlfiMPyyFSt8xBDgIvMYhZKqZ1/u87CyYpxtHH4mMhRTXCOsuL0+lJtONRMIdOTC/FjF/a
re4VvlFMcj3P3hRWqifWJj8AT8vvlQqyLALL9ulRsbq/a8IchcneBufBEwvnzdnAntaHoWMwO4z/
AX8oGP4tf0mcMVFLEpfnMeTW5POylBJWHQl/5uSm2NbZercSEmaX1KyXl6XUsW3GERgmd+r0xpCG
8VeXLag65+C423tu5yd0LK6WC4GoRaxvpG1cd72A3AzFoy6VfgXDO2OQB2pZsag+g8T+6KN9HsiA
lyPP40Hzp+Sl4Ci29byFzeqRLDC+sZXEtJumIKtzVnp//H3HLDqKoP1jCn+mVuGo7T3M4o8PM5dZ
rPLx90f6Y390f7wwSrPm84/7Hc/DCJqMwGI61Ualk98xKvE4JeYobNoXGFJjq2sb9Ko/zANsQ7D3
xcjhufM0iYhwRcdMjIBCWhrFnmd3prwlCef986mUFUcDga7CdqyC5Sn5s02jtBhBIyGhu2GLKQul
AdUqDb1UwAkOHBTw8Ix+v7ORdQoVZ6AMn1zHpCWol7eSUp2R2+A9f+RaEuuELrUaZFFt6Qt2AySh
RTynLvMwp9OqVW+52kW8fxhtw7s/PKd5BBEP94Abmgcv8HvJiESlspDayV6q6/rJc6fpiSeeysCq
+sOcKdn6j/3gN+lmjrtzkKKlKLo/uvRrEsOJ7iHac8LxNbW0sB4vX/KxscI+KYBpYHlKQnsckflR
quHSZFAVR/kBfB0k1aMN59eKOQVJBqd0uicHgBYMS2hu3SyDQplXqNKXAEtbY+K6ElBCsCyLmgLD
nVe5UrJswM4bUS/0UxhFHmfJhl9+LgKd7ihuxaJ+LGsMTndzsQ9VGGE5Ia+YSSCn9ht2u4XN9EIJ
e7oy5V4qh0szOZzF505WT9f5sQSWIjKGjylbVty9IbQvmFHLY7hqCTW75+b+oa0+HAACxZBTEF+M
URkF2f0kfuAOfftXnJ08M7i+KfM3I92+53YUX1a3wFTKZVLgD1tWWKcBgilUpoBqXBm6XWh80NB/
nflHHyKQTXmKYrnKJWi0zqdWeQM5EuCuicc3Yf/Ktk+b5rMZLT6yFJo1gbIiYo8fC48O7Heeh+ld
sqnneTuHM1RMQlYRgemOPNUax9Yqdk5UU4Xe8tbVBLt7/RX3pFO7i0h9F7PrxeiGCbp+dJeS5s+W
ekaVsH6h9xfsWs0y4oxzqAMh08l2jrpTzPRStHPrBgsKjEgSUyyPycYIxncERhekTK193CU9i4u8
7fln14BotvQXyI+lNXmvIkvd79Z1F/44CejEVfk3pJfds6Lo03BDH9mOHZ4DhxXDexQJoj5fwqJp
DfODjhytlf2yf6TUfMvzkAFHNlh6ZCJZUpU8PstW44hB+k5WmEDUThba8jzhawckgVMNTdZY/CKO
vZzDGcgY3e1T6eOiRm5RR/m3+3wp6tgZfDNa7TDi0gg6sNVmCYYnyvWzvVPBvDfymzO1buDbxFdi
9seixgwv6xUWvmpNcZEy1TMELfIDRzvnG3SQfwnbVlCBEOElLLqQZbQ/qZI56V+x87bmFb91OlEt
hWcBnA2ocE4ud3ibC2BVYy72zzxkZ+u3HbkovUJRhj7ARF7euXJZnOz5akMHKa4qDocEcxiidr85
wbn6ym/Z4Tvtpyc3YfUgipBOM73znF3LQvqdWIxxfkYiV5rT46RwZtl72L5PmeOD2bCf/BM/Ud7R
5MiuVaPSc7ppMxIuPU61f51eaw0J7iTg7fTBW+DStSp+fv6B4T1+vdpYS2wuzwUXRX3g6r7D785e
JHXYJKFZ4inHEdW1anPkgCMxSR9oWdcTUq8W3223DfXdp16aX+KAQiEbahjZWH0c0iLkx9OzUw1V
aKoPyc7415qbnIatgCTgUm3fx0OVVqYZeV+WAjarHct6t1ey0JdgeIe8K69O8wJpau9MD3LA/Adg
yM1qYIBWXNc0+2eHQ5pahuvb0KV99AWOn8KPq+hpky1Skk4me22Xv1mwhcHVC0ib1AiGabaFYj29
SXmKaPY9Iw9mpQCn3IbDphA/2AxHWhRxvZC6kpSTMSG9wBSkFQx82CO6CjTLyGMFwsBgHnnnkNb5
sQA9/Tq1z7BxNBpzvnSSNX/Q3izdgUnyUF2POaZ9guz2Ffa4fGKa26jPFq7RKFLJC5Tpy58qrmey
Frg3OItGGPnpE9NvpV6SwWroDdQbntqV64HsGUxY5Ni7V/Vo+yn0oypksZTWRIPttRzX3SGU+P/a
Dpi7p3751YVr8eXIVvXJ/FNzSEVryCnOHstgTTKqJ/H4ShaHyHyTdfi58JajkD7asrmrNS8VgQga
z1F71BMT5jkqNl93YmCySbiEbVdggNV03Bavf7JfYLfbT0hGiSLop4zCXKqqDCSxFR7neFoeK+E5
7FcmAY4OcA1aBhtXTBaKgDUuHPwq5kvbGk8FH0kYeqqONNiW5758Utdubx5TzKTo5Wvep1WYruNg
cisCgFUGpuuPt4JIh/YUd0ZaF6h6j51Gm9zqgZl0/EBWLH5r1DjiM8kWjaKD0Jm6AEAX/+qQ3dMe
bYO9kMVTt6xuqHPOBiRx1Cy/Jx+/nQSR75hrPstLRWoSl5cCWOk4TtQVARm1jnkeC2yfEmS+a7o8
XQtFDjyCvPw9kMREzSJm4teh1wsca227tBD9JvdoQzDIE1SoLKmHXmJPxm2TOYtYV7VJ/wg8bYXN
4MbiRkEUmz3iiQdPgu3AwFtF8mNZ5cMjf0oDp1eN4xZeKzsHn+Gb+Xj60AjxtXnV/UFrbSgtPNGn
UTB1SmAOSp+MZMqr+myisAVxPymCZDuamY8nnXqESZsH5ULA09a4iRddVQ9MGMT13v/ge/3zXfNm
KEojyty3bFuj5ZMi2BnS5pny5cNabla0gXT/QqUjQIRLjDH0EiSrR2P3y+svTxgZXSglg9xAMDrM
JxkNSl3DY60fChO6WfRHJJYfeCkVX00Ux1fAEL2oIcu3jBzsQqLJ2XZP1BQrPwSqJSXhD1hXTe77
KDyupvfh2TgkR4XS62dEEFat1oCfJuO1YO7WgGXTr/FOMlEoAmMxw2+K7wrI+BBFEUFnJTcRMhFJ
t4GajgWIlMiNJ1ygA6gdDOeE110bcaEMz7J/lFpW2II/i9UwoTU+z/E0ojSlgeiMPh7vDYpYYI/Q
2tkMtlmf7LSUEWidn2QKh3/XDXcZp3JE9jopAxLUvQUcHr4u6KlrTej7Qz2xWqEvdb5gmeCRPfnc
0PfLEJOEMDhKCkrY8Ox1zH9yD3Sc+Kx/tDHyRMgztsipDi6JucAgTcczQdk5OLAEgw84hUrm9+Ag
/Y/DdLX9FwpcQbiEdrZZmZrFClTg/O7TCQCQ/oTAuzlYp/ZupUURJFEoCPr7I3/3AOhfVq/DjqAM
1bn2f3OZmOy6Wai68HRG6LvnqW26M1np9UwEBwkU7C7fqIpz68B39Ls/VOwIQVokRsCyZlmNxR4f
AW4pAwlyw10c3FX6SotaEbgqjxA8Ijom3FkaKZ6uxxow2J48Z7sEz3Kp+CrSTsYKj/gJGdU/hhYN
l6/jPjIVsDvfI4KogpXiM5YmdxdBe5bC7gELCI+DOHFEFAT2kSxIk8sst67PkE8ZRk7vCbpPfKXX
wodMko0NHcN/5KmGayvkQo3EqfIHyI5DsIzuGOTT18bYnRmXzxsKLjom2KKlan3bTfuOmrx3elQX
DNrsgiZI62pude4+iSt6lYi21Zy+8FXFjmF/kV4yXOV9gn9m8z0nkS/FpSsAV4uCTnphQR0IJZxn
dwt7AsCLEw5n8YgeQBPHaB2YUzFYF0omk40eRFuRvMqQHomP/URHwm0qaOBP+4MwCy17fGRci+hM
9lhcMxlBdq60WmEaRtLQ+JGLEy3vAxaKM7pm7V9GHaWSucOjzTJoqjXzac6teMV9fzMW5+kSuTgd
gwLezkuUI4luG3oLmk5KGs8PAKv++iwWv/ptcUgP4O8yG0m/U2kECPlIGWkS/D162bLW33lmJtqK
E/XSEj4w4wlCGrFJutoscmgo+QD/oPw+Jph05j8eaY7hHU1utt9qN+b8USxQk//g58jxvhIZ1FDT
rV+QrOuLPTIg8CC9uTu3WYRjP4j3098NFJnxg/zdR83pZqisIA80+zTY2LKc+41/89rKQjXpEPTx
MI4yFZ0s4m97gMAKhyrAbTZ6l+ONNEUquJZ6HTYPvu4Iu7Qf3fXTwctBA8a9lkJurcrU5XVvk7Gv
o/1WuH7Cs9qSpmrtNGHmNs6dtVfcHE8g75pd4SeKkNV6crj8BEShRJ8ntWLDc7edsJ+1sPcEwhNh
WteIKWX50ciEElmLxz/JWZEHSnuH2r6MfAuFx3s8udbauefXppQF1ygomY0J/WDcuMiS558iW3j1
gy66McVhY1KsC+XqiDpSrlaiJ4JN9KYIYAL/ba6EZwxa1WMXLqyoyXGjALqH9vBxPKTUxfeg9OAi
qNiiDEgO02voh46tskvo72DmadIRVOTw0H6fY71ZSUTJv7Q2YW9Vu8vw+IYuooVUhmDppILcaw2C
59tYuQU0NMJf6TJlZLlUAy124bzyHgpGeFAJGsaNN7YFqIbPRXNfwU9I5ALGxfckSOx2HQjC0K/f
KQCkPpdQPD3hwN23haPOL2NCPmCT43JqGNgM9bLDQG/vWqAUC0vfnOXQleTuWG2agg7TfIYrd63m
+uzz6bdpjZYg0kyFY8zlOqD6I/RFmGiQogTGQJY5r6x0XgNIXMvOQUjFf8rcElsPJ8Dz1xbluNP6
lga0pcVtYaLjtREELnG8dnD1csPaFWeoLZXDdV22v4pthIxsF/5PJpSRFIKAIY7T5F70JnmjtJyy
eev2UxKkpmWaSXBKzC9yL/WWOhYwIB3bmQSNCFuNfZ2QjqbFhWtwIKifm8tHGQJKOCwlWVNJQgRu
OUUmMhPsHcMHDI1xceR7e7tpXzIjuxaoRWY5m1/CIaIi4P/EjN9NNIY07Pz+j8Kbds6uSUIMLSFA
itLEwT+Fx8SlN/z0IWamJ+LILjsJ9Iy5KKyHHkw4GmzETx2FXqybt2DtBVuOFcmSunuqJ/TFmfch
M/FAnBTQHgO41+FLxatFm/8iMP003BTuI1yWz1uk0X4XQdzUFp4VkKZK/Eyo/dTVo4Da1FvAE+ZL
sJbj4RpdAkuVwT/X9wTgWUCp8C0c69xCuEHffVkCIjPqcl8gFuzA13bEteitiJ0THAsQrisJ5tWW
Jh027phBbxeYhBJLPNVxE3Pps4fB3MAiWpJ0kXwYsoR9jqtE2vLg5YMKK791dP+OIgPB5G9NDXt0
jk8gR6sj076aLtZL4rcajf8h+PC8UwdPRNlrwOP7iCZeKCPp4HWNkfkTOIa+7E6HRr427zh0rXSO
9ac4tJ4eB1U7hEAWtmZFFhZqeE5AcrKSHy/R/AzTbMiUNBY3Jznk00mta1DvqCPDtNhmQTM1pxJj
hlITj+oNjjWcqvw4ATHi3HLMZWWpq+LyvPmSrcOCd8hO2uPi9BVYW4StDShYWDnAXkrREEYPeJL7
o+6oeiVflThhNiA+bd7XHOYKYLsbUT8AxFj/JLOwWaiRTFe/3aRS0k+9d+/o5whNoJXIYIEuiTs3
k2jfuOhZhFliye82dBRXZrxHraOKsHIiIEJVba8DogtKM6CmTWAGO8xbNzQ7dCcd7JbBVXpG86Ov
2BVclg9VWvVWG0YNIlO0Cl+LPwyncS5B49s1gUzyLeUyPfsMytsiAuApDOVnBTdVeioRJyd9z9r/
fQKKb0vOvwRMG948/BYt8WNnjbEDX6AO7AACNaEhJ5ISdp0QyvAyhwOfA2RK/LugrudJ+ojc9b/e
u+oMy96V5lq/6coy9D7Yc+IJJ2TEmVUdcAHSgVdKRIZqbEntqT+XqCFC3pgLq86LPkej4HcSxDPZ
OnMhOYcDCwaqItn4Dnry1IGZMqFmWrH54+7P4Zu4WDTRoUQx3L9/SGYoO5DOaSCAfT/zNnJKdAnG
wI+jEoV8dOl+nkg3y1gheuHtg0FctgTYKHGkGdkEta0oBe7tYwKn5+pWoxwvR+wA0vT1CWd33eLt
PP61kKerr6zoDY3wL3zbwQgEnje1suHuFnfTCtTJtFlJwQdvytVc0qmSGpYi8e6Rz6SVw3IyAfTH
qocU68+Guogz+RaVHSJEW+K5jlz4E+fTjwm1soL5rdUfv852tnULAG2Kksi00u7pE/EueLAwbNFU
ecEXRJmicgeMpBkxqFMR07OsTiGO2HzOWv8p/stq0F/D7XGeiSaJvtyaF/L1RuWd73EKwRuLH7L0
smMq8wTOWVC3vHIYJslwooMaayLAsFVmUHAsCS9PBqELOnDA7/hoJwbS4p+3D5FCKd8dTLawbwoC
VFQSXrH/fyVh0GY8vRENEWavH6H4f7kAvSQqg+ShnhgCYYnZ6wfZhoVb3qM5xk6Yi2jb1CuawVex
HRgdU91ILrENNvv0OWgLgp8KHa0xtG55NjEKkHvuK+0XQBDOhW97k+5O8kLi1FQHKwtch/YycJ7w
PWWwISX1zaaEoVRqaMXt0tCN7UT7e+XRAuI/TnXbPcCYysHgheFRPgpH3Uoj0nA0GpuPo0ySfv9F
GeQJ/S0UwZEs67jsqCnpauKa0kdFuhItM/FjOfTRxWNRXdtb0Hq7S+DjHT6oTBVucc2NatHnZZoz
c0ycH+b/ImKkmW3NpqRSdjsxM+xp8jai5PwexKN3/aNj1COW215E1bBTsW7o4x8xhsD3I8tVb7q7
iRUXDDLzQII5lNqnhpo2dyDVjifC1T1iauGuRbHBAeoPVQhLOSaeddXfFPMarOa5fM52QKs87XOt
LS5LEbvvBiQfBOscZdOk5ysn0DyqPlxQcifuYNJQkX1FA0gY8/uzZ2sXYQjiJtdVcW7jUpdaQMWc
ev62GnN/D1ctKHK09BsqCKv260uHFRNu2N4qEJRJaEF8ITY3dNUZlyuT4VWGxIZlfSI6lXgtzt2c
3dZAXymfkoSNBn0J1TQYNjunyrpLHJKp6oFghNSulLriYStYUPR6YlZTkKbBDh0b3s7nvLvS+y+m
UDfmBBK3tKEZMf3hwQLiU0OXgXPGOb82nCDDhu6WL2NhVrhmX5nQ5tcBv02CrUN4b/tUBXuRgi+C
WZeQt/YpwzZXzqIl5tKFr64svVp6p63Z3sHeZF5rJg5078FnHFbx5i6SZOv01l2lPTP3QnGg5KXh
PXeDouNWwZ+ninBAQJrP3wOdVho0CUe35yTEIIJ0mec5dq2JWLhiKOFGD/KtgtMkQVmcB9Yvpz8j
3jh5aZbhK3/phaMk6PGmrk4mTYxDR8rMq3w+gRn9QbuD6LvGcQ8SIJ9TwG9XxHkhnoDPfiJf+7ss
ByM+xmU4/ue+ek4Zvj+APPBvrivQG1CeXPz3EJSO4KhEMsWKEscmu0mTtLV9K0ALvaMx9xC4L7h9
mBb9sFxWrR9TixDsJVpeZfN/uNOovjJZLK5yT5gtfnBRhnjpZL0mibgJQ9TkvIAE2KCqRzNLEimA
ooWigQPpTXKYzZM9LHvlefXqeVDM80nP97FaLh+ZF9Aqa/cWzjzvcPDNMkyp6ydGEO4nEXcxuHK+
GhnLLdiGw8tdpRhgMYdFGkeJTtfxI7T1EwGLNrH0NoDWFuL1oWowBSYtpSCsTVg0aHlHe56/AoLC
WTQUQruq/mjdEJsu7QHwmqEo4AlZ0h/+QdrNFsSqRFIEdXt9JOCxlgQElVI6QD0RPTDUqkL4szAE
BzU4lbQtmmelfZO2hENNTsPs36sdW9DsWAgMe8lYDoNK0ltzW7VJTK73nwYE7hj9+baLY4G4kxYY
l+4Vt+UPDOl/Q1gXjQk+o/oOsgQquT9LSrBTFiVCjyQbVWc6A09hoGuDgwqLGrdg5+S2tdrmzmfV
GtkREJr6zkhTm0nJ58zZrGbnoNJMe+vST8cTZUpioCGYo5cc9HGOdxKALKoxJVlQNpAuJOWuf/vl
atDvhSqC0Ep/rbnqxUjoYtVukSB45486UHG3rPZUphj5ofV3yNXgktapz4zOUpRDxIFFax03w0OV
ogDJUbUfq5b/6agJp1tSdnXL7oRrMGHorg1/dtYnubJ4CevxCkLKw1dLcqjYJ1tpUsWz2r1QCpFg
eESmkyPzTbtc5OjbGozW5y2YCoavZ/QS8aN+b01p6PnBBa+Qi9cK7mNPuiJBg4mAM97falWKc0ow
ddNfQdCMpYpM6x1QL1Eze76c8H0iORcC52N+x7VhLfbiG/vg0AwgQORSrSog9HTCOVgKjq5vhLF5
mbVHpIvXvG8f7Tunxj0jm3M9j7BquNblEMN3uGyjA4fls0Q50ABMxjpEI/pTSHIq5ctfgS1v/ZUF
nlumCcZLXpj/+1Jl91Cgz1xKGkbMJ66+0GGL3VoSzWJRIX/lrqDc+O0bxSFBVeH8KBYvuAUWVFu/
iuBNZ6PnzXFyTgaeh3KHvS2KCcqouT9lqGg4K1Dy/sw6SslWGCISVoBNw9XI4ILOZjEY1Xq3XBSr
V3rsxuNrhbPbVj0GMgcDaLvB8eA4/YEjk1Kg8carKAMkE7Nwos0tPy1s6ZXj5WxoerwcyiYLo+89
90O4OERn/egkwbcvHvIdhD82nBvPcR0V/LaNR5q5H14eEurvo5/rCKES6SZU7dckZ6MFhY3Hu//c
GliE/g0p9RlA8El3WR1eFSCfZcBEXvZ86e02cDMboPGyciIMNOaAJpKdBXMk+xcdRy1lAz4ikm2l
+3dLoGEBcF9AZPsXNrySLJAuEp1CvE2Yw1R+vus2WFbzNqM/CDl7TrcAoSloWcVPVW9X9oL0HGZl
1ifXRFWNyNITlEy6K13fne5fTzGX/YWasPl1+oN1bsfDwDcsRmn6WS7pYBiOhNqEI9BdHgijcz81
IX/2EqF1RoXMarRZN2nQtLrvH1D42Dmqmgp+DE7zUq4qzrlMFwTexdldE5vMRQeG9Mxl+qsmnXcm
Y1TvstVfXxEwErD4m/SwxYBGvAs3RPq+ujTXqjoNaYqYHvy7dNL07ar8PK3fLNK2kEf2kMrhX0Hi
C2kIr+7/G6oSHL3eQpxv53yXZpyrRfNcDGGs+OWgwGXoQlDVxFWiDQOR4rwMhO1gEACC+t1Nxc6W
Iye4j6/F4fGCOlKqvxfPI61QWPvtM0dbxhALls++arHq/oC0wyUB1ty8EN2R5mDRipy+KP0Dcyb6
7/2iaThh2nvGkUwz0HLKs2wyYlDp8Yp4RSEd4e8rKq1pPWgTaP+3Zw0DMT+qdrTIY0+zYhEciqBv
I8HWyRDFvAa7tnCP7+KOfEt11qiZK5gRuWCH386/y0TkSLdmpBO4wbg4S5c8bch8/MIWWj8fLTQb
07j+rgRHdiZI4h4K4SnHBsjYoiTl6z2mawla3BmM3dz3p/cekNLsSydFpCCnh8PFa0nCfIlKvdIv
m7704j5SGhw/gFSgbUxGZZEGDZP2vlJvdfrDhbrJiFCvIb0tIyKR+QL7v3Ew65CJU0H6JIiE4ZaY
jcdoXJIzxRj78yfIesLNiBnQjTnQLHQX4LYelA+tiWPiaNOfnEqwH5jmgxxn5rrp8MI8g/KXW/mx
OkUmTl2v929lRMXtbaoKaGDss9IA7lFBVs0b64PUeAVgmlyIm7rnNGOUZ5THcYrYSLGNyUPsWPgH
zAo5ANz6Rqg447lJmnFJcRVE6+XZkQyaKqk+myYeiK3qyDFUhc+Z+sbX8maDYknj82CYfpQlCB6m
yF3NmXkuihpqtd0dpLEyAzV4AXa3qFKqho0t+7w7bz+c7+Kp0lCUpAluGRwDEh449qWuMW1mVEF8
WpFlTuSzbqOy8j5QHuQHmiu2KRWfIbHv8WNncP+pu0SWg8BuHHn/8uVtjgkBQ9vrVXGPV4k6gDn8
z6l84+1Jo1F4v+hjz1slQ3D6KC85kjO3joYvNs5Yj7Zsb5fkcG+qzupiC9zi72ridDMnP39Ac5FR
FAGpCOF98wLIexAy0lXdEwt4cOHe4ouXYfFaOWxspXSJ8s0oAUYljJ5hpmevGxSRys/x8JVp90Dz
ll2QHzdbZfKTu419WWmh1zjCQjvOaTPCRBlj6qwlptsroVH6aT9bkaNXh1ZWdTYk7F+nObphVr4T
WkHZv0/VdmEhRnZOgwJi0TxKF0fO2T5DKT3vSs8cRzb+weZ/fV3R6Nis83WrF5ku8SngNPITSgyA
EhMfWUlgFlAbvH8ilzViz+4Z8zzhaAjHQBJJBd3zItXkgzgM+nzyurioSbX4Z+KePx5/sOf/N13x
7N7oDv3a6kyZvIMjQHravbtO3VOqYoWGnHy0SwAVVk/9ONuQSoJV00jBDUJTR18MVpvvfRldRqe/
7sUyzCa6+X/mujzsL/ptt7HmvgWxJCeOikRtNOXjU4HJmtMrG8dTvuRk6vbGQtsVt0De8Cbo61Cb
lVMl1oQKAO32FO5LongMgZEDphDTttcy+P95lKzBbP84NwaxloZiuQaSR3WMBKYJ4pR0lGT3OXE1
pBJmKPRL7M2U9b4LnCduzJY4GVjB496ChZ1S3uZW1SVefPPVMoBCzLnclz22kAqjTOimdo4EmxBE
jv1fvEjXIHmjIp3sk+BYiqIaoQLgYACkRhaIo9bwax/gAm5BVp3swPShwJHXvnVYQ9gzpyiSR4fR
7Wa0awp2vfLhCFgCh+q4A01pElIxzGP21QVg+8Ehx15nLq3Q25As+Yc8izWHFJnQ/hCBj8+UflNI
N87EAlh8+fOrVKFPUt06JoZjUiWXu0fO6caDkeOMjvLYHpjRW67+teFiBNg7cUEK66B1R5jHQEEc
hLx8b38Jo8o3FsHiqRtV05zZoE+xB+9c1LYWshsCxzdV/Sp4qZ53n9EnV10ZA04wj3tTkN1HIzYu
7OoeciyGGxNqdaLEpKx5y1PcV695gDjf1O0YTaxRWIhY3KdbBEsa1Q7uayAXhtkdeH8ZPMYkbHgj
zHT/k7SCi3j4LGyk47P+dbBRxuFeCEBVBp5RQl/zFIAdDIIShS2nT7QmUW1ROkqwV2obrK/8zqVV
cKmMmVH5u4vgfoPCX7FHmiE5iIYFcSsLO5YezyWrHo7mdbm+ITvSZRR5t5Q6G7RBfQDcnlsvHM9V
PZW2ud1GLGkRiqx7ZBc8VIsEegH4vCuv52ffQgVT8I5e6amxFRsYlOS8uhNgKrEYXl1wsn39Ayjn
GypsUdKYoqKMoRa1u2bCOe0eqc9dAjlUlzX+RPnNmfIzklNF3bfjXiqg9hz6mt3+YqIVEFnENw/a
BnwafI5LUlt0UBWHg6aVTPY4jhM6+7WRoLKPqNyTloSh+LaKvr5MO9SUBIPJhdhCVjx6AP2awY6U
kwIqCrbBHqx1Oa9ZWIVU2wDgzZmWrmjgDiXjemVEkk8SzovJIxZT7D2id3xiT0FnXqH1ZFWOXuc8
fbnSf3+9ecQe8EDMQbq8CqEEwXHbcB9zglRSztvIWZJqaNr9Meob2/ZVovof+7MPUOkb5BXbHaKv
k5R9pBaUKzzPhGy1BqczWLSMNbY/RGw2+Uc7jzwBHI1dI1jsmVAAd2Qom0+oQBjZWg1XZyoch1cV
3xJgBbR+8CV+BcjauStQkTdyva/VQ2kC4BjagHgMxooo6o/E62/ZobZyCVDsdidcvMeysyPm6yUJ
RkP6DC2aQSlt4GZq+MQjmRn6HnMlAUJTIvTKjRT0fYR/V4+05PAGIiOCcb1sLFwP3h37P8s7+Ld7
/7AH19ysRtc9g16gBvqHe2suU+NZHbJ1oYGk0B9rshDKoLEt7jKM9r0amEMYYZm5pav83j3Zr5Ft
j6S0TDhrtGdaBh9JwuR97vU0nex2v1ZzBMUKnh8SlA30lGNdWx7rbqcGIRmpIZljcHox2i7pJhUs
6/uwAiT+x3l0EJvGhjUVkKcoNEPDtAg0esMMtoYpktu1nRrtXOSpF39bNoh4z+62HAgx9+C9P9xV
OArCdIXnqbIdWL8kXUOe/8KDqu0a5zO9bsbCrNbHTlbBUfNdAvdCCAVwMVaIeYcpiXCGKzReAqOy
X2VZgE4ewHNphDdRt5f3sgpMDcRV4cjjhHHhkpthT9uiEoJjJhdxfrYkUecfe2VyMCKi6QqXVhMR
l9+a0EySEjJvq+FbrksiC/GN4x3DjZa5szzChpf9s+J07fQALgB6gWdkaoSdZvu0b6mfneB9n5FZ
HeD60qeKOYfI4MrHCztvfsM72gLrDO5pW/ops53EVBz5Wd6pKYaSMP+Yro30IbcW7VF/AoOyjy/R
O+3cwm89z845eBNAY70J2rSdu1NZ0c3/KufvzX9ZStSi42m2GPhBzdXhotonISuis4QyH4oWOhVx
mUyfJo5J6lzMp0NfeRBwiYNv7Vt8xuAVYwTjHx33iuVyLtNen02u4bU8Y+Wgcm29J586ZPC6FeAZ
5m7y36EyyDl1E2Put+FIYN6gtCOHAs3HGcJN+KA+Pp71zq7elDJqwLf7BTGZpEYCI9w5/WBKaKBB
psMW72d4cs+Exgt2SJW3/m8km4vE88g0j+CmdD0Ym/GuCd+G/RyEjFrmkOGBvs6HXZjor8QpkfXk
YtdXi7130zHHs8ADOcOgb5sPGLtgsOqMfET99oeViXNA1L5xTEEUyS0lBYf4PYHA7QFrp8bDBMXZ
5ieCIu2tnJsmnKkLydpJjjzjlviWfpEyijrzbtE3+DKvjkA74gtrnoqYbSe2LxAY0V5dEBXGkJ0H
NYbRgpT9CmQwInDx2/SrAwKaRrNXHMrI9043buR/uJGoi9xeCYAe55qzINIjRNe9oMZoQ54sSRGo
AjQAlIlousmSFSK/OweJlvw/kQOGe3xKJ7DmfRJQitq7bylLLDRuDETp7f2rjfsjT04BtPppSzy7
fpyjKX3QjBuhgD8j23SE30o2DOhbhrJhz93eOPCj+edJGHgW4fNdtFYhtTsXzkZ/19CsESyL2xMO
QlxNpZYC32K4tG+eQUFClzPYc0aT/LhEWohwxufLcAkl9e+xiGeKzIQeCWAVJGDMcK5igfTZ8k1Z
WHAGPWI5ceCBRVQSVC1yRaUpTFMdjPCCCpKUgIZCxhm8IpMzChC8uNN5h2S9Gh3JUIxERylBl5M2
/aUsFTt2l7nXWFqdLS5okCmJkDIANt5pzXk6XZagaObT8T/a6O0Q0hOhJ5MOily+Sp2e3dFpp8/x
ONv8Z154R1FDJ3g7cZOnLfgqNFuqGF1DG4A8ghfU0ZDsThIVNpvO0tYL1+RHGaOwNW/TpFysDwzE
3HQjgnNScZxqIXueNjJtrO0el8ATut/PxnDodMU3ogooRLreM0q+ITvuSccR968zjoHXcyyj2MXT
g4+MdW4/deC694MINEFXckYFW6HaJHfHgXfNGGVVbQBpzj4GKuzrRXgkPk2FHUBv4jkpJ+jitXc+
LDCNiwweOr1T1oWvtiFM5e4RNAnr9ndJfmvZ3b4k4cYSPwOHWOwVrOavMo8JfXg+XEYUYx/CWEKE
94fnfeK0QhHY0anVuLg7hi3fCE15AYN92RDjoL02xxxVG0npPnfAcU3/R0c+70VxV+V6utknsxse
eUbh8afv8eS0tFSxiGUAhKTesE1DN6vE3rmd11rIJIrT1x3EPxmfWfwn7LlNMFWZh8k7kzuGZRZV
DlhhA36JxaFTXcnvyZQdaVTXVoJRV6Libsl1IAZm1p22neRv4MynTj66IR3bN+lUjTAnZc6lLsWZ
NFJyyNr+vPEcHK/KD/YYnz1K5EKjPKpxlFl4LI6Z5GQi0t8EgVezaL8fru/pO/T46TI4ZYoVAHfq
8ArgIJyMugpKmlrYO0KcZZkbyXWLVsGcvEkhgXjLyo6l1mOzveWu7bpR33iX8AnKX1jUB8Tskckv
38Bxg2XkkiUaZgq8MFk/ozKgojdlz0+pQ6QSGRpvO+kDKKvuSpFb8rqWtL9gujktKuQuXjog+Y7z
l2zC9VGO5EE3zaxNk+zKtSis8XEuWm4dL8lwf8JBcwopcQ5jFT3JsUHP6FarlIMtoECpA2oa2Rsj
TyfWNqKg4K8KYULq4ZhA032K2VNLk1nXsZGT3aj8nouK0lXLvFa0rLudwpvn3yWO1MrLs5druoAk
XAJnQ2pJohuDp7YoAFFUOEsRiCBl7+eeta4DUz4kj8EDtiieQS//vQIGkIUQ6E0QF4t3A/J4XO4S
CFOg9QVYpT5TLCq2tFG52nkHDN4CzByeVEzA/OdPDclvzRMS1dU2koDQ4IBtO8opRKaYhcUrSMUg
YbeqxAsVH06nOodjonj2VeM5xlvU/e5H+HzxzJMpANTFAxU6lP/51PbPDvmNvIpgny/38YZ5id/O
Dap02zm5uAAWdd6/m5NGhoYDrHBkO4nBliR5T8+anx4srTkr9QxB8yM0t1gZvbBmextSxiH2RApX
99dE9JjoQ2JWYQDq9MJP85xyuzzo1iTRfixp6zuFuMZrv6huLqcndDePTONg18hZH6HjoalDHIg5
AOKeInvmbNGZRraYoll7PHlHOdZbaRXjl34+V3mEY2RCl9py6O73Gpd40MEDGW0aVH+Cn70SbgVx
eP37DoumahpEdwuD3XmxBJDuh0pJzmz9oWRU7TvrrS8crovgpnX3rcxaieBbtj2vwu3Q48gBfdY3
aZbmNBdUUx1I4q41u9ETu78k2A7sW9yHO559/H/fysMs0eM8KRuh0gaPi7lm3FrFvBmHTFc3mWXN
WYmQ26NkdVdSqbyp2Z7kXlJf3+N/8oxd6OuDDmvh3cJM6oRa+623bm+7w+pZYqJBdOoByFQ2Y5n/
94R61wX2QQkKMZFDOf037+aTFmH1/dtsfOOcJ/j/KGFen1UGBVKkZ0CdKWTuXJ5NVtMFY7vxo6sj
hN1Mhv5mOIDjZYemj1hdo6AWqVm16d7/BEsTF7ciplEWiJab5stS9KP40RSB95BBfUD6v15g6t2r
oMl64THeihp2Lpw+A/PbvpHiyPQvQpDINwYYebE+l7OvvwsXL65c9d8ZvcTb3GYqaC6NPD9pXy3z
IHRZyOyRTJKsgaoNJDr1T6Pmgl3+rzyvTpPxhdm7kudvtKRHZWWOLHxj5ynwps2Q6fqmG6TquXUX
sFzeQqI+FcnzT2UJLB4tIpUFDyPsZbwkjAJsHI2p4c4rCWPIrlAyHMB1yjW/9LPAXtsWfn9MNRBe
JUCVzDK19CvA03d8LMAl+446PoVj62ILL2rDsXCfXwNHdPJXTxdICPPLDhkg8lVB4z+0b8iUhMtk
Nl3/ZMcX43cKPLVFwVJDV2yQ2nhdFa8TQyZsW932Bw9feCKsguSOfxL8+5c4d1uEzagq9KYZXEfW
Uu3tQhmTY9DXDh93SIkcxw7IGHNnCObvbICJH4RhJcgO2zqfe/ey/ni6ra+rGf6s/Vyv3cY+1GC3
EUmHML+UHuod1OyjtdCkj114Ic/6IJbuBZ1MzICi65EuDi/zMQWVDHmXr3nldqEsQ5Sy8ESg01kN
ipoZeQg92CiRwNJ1VvC5BOX4eq6AJoeZg/v8NjQ9oOOHQp/t1r5ut5GqYWesPeVV1Je9GsKUat2i
HC83j1d9GAGCJhOCQHnbsl3Z0yScKxLWSwSeqHxN/5cF9788V6iuDv3WNq1BgwCsmp/b3BpLX6Ul
m6Ggr7wU2C17Cj39vHPJZ8eLP+XTJK9Q/qZ86Vp7Q2ny1e1oouK2Yu7VdEBIj0V5JFLNmVZBk/KT
qOkbLx/jQUD6UMuMk8tpbRZe/NW2nk/M/VfimbGMH987lO7F9irkzvUtxRVoeC3aAsiK1DciSOZn
mf4XyfyY4CkoqPSA9KH7YL4AcmAt4SCMAh805lIJgELmT0Ot9EM6LbwqOczodgvUK+M7y+xw1B1B
2JL2ad/U8ImUimGXCH86E/MLSsduyfCazwado0E+RS62Eeaa6cPT8V3pF3T5JcaGGPJM563Tf947
n3iuDK9sEDGUP9KOBYpj5p6NYGU2Q3JirJ5CLJycS87VgxitEUcKoivv/aW3kLpfTPzSyEOv3Ri2
LBmkXZu4nwljSgArtM0cj/ildGyOz0dNCnNosxxVhc1stiLjNW8d1Fte5eooQvXeqGPoJaG21j08
yfoH1y3iP8zxKl+zhjMjlqbl9crUYmP2S+GbCFX5x7kn51yzPPGtuxV9Dzuhj101/8jZy3UHHm0d
cnz1Zmbc6P5ecEghXKcQ7eXGXP+N2+zEgsZA+YQwkGUO9dI5BOivGgYtC9ro6GHhzPIgugvVccVD
fMZ/aHkW86XeqWxuXpKAT8n+HU50TJ0ufDvAtkl7dTk7L/UUQPcUB3dB6BKUespUunyQ6BEbT4L5
3LKjXVuQP75KmqrpAZ6kGACagZ6oH0MeTLZMNwdv1xs6K9y+jodhYkZRf9cdO80fnZjJ+MZ4B77r
GYsAJjZP9b9gum/RgErpH1UERc9kRx6wLtqEwMfziixhoujFR9L3YMm33gonhr631qcCobDrqT71
m323n+wcPvnOOt3RHMZNJcCUYjG7dt8QMvgm8jhfpjaglbZIqJ8ve8KFCOMrIrLqLr6o/D63XyvF
cf9Dk+hIrcCJCHOjpGpBInHo8mOyA5hYjAJ+GwModfgeY3EHJq116w+lcKaJKRucaUkwF+/B9Zmf
tLIp31TGbJcYwkQosZwVnONhR7Zi5IIbGB9lgQemuF3kilVJMFKlJKF22KjCSBmg37M82kCmUPMM
YhpfQE9Q4N5Ja2TuOwWMpuo3215UMORnk0+z67c/BVYgxszfPcxYdNLRrmj5u77U9C9K+OIYOkRk
GLciPI1IOwP78Exd18oRmQSZmznd/JXucQFCBLqrHQUnXsWSKl6yHxEV/roFV6/dfIK+cUG8dfaw
i3hSVaeYPKKkiNFNRfimC0j1kIo+amRrl/klomKCzGmMfAYFDZS56JV147GDeF5qi4TWdD7/BefU
jl8tzZJe4baBz0mv0gNqeW3AsDU2AXQmGSIKmHn3mglJfMIDTSzwjg2ZFZg8k7P+EFIaNmPx0D5B
f+rJZdsUhkFwlDRAIlKLTwZ2PcoPEnd1Ij8pDMijs8OeLzcOVxryCOkY8qjfHjKV2RlOgGaXwNkZ
LuaTL7u27kCW8fq/5wGUbxZ/8oPSfn4F3G7ElruIByyQRET63vn5L5r6uVOpDzH+K9Vr//0rYhbO
Na70MZIIoh0cVTHwkwif3A3JXObqbECD/2pYr0NUVvjUFQHR30Ab4dxlLHD3GcO887xc0F8AqWDr
szYWFca94AAuy4i3m+cdq3ftA3PeVdgU3QJCPKvLdzNaPbjYX3tmSr6R+l/4gBWu3YyI2yuQ562w
zB9veq2+XlH8jHZDLlG6wXSGneKyn2ldRz20cPs+Qj9YKgqD54ebtVpKbnte4s9D/UEjw4XUooyV
1iRV79O/y/4Y+kjH4TqQWK7WuZdNUmVNDm3ay1kuH2e50L7eUX+n9aHPhvxxoar+mFYrrt3X5O+J
fzK6EEjApCFGTdOU1fl4gd//GtDmOeanuNbcUwggMX1UX/JocLDd8V1l8H00WAbB96jMSxxkgS+Y
DMZgvHKX4570Ezjhl8F9M7/4v1Q9ro4jr/2saQ6ks9VStY62zmsQbT45weBSDXuQi5nuK2JP4KLV
k1mOLtPA6LAjLi5iT2lrW0gn2FxHuovzuqLtxtBO396dLxAvYhZoB7mnh4mMJz9eC+7c51zeW6IW
Y0292uwe0W0I6PbtidLcIg3GputYy/x7zjXQc1hqvjZsodgG6c9VjJcR2GtAg/0UJbGJ1TdgCYJ0
8hDrJTBK3zaQgSdNzfyCybvGTj1OamooqlOki2FWqNIbb0X8hiCwh0RfGuf4nx0n+Uh/4IFDePro
+jBvoTtLUeEJa99D7G4oIXOcI+F5ztvamNO3+ROCTWG9NuYkkOFzqTq8kDGuRI6cpOlp5LL03PHS
tGVQOo8zphZRwEA5VKk8RbbV/jqNxOfhLImZe+NEA/GkfGaCWfxVwrK34dik8xRYu/VnldrQbhiX
kA72CmylDyUsLLOsUGvv4lRXa7zO4V3zuwFHcKJLFJpLUXyQ9g/rzPsKoohJzsS9mtw7SOIpex8B
4HdO3LVpN9MbGEDmhJ/I0OB+KGEj4hUP6X85/i5u65ImZq44Y9D4yTkibvFTTM7nP1EQqG2BzdnS
6CpoI3KjIxAq81mT1G/MIIl46KcDUDPfZ/cXBZ1pkBd6CxZnc4Y3/LddhckYwFnwMQVpNZ5W2aDw
KZ9vqywJK4928CYPbtkwn61VeVxfmaaHlPqpzP0QgPfbp9C8jp2fa27rkKUa5DJyQNxohGk4YxWN
86OtRhJsk+eB2SNW500jMPOjulAhHr6so2Hrusr1d435J5sw3GHSTclwuXJfNX4F64KLPse4KAUo
yPgbcTEdj4Z8ftC8NjhCr3gfKmvNUna9ZgrGpsri/SHFoUIP7Qm412KelE6vnGcI5po7s6BGfsMu
w4ltA/1kolWZQrkVcyZvgJf4h72YsktQHvgPM/vhLWcoo+yiCP4GVdv3l+5RSNJN1BI5LAH4/J4y
x3aImK5vQZY+5GGajGc8ObTbl5Zbn+WaQcP6+ofYGJwQ/Ueo9imZTwtrTAw8t5XSgklyLFwkxa7j
1OlGt+8c1rYhqey/miDgYvxyrn/J7OcJWPKJyJDEljYVzV0vGSequHgbMTCIDWtxuywrYNf6G0nx
TB5sY8PxeLlYg+3K1tTJDOb/iQDhjtsTDHQNCyzvxted68XBlUb/kQHu9ZKXbYmtVMNIRdesFkXr
f8Qffy08W8n4P3BcBcYLFIG6pjvkL1kPEM/Azs3Oh+k+Rolh1zs9ePTamS59O7+wyIntAWJhTHvu
ilVy8+wv59o/BEiJfSZSu34ZKIAw+wXdkap0KarrY5sXrHVIPrfej0PbHawGXrP3DyLZzmBcK5ts
oohPonv+OxxcygCREc4cazAhWSRg/umKkNkOtIqkG4oBM8GeiDpSEfSCELR9sR/ja/yZmvcn4wIb
vKZ1p+UPcGJdHPlbV8LHXm+oeXPJ4DawgpFKIbpbv8ByelYMuOM3GKaKVOcRHuNoIKxblodMhGCS
7Ajn7hUcxHrDLTYYV+3Qy+9tXajcgvzDdeFAAv1qBJSLI4wA3sozar3YPpMbUDtf2hAUNmOzSELo
B6ThIvnTG7ww5XsMBMADjhlhbmDL61cBEOhYFJolRJpWzu6PPuNu3j+98seX9MOa+U7DhUu7Tr9h
G7c2wtKfUwr77M28hHojxHLgT2Hq8zzqYCrfT0cYVEfRr5R9hQCx1w071LkAK122orCKpWwtnJY9
CDCi5tp2kiwlaB5fQzF9A4IKLFnRjhy3iK3cs0Ot7k7XSqxbLCGZ3TDXn7tVxBiDBfI0rU3ocKYh
qaVBkqdHkOvE9ebwz9nde5+dsCsgV7655jJ7Fj421cL02MwZ28cX3mzoz1e0gcBp2Y+aZI+wSo7a
4ItfDqJJy03RaT5EPOsPjmdzdadi4QZLcQ5RhBMfwuvq4JLqmMgDsu95yV2XTHbnc5+I1b1qR3PG
LtuyQRWxRDeVPaDXqIdeiyLIClITT1mZoAil78nMwjMN7WrzBr0EKiuV4kSYfU8mSeiMsnzkbG4s
8i/OiMXaxpOwh+PJmIqclxVrrttI+8dadxNbtK6b8pKR46k9gkfqvS6cjlLRM13HCWt1KmcwbMlx
Ytj7x8HIc75D7vmMa1mXlc5xqFFQKnquLiwaiR02MSzsQEjXMaP3Mx3mnYIJgO47fl2ZtBh8HIUZ
fzhfaun07pQOfmXGEZJz3wmnHz//St9chTspLwWH/qd84KE44bwh5qLsBKxUNcUqLLhoNyZwcO1F
tVfnoMAq4rpxOH+e9EmYM+1mRfKsSEwbXdvtptPAttG6oyrAy32dED/dS+/55vbBK+I96E1MTJ8/
b1TofhVMTxOWOXAqdR5f43rrIsDnBK/3P+StRqP7yyc7gUSMRmoYfcHCIHV9wbQNE4uQ3X+l7qiG
z0iCQTLpkFd5rJH332TDMu2yLZMq6IdxlL5hLn4CpOk3sFLmCP9CHpAZGbfcy+A/pNQS7dt4NKPh
fwbHXoawSIcqrbQn/uSWMka5/UGqlX+KSTRFgG7v6iwdfWMHg761X5+ZCnCTU0rMs7U2DKHnN2sk
viJIU4bTQ7RDN2bku+HVLJ4QOcJ2DjBYyfwr7dKxycquCg6Ps55L1/zWSOda+KfSuFp9wIMIVohe
Vc/gc3NgFgL23VB5jqTNnE1eaDmthz6WqWh+TG3aIjXut2uCr7PMlCyPLx83588Vj0Qn9DliMCHv
5WK95yAQnebbrXqWa6GPA2OYgMd4mhFpO+1sE6592rcNsWilwEJ6+Xfp9pBRqsmjT4ja2+JsgtUO
Q+YJdIlOXPcPBWCsXUJ7tmVwpyYWn0Lk4vySp4gRNyWrURc0bQNiTbKv4BD1WmdIvfKzqrbn6sp+
Y4Yh8JKxkfy1qM9DKWvNbw9DO6BYDD0s1kA+eczUAO99v/vOYqP9Js2fbB+bJDpa8Bo2DP1298MT
xfRdOhSpbB/U1PQJBcyCBU9LOE9PKpSpLnNwttSfcFbG9f7pJmX/MWesKkf/IOaEQ3Hud1TyevnT
OHeM1yVFfz+Iw6i46/zni8M9u3fMcSNt89PO0GP3s5O6G1GlBnDbi0VzthFIk9W/moJugq0yMKAc
18PgaRyPFSfmKp0SpBwWoCsoM3qgGmMxWhqunJmiu3wlaGFSTfloOjGPiKgA8ZLhJe6tUTnRhTC9
O1yk9563rZV57jErhhD3gV/MF7e70s1hkhUO5rrYUd00BXGfj1/B3nwE/6owcaJwvVrA/KcZ3Ek7
ZI7eZp8K5UnHG5qHEpD6maHSi6tzpaEhhlIzFNf3PViDcczT4QUxu82ahbg8ymy3w6jCHh5rdvC6
pcgSkGGf5080nedR8ZAiPK8URKoNxi/JK0gEv2i4BzhfD5ojJIgM2vSPZGmp713HWfR2GOB/21d3
8LjkkQmf9eAvdIfa4GxeKTiWdZtIH+zGeXl1wZMSU1giTt3znVPhD/9KlmqhFXLEecSHXzmC5PgO
1FBbjzYBRjiRkKSFYXjRf/6HAouq6RevUEKXpsjQ7xuXmTvURBbdmCQIyA3zUxw+qhbEbql5FphK
89SIrcR0G1M1vhIT1oEWSezjYyjVnrAonca5K0tTCo8UkWPuSaGBxHfOQHcnr5/lnRRl3zk4fODQ
RVWruw+YTdjyVMBqI7h6gjG85RXblN7QiwLON5OAQ2rv+CALPAqLBkNpPv3FUTHlYS3fhILF3Slg
8/6ThXpYtClIS5gS9iwDJDAMGS5WmQx5f6Yq3hYtlqHQFiSQyAjkwR0WFaY/RkYRSI4t8hoXdYs9
iQU1wxfQRvFgT3wbWZKVlJ298TpXFQpdLEVqaH2sH2DnSvCXYvqPkVTlp8KZub9Eup8PmULXPgk/
8a9kECW+dsVyapPC/zbXEwPugrWouu+RWqAQY6hpQ0b3BY6aMD4K8XOYLrJUAJcxlHvkuyDaVren
eQz+o/bsS8WyRh7CTbrrB3zxYgl0c+wW7SCh5gQ8uwf+Jl5KqzQgZjGzdRjg29vulAX4p2USJB7Z
SV6cnIfBpsZBJKSVF0WofIBUtE/SGsiNRDTR+0tmotN48ZiC9FSLAc3dap2lImJ5qp5/f3WJJPu8
FN5OR619eOKN7bUDwCnDABLueZH3HvK1Nqgi1rimQXKHJPhS+toXMRkASsvnkCqjvWABQDLjM2Y3
0PpCDbxQzGlX2YDnDJ3U0joHFxdVk4UPer8nKzUY9JfICWLrOKIXqjY1X/Sbp9rCMg/i96F77+m4
ZjGcnUSt3rnOOrtuEBqYV5T4pDHbsmaeedxX8CDtxlqDQcN5jON8OOMvR+4YDsxSafLziG+G+uJ2
BA+RbY1JbtGQ7Zo0GlEqdBGwCWPwFCVO2QVbIdwYUb4PERgZg2hBupi7GWjbQr7Xmrdm3dlKR1fn
Dh4MQgMRHEn8F6CEpjCDZ5g0fcvPEazpeS12CwGzOqGQtdbIgBu1fER+57frm3i+4AvQC4fHD7d7
foIHGTkRv32nNlPDO3Vso3XDRg0hTJxQl4zhhZ0LcCqWhhIihpHO/kaMJAzY1ui2YeLkCvehl181
JD+EVWcDO48ab081eDF+CXNkV0opKWVe90LA4G2DM/1pkCkAtoETs9Olj77EbDmaJsYZ3wKFLHF1
obzynPow7NWmndS1tGxOBbWHoWF7Z3MTrBbap52hTApTdmYK/FdVJcM/XnrnW633cCnuxc4wyNn1
nbaYfQ1el45hFbO9XXZcIdLWbJC9EBKD/BbeG4AI/oh+02bZCJSBC/tsxKhV4pUX/8Dk1Ez7NpWS
Zp3IDn9NrcVXLlwwRKE8CyEsE1dm4O9ryuNVUIOcxnFpE4k1MVzQm+zVVqa+/U6fSrPJPDJBNTTM
oYhak7Fox15AUp1aq5z/KrtFNqDlh8HmBSmJqE2Yc6Zo//dhySRa55ES283fdzentiNLCkC0H/5U
XGUNBMN42179ltPwZth1C6mHy666V7YbzfH8EJGPLDWXg+AArgCXLUZwBQfrOQcqg/INh6UNhYEv
He0YFqOH1bZYBaKoPXK6wAgBhZJxOEhCUYWvnJ+SAuLOKmPh7Bp7ZjCUvHV3vG3MCGaX9ZxoNQQH
EjhZG8+Ju6hQX+I8XmeSdquyEWWL6L7yPcAQkNyPG1nYJ1imV7uoY/XrZ05MXYdu0+pj7vZi96Kh
niFB4MMs2Eo7zgcJAqIE6MB37VB0/dxms0pB1PAOYbJaNpejIz3wRLBmXfxof8nIExnxSDo6C71F
YipbqEU2z8cPENxd5Kd/tq7FxlK5b8pqEUdHVs2xljtCBGDSNhWfjZJD+GDyZPr/ec9roUyuOI/U
v/IGBheZ36ZDYnrujeSKfAojeaw7GlFEGmcotKeQiKvRG/dSU/SwmgQId46ojTAj//wAq41z2pvX
QAlvgJZVRv6RZFAdcGG2AqDceyVUk0GnnBdXD+Ihr4g3wn4jYZHagW0vcFPOcIbGc9VNsH1U7y8G
CT76lHlFQzSdAOltZunKOqJ9ndx+iLV1Icv/JsHhCKyiseqBrMLjd6BJJhfcJ/U9ep8HEiQHR8ag
QSSSULPXACuf65JQ7JNaxx6uXbotuS/rw0wZ1QQ6qDunMZllI5yLWD4O6Ztvi9xcZ+M2LrDNI3YQ
IhoKbOwSoDVhY0eO1Zxp6vGCiVi+P6yyduguUu+vFLH0qWvup1zl+4n2Hd5qn7rcjrxKQFH5xHYz
7H3+hckAQ3YO79a1RcHFZM4j+UZPV0DNzqNS0u36jO86z+SfFuoKfWTVo5nkUA0B3lCJs9wuH9OG
izH0cc+Jz6w16wtZx1jUPf3IVxYjqRHehCHFt0kRo4utXflMyChlRFseuDncQO4YvG17kiaO2wZ7
Rjw/8uaSTHKbvd6Dk+jNUIEGm4nTSlUUdFT+VbEXXcoTYJaBkOlXopfEnHmjFeUYPj/JVeIjGIi8
jxWsaXPmcGQX/FmTAl0g44hspFxgcPamyjiUppRxfSqPcJS7INtjy/192Q8iZJPuiR8aLsBXZQR/
dgwcpoCEwuRb91x2qdr0thM/kAUpDQVWliMS5+AU5TqkiZrF1028RLSvx47Ag2ZSPzGxHB/iXCPI
WWXgf/lDQOQfocB/PeR4EYkTg5pnno3RXGqIsKaSqX8osjNbu5ixPmY5g8SJIQpS7TR4KNemf9Zd
k2v5umhb5YFX3WymAmIy/IPKC+bSs+Y6FzuUI3SQ4gRkwTwaS9XDws0hhAczKnFGi3LXOoNocPT5
8Vt22rCgEg378T9MywzVw+sBHybpJ932Gm2LGvhOFnaWpEROVXm/xIVuVrc+K1nHS6THsDkSAxQO
lZufuZnasyQbzaItOmgsRD0B62qV6QDZjMm8PfQQ+UjiWs2b1QI0Kq0asbhObZlqvUsbRtFH3iuA
3Oa0nkiKiMf3FBPFmM8DCP5TK3S5HRymOvAmXGgeGDtSAxC0EnYsnFGXT8k3wwZFSG1hlBen9zGQ
YzuASx3RHFlGo4mid4VYQXsa529/7PPw4BAPypdyIX1Qw6WtJG0WRWZv/3UZfu4D2L4yVDmBPJy0
ByKtPJWLyAb83vPbcY4Oua+IOVPVPkk3ebbqo/N6Q68ulMD3sEZIzsIp2dC4BhVRNHxU4WseuTy7
TQfIRMkB9ycGuIjMCGjgYrg+p3PY3oDUTkS99G+pmPzE2TDQBjVMg2IqrKcMJL/zzTNzi8UxhYdj
xgUmY0elxL+XZXCQ36d+f531Ktp6Cmd4LREBUnwE1M7vXDuXmE/UyTKGnwrS/rDmhHBRFAO1g557
YEDTFNAtRvqXgRVPVfvWFYBOVtcuPY+jWQu6ItoJgZwl0yHLY88kOP5oD6sRIj6Np9MrP3anHHYr
olp5JEPPMWuNACtkZ9R4o9Ytet1yIS/GfHHM0TCw2Rraocwo2WlpW2urntd1SRrhc+R6hvhJK9c/
CtZDvpSwxoEr/PlMcsHusTwP7W6Q5tuZj/GJQyPM4hIJSLXrQsgK3jQ+BP4AehgB1cEvLbGtcz4B
0inYLGvvHKU8kwc+gaX2cg1vvdFjN4PmRHDJl8HLc+mOAuUH/gOaFMOUXsc3wJ/CFPce0Tn2xPfF
B91WFvCcXsyMfCLByEiF8dQpyVb3LZ5041f8DtZIwUMyAYKvzv/8aRLme0+/ZVCvf43v1O9ksSQd
F1xPiZ+S+oW+EEThOTch1GKg524G4CnlOOd6YSP/HjXuCTbg4CBKCDzSUwJVgN9yKvXHy5Igd8wP
r/zIdhm4T5mexc1yUgKIibtXsTJTgiWExnNx339n38ptCgyArXo5Z6spVDe8vDCD5HewvOuopxOW
Io5Ly3bt+A4nChL29EiqGerMb8YgLS68cX3qBGcB9xIswF6dMMJ2gucY0N/Jz+CSk2Hf5jRZTYk7
maTPvke8Mw3g2lsPzI7xfHYRVt2SPKI1Y+5kFdil4o0ThBAayo0ZO3vz+Q7GdNKxnQRBY0lE6NLt
yRkPeKtnKdjo++lL53XZYS47QEpi1wphbsGToZ8T43dRZEtlx76OqFIq6UGwZQvB+NRNxups7AzJ
U7vc58d3aoDjw5UXmhuRR0G6hRwRZgR0EqMo7zYF0PzsdxYDWw2n6HhVR4BX2xaEPrszgX50jr8V
oTFzdg9TLaew2CvZS0EQEMbwK1pVnThT6BZExA7Ec2EDCCEm9G3t5ZKf9zbt2kZ46vwAqV4r5iPs
R0INjAq/0bHIaqmdxBi+LW7MvynfuGb8pF3T+DmBJPAmZ87rp+fkJ8yJVN9RHrVdizcvaoo8FkGk
LUeVClVf+15qZ4Wob/MA/7VpKWDfho3ymnb/o3sFHaoO++Zfxnk6lDy4WU+DbXHs6yqd1BGL0crM
ZBhsth5izC0PT4OOHFLOOviA8UHeMD1/eUfjFo35HGJg2M0wXvAi2Y3aUzD9oSlsjWKDyZW8Mgh9
GgY+ikanwi+DGSNBp9VVW1m1SNNCk6kG6Eb8Gw+eYHwpIDzvekJ8ULDk9T1DHkZBX8as4wvPrNXl
rWnslLcd8jaFe+x2gx1tVi09pKRCQoGsO02DkLfm59S3TrSTyyUSb89o21RSgLYrVUFYmdr5zIC1
uzG2kQ+9mVsyod++X8moMXbp7H+jk79oGuneE52RPWYb6bRhnyHrFexO/YliTG7i7bz+lpuers9q
r84DzM+VobVNZ70i6nUydcCcTqJAzBJMBK6aC2L/Q2eASm8GGs0/iuELOtagzJlg7ENZgta30IAI
uYE8Q7XeHILMWmRpBT0vmvRFp5R7TMt06n160luJTtrYzePBNVI63QC+8StUJyUD9a8dgUJUUf5+
8XWfitmPrcG5eTKrm2o6e3mg8aKykNoSG1mEgPB759r/F6dUDSXy+wO0UW7I8pfYWtFN5a901OpW
1nQr3TQIJXhreVproSOORqzRa9L35pPCV3SLzazum1UX6vC0w/63AZhtV2GwpcELIJYKbbr8PekV
STiqtmq9wZ8LcGqcU9QaD3SiuHDjU4Wdp4RJLTgY+6u9ZbBi67gCLC81E8vjNqx5qv8v5pEDpQ4q
DNSJa/HC6RGfm7JzMMVWkyjg2chIBaZcLEM8F75MRXhspR/DcCpEfDh3RIS5Ntc21zfl5CBXg2sX
htsmg8Ne51Mkf222yHvZvj5Y2qpT60rOp9xAtxrLn9YxbBK4qNPagqYqosNSAwI3uCn6T9102Lll
aXoktiLMEipEXJaztTPq0NQUcyNc9GtoKyVS6QonoWgHpXDeC15zRImOJXmxg5vNahZjs1Rnf+QS
GjO0bZbXDsyptQyOuPlkjdXD2Oaf31flavHQFqMzUw/QlehlNbjaHE4sq4AwQHrYVIfyFcwYI41v
xVdo2GNbJGUic15AxGKD4fX+gePAXE21FB/qL3z8uNh1/TbSfMJX4TbGHAWzIPMBTGgFnvQYz8VN
kAEzzAwOm39jlYXsXBW6Asv62LyB7ZQI4e5Rs9be8DHIVyGiNdNMYGonhgN80zcW5/G9uxgVtq2a
2YZMtlYdt1i3DJU156jtwp68jDJN2Lt59ghRQXpsq1623NYITrBxvDLLI/+beFRO/ugdUnWEnJ5f
z5BEeRwUTtiFajQzjRLjzhkYoNFqJIzNOy3ZN1+nKTStAOhye/0xUw7JKA0uijIP9K4k62UCylRB
uG0AU7CS6uTKZ+GuufOzKEZJZURmiou68HGi7DCdeNxfvGxPSQhDxODc6NlF4Wy0/bldLSiJMAc7
OUQhJwKbdD1HahlYSwR7T43RdLKi0RJcOpQKXsGPvby0HLMzxa3FrD0IG+ECLFLH32GkKFcAGJxI
wTmhlib4Rz3UNq+PQOk79be8Dp1mNu2LTydW0cJTgOpB2+u2oAfofMG3IyOv4nqPy6bMPEuB+tat
8uglSRM4cZC63XCK3Mufb1dpqVqMgkwjcnHis+OULRG6wS9CiLK6jNNy3iUsZsUL6pUCiMyaLJ5H
/xhU70owVJofGN2wwUUNx+2xsOA8GmqGwIcDXDttrR/PT8cegI4i8xMINNPg4+rpgheIvaN4CJXV
iRW0o48kPG4yk/hgsHtvnnWvrllZIY6a0UMHdZQFRMEmuj6Q8fRIMTrMQuBQcLK0ekrNRLPLkcra
zAljFHvl718oNDLMCv8FBA/RFguMiLmuRwTYusMwCJgqUYG9hdcSf7o/JHfwkFUWQYq0riNC9yqh
tzJXTx14P6uBFMF3U8Roxr6b7mPdwJdkW1KRW2ryzXSM4kure+U3yOJmaiuZG69HIUOcytsaGWkp
k1w/HnthJTykZcZFmSrMx3Khy74VQpvZND7rVLrVIszm5RXB+MDf00BtMBLFC3UXB5VWgxFIM1d/
0dzKnDEgTuSxGgl6PGo1pVAtpzdTPkN/cwJCwYUV1B1/aSVa7IXXAIfpbGntJWih6Pgibv9ow7i2
4JE/39jXkw3dHc9hlD+V1ePQafz9Wrm8q695PsdBpmtufQa4xKqvOKn5d1E3dQ9FzxCXf1Us6rrb
yM3W/0bWhgoUX5jao6cdycsrS4qKQTpMAuNN5teqTbTKdMOBCyZJsjR66XvVnspqIdNyKTR03baJ
YOzLtHq80ka73PI72t0MTTFQFwSqBmS/LjOtPp550eo8YahUcyXcH++9RV5lWsWYnVYDSWApJBo2
x2daTbCmHLuoQArOwrQ7XOiubbwhFxibr6MIJs3EWdHPVx4tC521rnHe+jVpzPgeMgzV6wiMwGox
6EYwU+TXfxR7OcsZDyW0h3XyTdaWIyxbvtty+tWDWiM1ocZ7F9gQTQevoFO8QsIdiOOudpLqb0wN
KZvXxrgXzYE/06LXDEKz6m+5qPr+hdynbKlIaCcelIsVOlIe1tC2VL+ussGqHBjRAhGZN5w/MUX1
exbsRjrnaEOf8FPs7PwomzD93Tq7Rea9eayl+vulcVxbEWddnaHxq1LoA3kjL5G/ykVch1D6kM22
DdeLxsQpq9UbgEYmfNX3ylmKyK6klMxOBzgzLELLrXYOhBMyqr/NKY5dVr1iJi2ZsyI21URNe36v
P7jE8f7mhjx9pvUOQyi3tCU2Eng+7jRXeCZxoCUM4htwy+oZbygDx6DicvXAV6KmsfldVo78NkmG
ZrloNrezsDGtIHsjEtkS/ztdaX+aARQTBsQFxriB4C6E5z6A9Bb6uCG7epAAb03AWKT0vIIsVNmt
uJ37DZ2Z47s9W2/j+Zvx2zmalHVfO5AqqpEYuWFkr2yNdLE+9Io9M/ivlfCm+zXbnzmL8OKXwAYr
GTJCCUzqGoRsJiaWQ5Kxr9vG9zXsQ3+gm0EC5a0+DhuOUTXrtAv2EYPDrcZJ0b44XwBDORtNIiHz
hHFvfgAqlxgW6J5qYH1x5dVQJjTNnaHWDiyl6KFLiJAb/UeFWZYh6R1uOFq9+z/935f24T6+Pd5l
PjWbMeKwniXuto8hI5GWYAbI4uYEDY5bBtKFZD6ZLv3eZeqrr11Y4t9DWFm6wfUQEz9Cck8SHSoN
vFLu/6x1jufTRJP9seOkGtQRzl+D2hVO9iJjhYHHP2OxJi2bsBPdpeHrNjB5PYe8nq3HuhLWOM8K
1FW7DgdwWQfeOmcKjdcxglWcJC3JLCmfsb9TUqoCvjhmjGXN6W/1GkqGjiv5LH81xnG6voQqSEBa
FwspyMYBN0cZr5b8gMYssORD9GB8OPeEiIEaPep2SnssZGKlQauJc5Sza9c4UgZtn6hG9CEIgB1a
6zpUt3WFt3jgY8G5KR23n7VqJ9plKDOyzjGKs4hIDBJiaTyFi5l6e6TN8jfOi8Kf1StFuWkxQP8k
UJjUCjB0EQhCiawFDUatMpA1dhR0tGb7IOJtJRktKjYyIOP5C+VHQRyog5ZTS3YP+jEljMnZWdYx
s9BdjMt32thg3junOC6CjB+/alWWo2JJlcTjwrZT/M3e/NTNsxqc1ukypi96eP10SKgZaFsnNfnl
/qXsFWIWrPfbu2eLzwYxjPyMZg2mUVDuLbF1SJ/fGHmfOtAFad8U3UC82MM6Zbvou+GF71Xj2CCp
w0yOeMJpxC23NjnBojsv8iNluyZ71UKedpwKcO9La73Nu9YHYtJiSN7/yamvs/5tsL8WATtwFyJf
Xst8jnWK464syB1LUjZCmaZajldoYTXs6SXN54ZGfzDMJacN9vorruSKE09XsJu/vTerKMkyp0xX
jz1cDswOHSVw2P8zF6/Evjc0iA3h9HYYtF9/zn3VhDkbaX+AxaZ5M/HTTpBSRrwq6e2drDoiY9TL
XUuxVEEX7ZETvOoMZWhIVeVmhCfBPEGZckifRUCpJeT6xk/ahxiOLR7mVnYdq4/ORHCzsNLoff0Z
hFeyBwDH4eIp6UpY0viKaUwZoUgl/EbEGNzzqgeYmeiIsbmnpSUaCDfXY2D+92GfUL+1J9Bw4SE7
1uEmDM3ctCFw9BOtoZuKd6qd6VA4HtMsueGwpXTq/eND+6fD2r7UE50QXVbjnjjEcqOHu8mt75nP
LFRJfm5xUexhZF+NdNIGedTukQslVjwrhMnnNCYyjUePM/4yqn/QX5FLV8D/qlPkSyw4P4F3ncWl
4cPcb505dL+Rs+anL/TmX2t4lm/molNysFTEDLZc2G1JH5NFFuvyEtfDUhN7Tq5HHqShPZZ9y0OH
MEbAwWmyyutUPLewdcc+4FuA1zqfmznq1Ufo4M88gtIEBIVCFtFMc7hS31laTmZFVA98W7qoZNVZ
LNBDzTJvV+z89qn7eRf3l26xfxFHHbG++EV4XW6ea+7ggZP/+u79tGXXw3svDeBoTTv+C8rzz/96
XoL66zF5X7kaNNzXcJX8YPj/LHYaqvHHfH/Voptnmp5w2DU7iSx8KvGwh0JeG34lDTuQIHf1Z8aj
PoJ45H06VnDbxUqxJoBbzUrzzyxkIUQQYrD1sWFiwU9vqDAonPgdT13rWHQjrXT5nnBJHZ5/vJGj
XTj+6SvOwGYYQSPj7xkuaRtU2aLkpoGdlEq6Oc3OTKsmD9iOQidHZdzf9WQwbPPLkuyb3kPm01TT
LWOwWuPss8qNFhfnYDzVdJxqYiPhfOPFvHOWpNwZV/L6CeXuLM0K99DfC115FuiL6vltU1Y+ceu2
0T6GqjHuH49s/RCD0VmWAJF/kVAN6/aGNnbi65TqBKyutqXXQOyrDBjaFRLjCfa2BaGIqEm8y7MP
Om4XytzfPb8CgaqCWwbVdTRaakKWl/tXNl+86zVPm3cOYXNceYH3fR+Ldxr0l1hibbRjwMb6kjlS
TGrrZB0W/O6L+3RYSVHP3PVhjd4931HiS4S6RRmjfch6nuD6OPi4yWT3ja4nn3IkEMzoZSBRKASD
i+xi/+K3Q6IpKxeZkQteemToQ/3iPs+nxGFyJBT+9atzIPxO+RD4Idb3OG2A42OCDDUY4TcunwgW
dP5R1ZiqrRCPM8JbxfHn8oLxkeFrmUNf3YrmMwLKutt9PrRwWWFwx+5hyouhlwUynmtfrair22nL
jE+HPciA9KiK3QSyZGkvmhvBLrb/CJsFAPjqjdMgLiAJw9iYK05K/G3LnUWcUIxkxTeWpxT8ToTj
tKber25rjwiRlKMrUH2T00Ezq5LJjHpIb23pgYnvr80l7PgZcy/8sdboMQAEgOX6HGG6MJoEAEcX
sHWp2Ixp/vPvesgHVsiZjEXMCvOxxecnMNUKP1mGWdo6W6r9Dz3I80wGfHTQuzIKDXPEEDOSB9wj
wcrUEI60dKeHtm++3Us3d13J663QxuHK7+mCttERjXSxpZbc6UTRpZ52ZN7MVs3YGFhjtfjW2re4
e3IZiui7CnhKO8RWOJkWvnT5rml8H2ABVCKBVlHCLLvuMdNgOg8xHow8/GX+3IICSxl0XnZmCJ4s
AZaAqnhKOuWGfKbjC/Rl/sznY+VHNEM5HYqfmfqokKe9Z+nkzc3/+AvaqiWr1IvkiWjcFjIB/loI
DkG5HmJ7+eBYrx8Gz1JILJ8SpK8D9Pf9+/P9ox40KsCJDiDEagZ0XHUhp5mpCYlr+vMdJnK6fLLG
7LmFDI+0Zp8okguOgy7ELW0uZ0tfrU38deburzdg0GrPmbT2rDVJs0UHITyrUdBnkDWY0c5G7hKC
ZVebjSNAiilThCEruJW3t/1qcesq9djAlcDZ/CEQxdW5Q0X8rcXkw5fMkU4aUsc9aZevudXtpMXy
17+CBwcI4N6hDh/U1TjtwfNT/hr66YTUPO6aRLpvY+JgItbvjfy8Rgmlod95o6fg61FIYIc2ndjo
hIw0mE1DHY+MIhf+cmBoDeFyq3kX366vU4P0tJW0ltAnCRct0sg0ZnoTJYB2fz4d7QmhWHKyBTYR
agY/aERTfvjEqeQpbAhIQiwuNjT8ccCGHH4NASxjvUhve0mvMgiM1U+CRTiqqf/T+fsrGD4Zs77O
NU1SZKe/id2bXqHz8JlNKMJvXETCMykzSx9OqOS/7AzzZkXE+rd/6uj19QZssVWTXAzTQHShJuL8
BCH4D3OH87eyssEvD7joof6W6kTzd1dIHeRTi1NXhLYhIWI6P6zAITB9Pf2440u0lkK5/yveF8V/
Sb10n93DDwJao6VQROm2HcZUWMXtcjJlAq5aDhIqDXb4jVkB/IoaUTvAQyke7CtceV7ik9mt74aY
BkftFqQBbaffVdRRXYGl9+ydt0+Hu9kobMS+P/+h2iJ6DtOtis7p+v0HD7WE+mTIfgQ97icKI2SD
Jc/XEiZJXodKUIVhndDWLZS12XWBY+kTZHDijndN/9IJ6rMLkManwPseHwBKguDW55s2cAW8OTP8
yMIcOGMK/DYlT/15DAHrgTwrVPr6ns7e1ZwbQLzqmPtGmDsYKMRbp5dnZ8DuStyPOrWOI2set0Lo
7n/JUPplBxNGSXYmZs/5y1H6j+C7OlfnFF28FWZVacp/Tnhz80lzC6+k3K5fBBm2/Djj76f6DCOr
oiit/DFjEQgTrfiWRKPhD0nWR8hzXcgLXkTrABBdjJ1c6+9WPRv8MPAYpGbfeeeZrJhIJpqHb1EM
ISTxSSDJsZRbUkGfN2CFiZzAOCId5slSlGu/32fmfU9bKQ1Dy8hKBKa6t1GxyWyR9EKRTq9qWCPp
FBz1Oqq+0jirtcUI1EOKkvgE/hqLQc5+aC0ZGkx5f3u6/YSpch3Y6aoTj6v7liwFgq1lCe8T7eGa
I/B7L4hWVjfKuWFlzALNORxkDbl/ZJCuAWJPgUlT5llakZDWw9zwt209BzjxMTuyjPOWjl6HKt5j
8W9vRFg9uEOGksQMUi8POei9syKECzO8IvTLltXB6f4nEMwU1OilgftJdD5lQl96/75//1dg91mf
kcaauM8Erl7hIKha3NwdzN5UudKYHrSQk+726uvq3jhNC94KM8SQjfbygs/2Exn4xP7CvB89kMWi
BBzJN5M0qmO/oKr8nGEdQlE33GDiYA/Ax9q0RYIkhrtp0yc3U7qG3j4EKKUsdeubZXlf60YHEi2L
R4kaNb7LXyASrYuwaexw5mlqn5B7irrMxHJVkAVNqP6kssI71NSQ0Ur5BzjpZyF40cQkqxuRf6Ts
PVkdwGSL0dmBZrMYgkYAkiOMOfjXM2LPycs2BeNkhYcrwIE8Qk9H/h0RRu+3QHOvuq23QUG6GWRg
1wW7UPZBBOURJS/akHp72VtQdORjFCxakXn9Wi90hckMWaj99uuGKMudJydkGHwHRGb/W6bWJACV
3bNQUn78qwGrLZsAd60byh8U/SUZ0AFQcsDLIHcdNUVGhHMvYQIoBRCgI1eEv1+F4igEREkTjDWJ
j08CL0OqggKjBzTO/SfHCIubZFZ/vjVHI+//3Hebkbim++YlqhYqZbiO9vZfWFrfyXUk3+2DaYqJ
IqwgWiF0Z5qX08g4fcb7xMQebcxl3OM946HLtpJquZvvdYoAxv1FK0N9gjSDFSQs5+21Pm1IWoP4
gr5zMpTw0+rp9i8jmhPTRXCYlBNSW10q0GhyxCCpgmsyQ75+C4BIU9HQkoa5VrQigD4yKQKuf2hU
QYmdIGciN+nxmhT5RJgX8oSLdTW6Gkkn40LBa4QdfM877TIENSDWt5qbRn6Q3H/5s8oXxuJJDHVj
8Or0C6f7Ls0diCn5bQBd7GtIL3WXPp/Z08yv43aN1nnLx4vbccoafgGM0gTUhHbDIzGoPOH3UweT
s6NuQ6mhjo6niTCujcNC/AeW/TEVCFfoPtVtiwmU+MXCznfneiirOQqnb/kNVpldg+iovLfCYYQ6
zYCjMI5rk17bVF5z8Ymo5b1c77X+5Q54p0haLoSPAMpcC8WwKQj8ND9VrVYW56vUJ8gr+lY45CUC
getrzvwGGPul0CQO9LNGVmZqp9JTPk9eaRwYQTrhoBYFCDBUKyA3UwZZKp/EeDPQRIocTiOoagdf
14v7UsKkRXfNV/hUh+1qNCMx485T9Cn1jx5UVXKdJ/Q/YkvqoQ8JLMaUvj9HGyG1MKGfoXAT+TKN
uC6llfh2mIFH2hs2Q6HuAGH6XTFa4npwVSiBhxksFEgfGLQtVgcTyewMeQrVlPoW7WwBbPLZgTpN
TH9ebAwtDMN/owNE8pVDUiUfvJyu5KlSQVeCY/WCYTCteg96ZDFfayeLERV378dnO6ayUCCluEX2
3tdM5HQgpfZRQS+6160y+msrZgr2yLsuuf9sE0sKRCB4ie7ecSNEfymYjldiLGEcDI4IiCJ9kCdW
Nk8SvvvGwZ7FZIEpRaRr4b4HocVY2w6LbUsFzOq9XZTVe8/7SElSsl6Y18TFO11n2KwYd70Tbc0Q
+yk6QLGrHBxcfPCmIVcDo2dtkqCPwJTCYVZ6m90tZlMVuDdM7LbWlM2/jiQ8Q8kKj9H0rNB5nHdn
K/QAt22rqImacjFdTqeYP1YD7Lp+aX7r0fhklX9Oo3NOJoS/7hYESpFt/cN24xEOJtfBAfgfXCkE
YkiDuvUgtrq6/vULqOcOKFBq7Xd6NN1yetEbqVVSKDYEOyGFb2CwaM7bxdl8jnNvT9V6OiyMnLaW
Ihm6IC1FO+A7dvFc9/pvqgbczOVs99ZZKGihlQOC+C5QB/RmGEATqQOs9uUHdYbk1WR8K4bUlvvU
Jt59iT+vfFWZJpnJREDxY6xz4Hs9M4CxUZjoRI6kFz91T9Guqa3SvC3hcr/YbUZLwWaojKO3+d+G
gqnXHkuTk/kx8Z1KAoVVjjWvT7jotrf76k1CA6AXFsLhlwOViiHCJuwkhwZamtlzPH5Xd8adZXgK
TEtznnD2rjoYh/7+GlVnbMopqgFOXxZwjF93teAyIr5XfwrpH1/vxbg2ILMhFcszZT287WyUy0k+
9h0QK61pOGG/sZmXXor5z50XDDp4DvBBCtk3xIm0k8KSJ9PpfPxC3dd8bWxgVbaXXHWV20qSeeNo
e+/YaXsrD5xgReUs849rq8JJuQKt79LVVF1RgOuoY8vRTm3xO7H06EtH3WcMNMeZJ9v4UGCP3Imd
LHQYk9dDj6wWABwNzcsRHRarJeyL8i16p7qyJzqxAQ4hQ+FVG6x/xrcDz6E0AvJalVzfQ+JCHCO9
4OSwe3sznUp5x4P/S/biYSlHddTxbkK/OCOrhYk981fkiYMpZPNRiRoIH5bfdJ3fi3TJAZ1IGHl4
Fq9H/DHnKKEfIHhvhDR9aWBjS+QCkx9U0mJEIo0UQVe9XmGIGlZDopbOqXRQSxvSKaCrYqTSTErk
jNez6ttcOlvKA7PUrCGPmEc+5XXLLFcHHnj2jG8nLj85644gBeJl7inGhH2RrgVytuSMdrYtiwXl
CdsL2pwfg92SVgmGEO64dQ9RGSBXxavSgA41QcUb/jDkC0S8efS2VziDVEtc+JSXpgxbHaqD9xfd
40v5X3URRMjPohi7hLk8GJQYFKdmiJbrQPy45wYpnV/AShJ5K2l0ghm9K03J07H8COA6KxxhFpT6
04Oe+KfZaKyZI07/oeB4QCcBHZwEDaEyXZ6SNIlgBCU/v1f1up7hDUBFNQsmh1bnFocVvQcWNWbC
9caUzYHBLt6eJxd1h3T/GCDBwIYgzt3EZ4oSJyp1ROs7L6rBNXNUo9IFa8PBn44HjpIYKCt67Uif
x9XEI7FIShY3UKEZWh7Knx9msF1S7nB282UxDsRsAKb8vUrszADqyyLblGZuJO2Y5DL8UdAmploc
OeBbTPMst5McpFFr0v9upUkmE6p3SSA9Mll71cntl9rTHx1KcZR20+QMcWZED1Xtjlr7OOvsXnuV
qR2K5aJ5WU+TqbajjIL5BHRsjNymBM1u82Oi6np+ryZ3XLLaWyzjKdbYNcx4UmOxEMIRMdGDfD48
D5XapRgQJLCO8jsf8BW1wACyn3ZJ8d+EcjaISDKUqQVSrSyPxDJ/wNElaIfgRmnyaKHg6ns1xrWK
mGAOwGTu6C0CPcso8ElAoMeM9NOgMR3ZGpjVmISmHTxAtsbsf07/KFwYIfufYIWXahxgz/6a52k+
n4dXlXsdwPMwyQycsIsTCYCHCm/rrZ7WYn1RqZb5MatEOQAlnDNcHERepvquTTF7sRnkQXXGtnS+
/XlC39ManPpfzcyquG5OGLyMmdYDB9+P00S+ugXntaUSTgxWQmAiH1n9QDWyda7ATizXOFj1N6WM
2TJHh0tgg1SeSt2y66jMnTakKZDFYOqH5XgEsn0JeGZhbiZCzdg4UVQHkLMN3nP3Ky6LHStTejDU
QJmX9giwVKy23gwo+TFoAXeGw5+B9flPBebOQCZCP0xyL72QyTVZuxBzDwScg45PtoiMNLWu5smP
qaZ2i3tPXdZynYG98ovCSYVeDMCTgbHdcxySvI/xv7RaX4X48BzMBJs0SsduTAtYqMKSCVcL7Wz1
Ej3woPPQugZcl+ySb/MMy7SF0KZz8DbdBdW5KVI1J5Y0Yrdv2bmlLF9uVCsjHoc9PdArZsSApzlN
YpuJl0zogJ6eUggGDLoAeJo/EDV3cH52KZrmZR43VY/LabF9m99KddbpZi9d9qQ5sSsY0WsEekxj
KF7Naqw0/MipifBbSQHS7C0rc1RciAm4SZudeehnA2gJQeFvDRpcpRgQ/hlCsIZRqR2doWVrK7Da
m7BkEWaSyqIuL+r6VlpJ8NEs2HdDtLw6fz3RuiRtJnMYw2DAppwJgq+McCNe2XNtK+FSQuncqro+
YfV6flfHED75cvoDBg0WKsoiVu0YSygVzuSlRFxmYH/cCbRl5tOTfF+YdHhPgkprFXuV9ryRCm35
0PFSHCCtUAwThymO6Fz9HRIFTwIjH9e+/6h+HbcY69b4aDAOlmA0NI3F/H2grB5QcZUuu2C5o7nh
1JmqebqOcI9SH6qC8D5DfN+YtVm+MoRjvZhvteFaVHqOyTOhHS4tKOATaXCInhfT20udfjftD7Ga
ostZfLbJLoujeHTjZKHo6VoR7UexExGR2iXBIOYrYfM8YhUiNppwCOD04YIPfmmB4/HRvFU65/oJ
UngygBcV6dQzpV/TFuOy4xC3vLJV/nnxtepTyfHS+ZaxqF0UzZPflOLXXttdFsAVUaC1pDUJMpGY
RZwsih05qVkHKWUJgKSLVvtU/yeHH+5vpB8hQ/AwymHRwxROvo7MHnBQ3cK9svQwRBOBG6SZMQyM
5eOS2n7nWPa0MWMOFAP9fO8LyRp0FK/c4+dAi+omK99ekzQmDnYaHAJmiwHxoDMVrRehmPutnR3W
15GdFliDT/5XWxVK7cCqqruBf6nlgKY8DpgZ9dfuVSipySIElqXEJgMVGFg3UwDCeW6HB2pKN72l
PsoP3lyrgJr/WS/H1MmdeHXXiiZBPHIdxjfNjfi8n+6MkbpJkoPJ/gTXL0hjScnhSz/wTtOCNY3A
KWFpQis1tHl3LjacTE/zpJS9WtsBsURi2ASzH7N9nJwHT9+tUyT5EL3go2W8xYePK9zrowBW08kj
AjhBzFYxMhsZitsNbh9Typnl9zqDeUJGeuip5HQsa0843JpcjD8BQco/1p0paGR4xSneY20W6ZV+
a7ePaCs85+j/EUiBKDtt+OG4SVzSsp8UA0/vnN0Z//8E9QFo/9mCrIVAVimzezsc7GlrI8Kxr7OH
YaZnAoY2VdxxSvxHH8dKmH8jKn1Qwvsbx1mtNLr7o3mKqRNkp2IucoIFnMDL0w0H9PIWl4jxaswy
jvL6CcAL3NaSdTarfDfjp5lMr4egBl31q7UAKXa2GVvFfBESbeBTNRCvkYf7o/cGNVvX+lheqn9c
NXAsD7fgEWgvT3VnJZ/TwByxIeo7vo03V6mKbJN4v0t4wANdWJPzbe2tl3zY+Nzdkii4YcIvhk+z
WqpFhZHX1Z5T3eLyGi1JHxH2GKJklEGDsBvx4mClRKjDoHiN69ITGSs6TZ1LCi5kuVm7LUl4Ct0Q
1bqP1uP0TTP6DICoecsQOkqs8TKN3lDBRrySqkSUfgRRGi7zBy8fXFrXY5GIWp3UlFHQP8vnX7R5
E+wz13IeQXnx5URlZ6iRY9sr+0DqCqMbGH2elrrXwVSfvargZcH2tiwdyMvA2jtQ6wkw/rDLQ5RA
f6pUY9hkPT7+iNzp92xQs5iIeVSBZ5X4aGFGQMLwIxECpcoZ4cGsQ0YFpMaLzo3z6deTvYtPL0/G
7ArV6n2wq8uT6P4w0hYPXSzCAQRTmanoSr4uBy5M3ra+qMrSeyrAv1EYOHKbg6tBtXyJJlKeB5/k
8dct8WTxhxhF5NaTIozkK8bJ1KLFqonbHTWyyHm3GIMW4MMzvohnJtaXUWG6tQtDRrB2e66YZhO4
206B3i/enO8lIqz4WAF171IQk5sz41Djt0jEVQj4LEoKMoeVI3ouKvJYAphcxRKQ7ZvRqlziZ0K+
Mny6ck7Itlycua6uTJ+SGPBb3V34JhETyLEhWkyh06+QVmwyPWAW0sPS+Nh73veU2UnVVgLN91gS
Y+7XVezADW1+CiBNHeyZWqbEBgeJk6vw3RqPyH9yqTscqn0vb2KHWGwYnzQHRZq3QyCRZGCG29YA
dgMYUedbDfYGnyLdkDftzbySWZYMZT5ClN/OzZ2nDZ/lSi01+rp8N70llmXqR9jYlKnXda7M9Lh0
yb8NdvRfZN8juGcCEH5zYQEhJT7UV/whvEcV7HUzkUBU6I77Fev4ASTZsef//VJDJV34O+IKAN8f
NUEPZooLVIWXB1evJU6tf8instPlRCQ44rJlpnULJ9EupAlM7zTdV8ckA4pZHI3GtxUBKkvpYmEI
V5ahxhGkc0uyIR9ca3Z8qsc1gSelyZRLvk9prbSJfDJLjJ6t8MgP2PW2RB/5XrTeJ08AglKfvCZ/
oqwv4xDMn4Wsxn0v0FZIltFENXevqE73+W0CBqdS3VUSTCahZvbTy9od1bRIwEGghDb9ZdufAJKD
RuuPQtJMvo2QfRLMfkT6og9YM9NKsHuJuuS+p1u8IFClhBX0GGpGnRaWjR8P6TLUw3q5gRSzaOzf
gAS55frrd/MwGJehC5pR++YFsolnuAS2azBmT3GFPyjYTWcqGsQ/AJJoimbyaHt+bpd7RprOimPN
duIhkg2UFBcu8fiT+i+GcFjg+8sO4uMCX+pMwkKIHYAc3UzwTXXdRUkfGaRb/XNijvgHP8Tm+RDj
9Ki++ryIQu0lBIdvtibdElzqx0XlYls5Pk8N4fD6eUgQp9YCP1f1cYUinA3NZaLoc+Cjtj0SdWRG
Vre8V45hal9+6my+Psvru8kuiCjOLE2fqKJ2BX/wBI4AQlZiTCYlaqIvJJxXyv9ASELtGgGXqOav
8XxToszhf/qGf8CFJBPhI+z4IIAhIuEtvjfuruSFz7Eq/E5wY06kTumCFCnxVotjlfaU4p9Aix04
uGIu4gVfQTCIB5juLruJPG4S4RNhUi64lzzilD0KqyUKo+w6yCGhShFVaVjGSpRWDTRVTgyp5BhI
DN4/R9AU26xM+RDfShK16hMRkkcNdIL5iGocTIV24xj7pZvw5yIqZ6Vz8qADrDLPMMC75gup7kXC
ZOJTBApdxV08MCy4RxBfuk8xWNnEM0YtImAl0Sbm4FR1vUOJxRC03nojTxdHECVXGSRbS6iCT2rV
0Urm9UfRTeyU4fQ3V6yJxZOkGM8Jen8vmQ3SrlbGgIIFm07CXrJruvoEXlaKDT+KDy247CasUTIf
4jlWe/ZWahf13nsUzKFXwx1mDTfhQBeEmPGX/d2P558TsRxH24ir/GI7kMcR5aRAKLWoyX/RIvTF
UxS1WkJGOkmjif/f99Fdw4S4MulUmuiWQIFBOROWbj1+Fy4io82VTOXy4uyxSV1jblnIWYFf2BQc
0keRDcQIsiQIT2BBOA7R4JAhmc1YSt3h/CcNcjlJ9WGgjK4B8SRY3q4xyTYBi4CGbDGEWUwOAtYU
puyDybrY+oBx+4HKde5ZNxT+iID5L05r2E4vF37/FXhC/yle1UelKIQqCjMHAbBwbcAd7RSpCOu5
AKMjm6fT709qn7ef8/61jqNUTkAVgShKu+wn8XxjdFsSCArXmuLmbszffckP306aa5OqnFX0n0e+
8JijoOgxj5qlWCBsvEl5ntAUgSCZPC8Jnlj/t07OvXx5MsSfPrYPghTtI3jw9mSGS9lC9DNNx0+X
GhssPi/P/yy0L7s1O5vAY4AcdAk2v1etk2IEyYgDn3IPrvU+h0dkh+owXEwCKMnZ71jshyA8oylf
C7IN1r6WAYnvX/dbw3eSU6HIxk36EwFiXDsPNAErVfsci/p6Om6F5zkTz/9BVqDUhc+9uX8ZV9pA
eWDVhEDGC39K4omYioAFh/PNGgVPlogMaMBAqxmVu5+QlEDJ+qIkVfa4GmvvvM0zf9OZdC68EzSe
G0itAbr3om0mjc+UtaGXtSC/yC31/uxdwExuDzs0Kwy99iHaJn6ECVYjZ4hcWpTk8/Qxo5qB3i3k
xOncv3IiHhTVqy5TxYnpUnhT1FlTXjXLV5YOATRwWihFtqxAC89KiRcqTU+MwOCXu7Z58D23ipVH
GopysVGKkVm0PfHwdlYs5LTJlqvyDxYyBYosOSdLrNg6CKR+6Zbhe8lSzp4ODfhvDdqT8rVF//uc
lbnUHRGCeKGot3B3CEpnl8hQBYuGOq5ouwB9UE0w591VaD5/9v74qEFAobRfJCAxpKIxIi0TXGJK
3de8mzvBfsUwOM7dU5/BHhklr+YFWxaosPXDyN3gtJ9sCVa1Wdf0+2ZWUjARffp0E4a6dFkzZR2r
w9VWAiHmtDTg3sIeQdqE3jSJ1jL7zN4YqueOWj/9yv3pCxB5fQawKDpP6uedF9hJyzD2RIAywoEr
iryjQYMfw3W8ZS3+5tAhE7k5kUQBXmQ7R/w5pFZaSUwv3S2tPJkk69LcxrrLg+Y6mopRVwK1AzN5
bvB8/dyU1zSt7pIOiGMjgDsHZiu62VtpSffgnbTeqtBG09x/ylQY4DzuQO4HxZsXuTRdsXKu+f9F
IozgM9+OGmATHKb/FfxUlIgM3CKZaLlORl642x0TVi8X/Y8p0vwfycCwNebY7XyHtBEWStM+ZgWq
gb3EYWbFaU7LaQ3KLifETh/v3oCY0JXQjwFx/FI0jqWOK7qCzWH8c+ahzk226i8NoeaarQu9uhMQ
6yvhK1OatOkIybGi/6Zd+80C0OBx06WLECq2cbV4telF73J8jb7s+SzAkuwIEM8ylRYNNmkZo1tc
r7Bfzt/amfH5FhVgj3UUV7cq14Ts/HhmlNvNlTWWzHb34qjKi7foJbAoAgHvAseiB1HI4l4rfk3q
MxaBI2PgMDhQGGZMoTtakXqqLx/dluGsUoU7VOwJ+JE0OFv/Axrn7wu5q2yThVIm6eSt6kGzLSQR
xlo2EOuHnU69sEWJoGY4sDi3HhpPI2XU63uNtrucL04o2ba/gKtJBspDRZ/qDacJRksCbWr7fq25
UoPYhsmwnuyXPCqHrIFzP52+0vNtxJcZ60T4zr696OTniJ2zozquxyP//U5l13ZaurO4NjFlTxYC
+56BUZThY/NWJaim73R8IfJqtI1gN5FvQWlsF+1xCb+wNAEU3+gYbTIjYsGqg+5i+fOipqcCDGmc
bKR5wAlnzbWBswd1iPHcmccTigyn/DbWuIjj4aUI3mDH94wXpdqEF48ZuGJigaM9f4AQdmzeJFcV
pfuMJXwMJEGNaw0bO6ccs4EzYCQPR/HGf0J1nTg5uCGHQheQ0BvYVBffbiGEnp0/P/a+kv7aFZoZ
nLAP42GRnqIeeqna89u+fpe1CccKWiQyuGK7MgKwU4sEGra0+D4wleR+D057ZQn8ntP9x0KXMefM
j/KodjFhBG2Xdg1/H/VINIGl3Kh+CDyHVPrZMn9OWBE9Yy/yHeVlLPoFMxrXCVK2kuAukbFD7ahL
MTRIGdeA/Jp+SjdDoAFFPe1oqBCh4LaURP+odIE749+jSLE2iAJAUiiQygnjX+b53mQxag25csjL
2accZzuqy7ZhRrLTO5PyA2/3RA8OycIFOiLW3RJ/dnsaFHHsvpk1HPuiWlzt5GrbbSxedMcI7KEl
6LkfUbpQ/hJRL7DAMDRDJI92E3bHPmBptZS6GRvVlSx6//5Eu67ipTn9+evAnClLI+uaZwDSdQMu
2sGvLkqRzcDgLpsid06YxOHQpPHoK1rfeXpGnMLrhVIC66e3tJiliv87WJoHigoiNU6A7mfP/lpY
jOn1coTTgHHKToChHMbV5QIFbcZRs6qsx7PWqxPzGhua4E0ihrdlXMtwpPoTu+AV1FvxopqycSkD
C341anq+FrR4T7l9kd1As8cc+4SUtjPHuS4VbyID7KnwO70lWRoISU1GF491gSiH15GK1bX4Iv/G
VRD5ky+HJSLQTiZa+IfDbuwZANbJBoI3lj+ZiRlllguelXp3hku+a42fd3s1JMeKbNL3kfrT4pd8
XqpvN0IDUqNCv6Yf+C32fcCEOalaTKbBYYd/7Vf5fCOehBiaLSyVoqDTgQfdWOKUeDr5Ailm6lrx
j73gdn9GT+7Oyo5E4c6XFRjnY4KUSn8+XDDDJxQ4dnAf/o1a07wSs7v/XR94eeU6eOg4QdTQ4y3p
2qbOKJ44Qkr6TzPkea/xINCSoq99+hShrAd7UiBOcWI4MZcqgcd0X1mnZcoIz8kyhN1SRFB3un+8
8UFfMrrcqr65QMWQlSgXtprYYporDRnH8DP3KlqUAQT2+9GATCl/clAeFFBm/MzOKa150oEeh6fT
Z2tln1USSIjyJDCwX07CKJZadsgsaqX3CXc7Xg0ET8QeLIlq4ZHEnuPgrmEVSgDVMaPBh00Vb01F
Rk1WXsUAygMwCo0F25lSIdp/JqZDxEpUFByqQR0uT6P5rDegAqCcV/BEelVqiak5ajY+hA4NqAZ1
ahwPjekSSiw2RuypiA+KUa4HYppuAOCH1GnRTVGdd2C3vsK+cWrtL4TGF6CJ9LG7SMxZv75v2mov
2ig0/WGjExQDC1yfO+jnYKe1dETe68TStNXE5qEW3fRltYCF62JFdoeJ9WzdQC8m6YG+WvgUh0E7
f+mIw6YP64++zgRB/+m3cqBzNyRGiK1kq/k7e5N8DvuQ6+Q2PbDbb9wKX8Ae4+IvHHvTmzrWxV3i
vAD1r6UgN1EG6Cq28rS5RtRLIu7t05WWKXQtCEkgEpoqXu3pbL/NeXqoR3Y4ArDQhiyLoGtvCAeI
FhwEfDJ1ZdkE96P2b5YXFAacqFIKG7tBmQpMQc1hALzV2Ld1OsXQKJdO+Rx4pRqPCmgyp2V6kfjr
u/lI+B6CB9fkwWOHbkeI+B6P9NGrCUT/68ThXRipU/TM/VyHuvA8dEPuCJBmdBZJdI9lO3oC0aSc
jNQYgToY+zKSl8D6UMjA0OTO11y6fDHzdhQrGEGk3C9AjkbPUJAwAS8To2I2v00wis94rgIBIAw6
bdLBfos+2lLPWCpJEBwVMu31UbkRtwVEKWWm2VFBQ61FMvuYGvct28xitdTrzBTI+LWipsdOJ36v
EK/dGotk1W5kLOi0TU2JvXQlvqeiWu7psbVEDXAA9QoFfNJQuC6Vre6FLyJ/BgDJxM8VMNID9BvP
B2LL9hvvZhWGFYljd6dqNguHYj6Qb47GTakXUVBNj82t05C/pLvuEwb6qDFdSL5RJTKHo+Wj4I7g
PC0Du60+ouoziAS+F/hbz4zSyJgl43JTQmEuUm1CDlHJfG6aPBgJyg9PjfXOjmoJZH8PCEDexhJA
QsYPY2QVG2VDbHLcf8XE/1mszboFb+xKYNCcmz/Gk5nsVboPDSCLZ4Fry1TDiKPPlu5krE7PwLn8
KuCe41qJDMU52CwNV+rJb1AyAHkBmis7DmsNnvdA15NLS6pPg/sZ0ZvQzfSGXV/rtvek0F+/Qs9Y
AnVeEYUdwJGkfO2KMWgfR4ryVY8C9hTRzeDFZi4Lvl4af4kx/A1ujW7zIc2bE38ug2TEYZawytsj
GuzaSlKhNO4/i3JWlSPb+TPPoUVKyOnlvN2MTM/E5NWTtHmLpQPVCRG1S4pLhxcdMO9PpGIozD4M
Yazw3rw0RGuXmz22tnKO+bf2XYAuu34+Gi07SR3sWJEURAKeM4QhKuGfuk9AGPUqMEIk7QQXDuHg
0cQjirEpkIDBYwZrFL83pcoUkF1S6a4BD73NpKYWU8Ja/Ug5KnaaWXoTrTXNH50Bvj1H/C9Lu+td
B7id3UqSrN7UnOU8vAqnkZHjL6bRb11MvS65N9S348VgApnOeJnhdAHGKaSWH8g2FKLEeMsDbVyN
LGQ2PeUlyDWZUAzkby+V96Rm5naTHimWcAGm1l+TTQNEX71norP6LrRJendob5t8sNcCM6zNrOAp
tbm26oQsc/aNJpeOV/H9WJR2E5OaSQOSW8wc8JVbdnue8iUa4szIomMlGEGh46pqV9xXHp4bPnKr
uFSxwAFj29jQBfbVAjgoM1u3Jtz8sBp7oB5xYsEXETNkhiH49YbhiEvp7s45SZ51U7z2nCU90PQK
WovVZY1mRAp+nY1Vb3kkPApSb4BsadOZxQrMhr6/jQBx/HLNnl5dzZy99MciT4+wodFI42Tvgt7E
uXLqGSB+mu2yBECiCqv4iT5MxSH4wuDbjgLRrKzlzn+RWIHbjwPzoTS0/ZiQC+J6Dv7YZ4T3x2r0
II+zEYViWsn3iyc6VXX1ZJCK34UamU+BSu3EPVNSxm3BQYbla+FagoFN8a8aHvACpwU/wUSfuN5K
ya/vDtCwzNDZIN8AsKFHkzJ76vOmKaF1hSDKoUi5MADgtQQZq/bJagNyVuG408iILvKKjJpF8yWi
F8RXPY+zRD6uXhsSylNibAS6IyXf+ad4Fjfqzj2JrgAng0zBCN5t3NNj4mX6C2gy6U25M16AELZh
wnaMQhOHSi60wHjTiIwhA0/eZ4FEgTMjtSXcJVpUXQgUBOVQzGOIjbSaaEuSgU8fb8SBS2Ozi3re
PmQbSchesleHy05eRf6pZMLimBV0fvwUQWOK7r3y0zlaJymrzhjKk9DlGXTClKzb8yetdqVJEqO2
cugDER7sCP69JN3+nPSMkF2r3vPJPisfWjT4ZWpxC/ovq8NgXgvtF4MJVuC8gSRGrbQLHbFUGtSe
41bbbGaygMg5FRU5l2BO62/nTRij2eMOYoeCTWe6VZ3SxRkeryXh5nZzCXs/glnIdQu1a3/sXKiL
6Bz2gkZlz1oBpKXj8ZknOvy9FBlbb4DvGjFN7FyipdcLEGJdFWEHZXBBfIxZOi3OZUuESSMkEeSN
PWGzqnlurXHSOs9pWdCJ5MhkaBg0p07cR1E6NZBNn9SeVMGn7GbHSgw/NgdRufZcziF1C+ECZ2rh
1+/DM4PDaFklAn7H7q1Ya8e2xtEzZ9rUcUefioz+DHDMf/o5LmojjCLLU01wEVHeJ1/ZcI61H8xA
Fquhc8vowGm1VUZfx324zi36wtptLv+Act9AQwwS/Q8/5V+GzAB+9ZW/s1hcmpUBfQPiKXrF6VNi
5S2znXNkUDbHWOzkl05W3u8YL61rK2TTRyhWp7YpcJUu6BDHBHP65OVSFzfQsab4wSGiYebxPI3G
pJNJzO7/8Xb5FblnJ8hJbSwLfaBs4Ns0sGoLZFHFYo4Yxin08d4rpHSSlMC7T3ahJ2RQOqy6QchI
DBH5u4MCDf0Ro0L/HdCZRxJx8YY5kM7PcWvHH1B0CSjJMa81+eRRBQ839UMNHCJ2CHT6QqW9XrIo
Y3/7yGGnnFIJdKLiXaiOPcS4/WTDrpjuwMUuXLe+DwlFBideGe3Bzc3THgdNvoKn2ute5AL1J33C
Uei41kgpoY7Uz+A/X7YIDUC4ufh3nmTYr/YEz9iuMWfvk5dQlz7aB3MtvjEi4g1Lq5y3FhPDuSdU
/p5jZ3Xwb/zJo4u3atd2ZXguad+pTwyR5Q9I+vOKMplGTcH1+/9peWoPW0VDCLilP++qFS/7EoW0
E/bPZnDKYTXR2/kQ2CtOEYHEdu/DTHOUwelGmMh5Db5axLfqn9OdW0Dhs2zMCOaHzdm+GHltiRD5
N0A27r+CkbrFtq1J9bMKBSVBpOX5r2UKEMHNFB7iIirbDkd/W0HoJh39OgyrWpvkCvKeT8qM7hkg
gKwXogqSRvBoexna2y5viCDVEZiFi2zTpJSNkdz5le6mc2a8fSaW1ypdJ8am2Gw7k9wAuGn9i0M9
+EjOGcH/TbEceNj3LWjR8NATFYH98aGNHo8RMCOoQbjBSOGZ7vAQnHmGAdKgtuHM3q2XgJu3V0ZX
/bIjiHUb/jbXdCAaqAQ6aKB+nbyCLcnkEMvDMG/+/SiV5HKzShDdys0d7j5wMXZc3TqvKqPah2WE
7OPfVDdHwhwz0EJrF8pfAR1Jxsl4voxvP/uacM0M0ny6y9UMqScTIB76dD50QtwX5dcRFYJlIMKc
n+H0fB8spdAXLBA2T9Yc/g/+nBlIh2vOAMxxcTQ0AnBooflSSH40GplCr7l1kRNGmYMBY4XonELQ
OCCGIvq40/ijKbnYrcIt1CR7ys5te4hUugKUWKVeGH1bTXCAWINsTbZlfpCn6eczFQyTECmE6FJJ
QTT+cdL0WNlXJQNP208FequUfjYTQ40i4x8n/dxHHp4FN1RiZ9KyF1SsBnfKNQAX2Ng/FrZ8pjZa
ygQJmN6k+ym3steAedkm//ooCSgiQ9hoLd1evA27opcz/AIkpRlrcof72V9zXI2udh6O3b4k5g4+
CI0GEUQ0ESLynefhv2XKx1EN6+3zvVwT+5OBUzJprhTGa6IDtLIDYQlp6uSYi8Wz4CkLzMfwmAdW
rqfxyVUcG2QJ4qz9MeL24yRE6urTzX5NcmbCZOwmlPbij0nQEcGcV/vMuiJULSGLoUfLMadWrdEC
Smd5RJnODayZ1C0wKDMgUgLjJTVtxW2yiegB+P2nYKYXUiZjxhAYx4j1c4ExogpnSnzhBxsQA0W7
8qz9VuA61fiLYvI6Jg7OQXbCEygH8bKMl6s77BxG4sDYtwKGyjeJkuwuPg29KFBuLlC+0XlNSaN8
wbhRoX+7bR4sVA6xPQG7AkOhHfYtkxPqbAC08TdHgBEEluKUxq+jhjrgI0Nvg+uRysEpJtf+DVT6
3HWxsg6+CqoOyJG07NpoSmZe3s1p4I3YvYXNr60YbMEOpVKxdR92AnKlVZEa0+sPAuL3VT1j2jMG
07qSMzmuwpJYOsgSNDeUDTzOt7AZE625S01RQ9Jz684lyKp/YetO5tqblSwdantfJvhATQdc//nf
sR74IXt7FkxM21kTKZi5Lc1psz4E9NegIUH3gcudjathR7MuWJ84tgpCx4H+3FKT6lWSWMZYmVkF
FQMx5UGxDBTna77RTasu+O8qHUFOZhKREl4tuXal1MjLFcODpnrvAtehtiT8vPxRF6fgIIoMnsR4
PY4Eo0FngXOeXB3bThNILB3LaJtdIhub+GZb3oVet8+4mdPB+++RTbjTlN4W3TX4MAFiI1uSmvdC
sJDoFPgbqPM9CHNGo1bFpfwPO0lxdrhPLeITY7osr0mfUXKiDkHFlvk/pueGQoPA6xFrFhL5rxEP
Son632i+B/OCTS4aX8y7IRKhXGWhF9gQlUPmzz42DvVhHkw+2CWWB6AiF6g/Ez92sVQOwgrHzeI5
rZA3rdk9Q+vHH+LlOCT3wijbKBKjMLFIdRTng3GazmItVxD1w8iovNqXWL05t34Cg2VC8WRHFW56
3j85FPd/Y7w2iD9zk2YvvzredYe9z4yPb7+wh2pNIG5FRFo4zlx2kKW870VnKXfY0HdrPzXzK7rb
HC2aoJvyCmrjx+TaNsQ0JBhxIz65HE1O2fWxn7E15Yra1sTgqPjD1X3A+OuB4h0BGkaFAaz1Rry5
Ltgyl7p5GLcXumflSBm6rHEBD2LUi75lDilykSvvqZV7RlQdtp76mJkEbN3iFn8bCBmnx8298t5n
SRvcW6JxUnHCUak6dP/R/JJMPOlOj1fxN3AEzdyl4ct0CniqxX8kMMRVlEBEPDMFHVtyt21cvBqF
7niMUflGj+FwUbyItBEL4iK7eVorns5tKOVJWjinfZpIg+aioV8RemkvVndYCCTaGXEhpZ3w2sBZ
28qetHRsB34woIkHhUxsSk9nMHTXHuE9TcL+SXWy31+s+IPz7eTwcfECoWbsOA0QheCS35mopt/p
Sb0TfE8AyT4qq5mkN5VVcZ1XxS/bnI37nAsP04fAv7MGj7JwaPFjRvCHXJa6irCGqoa3cNaXGftC
NPQQ98U9JCGb9eaAe0CJNOVobX0UaRORD/q59Gub7yVGv6nObgZxWIvZV/J3hLmIDWE9UZ6MgFkN
Zi51ItgTE4U0mnRCSSzyTrx4T6Kd8BbjJ17LeSXmgY39L+qgfLIC7fCJ4rxSr8c8P5urhx9bxPUw
+lamjMcOtYax743F6TvFfAcJ2frrwtlcOfxiFmMbRt+JPAmy3u8TIGan05tJWaAbPHed4GiAp+Ev
hMSDs/j5gUhtKtJnAK/k2JPEczLD+VHTfEJUF007LCplpoyA2O0pDCnYjs/lhkrReK+qn8oGjnGg
EyDXj3JKK7cynZ3OKBV3dE9qker8Nyk80z4kHHwTVuBogS3kdhV3SHQdv3RYYcP2G+tyZ6msjE3R
uhI6MVN5wthjVG60x6e7X6JE1c/QHuYD8GGm2T+7Y3pEkPbFXS3Z7vu87OI+RHvd2uOY8n03ULjP
xzm5KJyvoXCT0kaa+ORaMeCnj4CSPaaBxEZM06kXyjyMlQuPMyJ76yWTBf/g9qizUI0B9VdQcJvK
WogHFIaS8jfyw89FiziDQFVa9RL/rS6bECgfejKlYy2Lr5N8w/ARX/CAaOQVcHNLbO1XRocz++oF
Topvl8irHAfmKn4YM+43kz2OV7xqtsg0zsaTHI+VO6Q1h7dHucB7nz7JwgIHF93RMN1SZZYkqKIp
lLseeHYX7kO0i0yqydNs1QxI6RbbrFIJFCeJ5MnYmMkKUJe6Depgbq5JGB4NvMECcbhokm8E00Sk
EIFoSby82hdl/0816/raCZDRyNlIK6N2vLN4xAa4bKrTkS/nU5cMIp5UcqVVjJ3cAqsp7aqBta6o
fET/PT7lxyTIgaMQQWyCxJ/SzCcxJtzJQJncsH3IgoJa/c4MYUoJa/T7RNKtH/jAoalnfSZJ84EK
nS6FTqpZ9OZugKJ5SixhF+vXLSdXb3cdyxC12a7f87xtRlESyk4Kh90MWQH4Pd9SmsX97s2+Ah3v
I9EXyCb25Svi7qriDo+PpHJzdY49o4+LK3ADkq38tH55gCdBfzsnhZGU2BF4hltQ8uy3E/hwYDPJ
4mkdd42muq3iSXMXo7apHB1jt6RVdb3shY5yjoN3KbyUZ0t7jcQbCHVC8PXLeMJApy8h5feqtFvs
N/SjJYojOTkJ7mOXVzCW2bvAJozh8Jv6cNbV8tbIhO0tivuhsDt07L77L8fh9x16eCiHn9rBBxyp
J4MKnUSAonV3PoS0FTXicb28XQjlbdKaJyxRx+UQj9qUfNJMbgvZLJDuArsa33xfnvY7PLGZWidP
sBf1R2qVj5790Z73LsxvS46Hp+S6ebA67gyzIDfLhE/xyxq7RzbCATAmN2Oz3ZAOVIFSmgfnItgv
PgrVHLT5u64bDXBWGEetIP4mAYsKXc2unIE7z433rAk333IHIMhwEtaqzBH4SOeYWbTbFFnnj2sY
fgYur5DvdKQjP+Z9Xb+zQc5lkmdt8Jh3CPpXTvAc6BP+ktGCSE2qDaxVQeeGRY3F+W3L0I/lmeA0
otIYrMLN5jVMbcKJ0Bc/p3/69qOrLv4wuyCzZA33gDXpkXqbR+5o7RlNhrAnrs2JXRi8SJ+oSviu
YqOPgtqwam4T/rmak5L8O4ZZLUeSJPpPbuQnJUM0x1H6hWoZv/R6BIeJEr7JA+n3TDs9eSFwomBv
V4SphD5n/6uiJJUEyYfMVd9yzPa17CZS7B227a8tY0/uzEFGx1z22N6Dq291EGNEU7ZSYbtsLzQH
getDK2VvD0oa7ofM2FdVheJQnL1p4LWswMsFpoV1hSF4t53z239ohRw+S9HO5qiFCTViNeYR5Je9
UPVJjyQsgwpf2opSQhM/O4Xb3ILUJahpgcoqEg3Vf3eRIYIyI8+aWG1wIv1Go5m3xdl/H7Eeg3DW
9jnI8WgHKzOTFCfGkdWBOhqlnWGZTna6vS9dEVmXFPC3KXEJ6gXVsqRWVMkgqE5ZuiN15LZSpvm1
NBWevGDB72bOaJls8zLoMGmXw3JVSC4p6rSQX6fkEFygkrvaxJaEpMS/jW8zKw84SXMFS0zEAz8T
e2TDssT9V6KCr9P+jd+Oq7WkiZzZyHT+D8qy1/6kAgG2JJyXLwz+JvinSKUp44JkHliMj7tdr9I8
VvYoVaa1xsxTVByCPbP0Avfoka64wqpm7nMYtoZvmLv3oTz+iU8OARf0WMs04RrM3r9bH7TmpBNx
zp0ZUA7TE5l6bMhC0ULCYIUlkjS5jg7jEBHStzE7g6EjO2OUbZdLohlGY0GAZeaNsKAbRSYGqBiR
ijt1wQSn/5XxXYkazIJ/IH8WFzzeAGxg5tEXX0viQXQmmz4W3lAEDmxbREJcAISlDU+jNRZbDMA/
BWcwqpi6jwX4OK2L99SqJa2uOIn/wYRajJYctkTaXhZHriV/1bi6jv3PIDsQaRepHH1IOuj260R8
4iNkc3sUuHlnIqxmcDaCs/dBswBxi/2G9TzTyKXgLiE9r/YPRYtlE9y7ecx7MSm0h32F5iJMK2BJ
LkTAqpdHIloVcxqtDRjQ8sEJpLL1u5wlYX0kxpuTdyoh8jyDFLUHdtEH/1F0IWcw3CTH9t5BPsDT
Zaz5FhKSZE5qNm+R1LmqGCwJtIiseVi3i/pOz0GrubyoUe+V4yXmtqeruIcRjGpmlY+J6oXPTyEa
5P4NXWKWnQeqOUjXbb4KXwTM3tb0tTN+LSmj8YdXfDvwGRt+fzwqDcaWJGRsFWvNkHZgkppwiv4B
P20c3stDSJTXLtK/8LUv6zR+ZPvZkCuNj02l2id2BmuXF/+G/VCIavuXNczqd1aTk2mVRuofXcKk
D9LQBv//X4aAoRKubkIgZDp7+WRXSfoQq0SL4LWTimyWYaKE6Q9e0qVNAcEBLVuFAgQhhl8elerV
+3Tp3tzESso6b3gYk590qx3RnVg5qf+jx3gC3HTPJ5O8z9kFZdgnzQIC+Egp56MRsqdae42kSTiH
wCnMDhsJflEXc6KMzLGAoMvUUrvgCP8AXTpqn52ikwRbGtt8+9LJs4Vkru/yssXklXWgNNT+phyn
83fRNNHNXbfhGiF6G6XDE1L9eeCLm/cV/boYlMfLV77SZKYQ9c5fSB4X9SXCnFMwkLJHqA1EBC1C
B7zho4fIqsvOI839RZDchNxo27Wvgk9FTmTCJ4EihBDZ9mYDIvaKwadvvAH8BHR5B6244GsqzfIh
TdIMiHGjY8DBGbhzwEnF60oxccgSJL/MlMhq9FofOt22OErHtUi+8XD7grgdB+8BNvPOeRZc0rKd
JLkXDXbJGD2ZAk85ZWgzJmr7OhWhPjScqygmPW2l634jw197GYAC8iqDg0UvsfsTi3yqK82wpuqR
6v3Qx1PdpoiobAVsEuxzhEBwJ2DlI4UAZMgCJDhiusCEorUE9RN/QFcCW7ynz/ghCKJ8wGshHTHe
6z/cesYkjq/y2pDxDPBm79vO6RuG4YQv1kmTnGjZnEtNiL9aJ0y1hZrnokI7qLca4lAxmiQPUtnW
xpFrDLKvXALq9Ta6V36R3jmP1sMEjseycZAPA4Sqedfnr+OJP4x7Rrtrqvvb6vbVGNDLDNsupD3i
L+0etaj3MRHIRjWBhW8KX8DgqLhx9kzz6f6r61Nea3ZERucI+s97dG7TjQig+s5BeSo9j+GJsiwk
Y0dtXh4hJndK0xySrHnDXMcGo0ASiv8DNcoCgDGCVToPCdYiIg6FI6Syb8SeFmK9IBxfcTFBIuTU
3hE3lcJ2WW7WNFYvTUwyHRRE+Wr90KxFb8RDMxFakhGrRUPxiWHbsKbNfZ9t8jRiZnv4jqL14VTh
y7vfYqEqstu2oE6l4WfMJrbxeHYCp/R7kp7BGvc6IDPxZN6tjeiROa9CbfJj+c0Ndp/T5HGSsERq
Z1O7RmwAmE7+WHks30dWr9crtena3iip8aG+apVzvY9gENT2Ng+hL+PKV5LT8B0rsk3UM3xfFX7i
mw1cCojtVawKECYuj0agT7v9005l2SE1QfCWWEkU47vpbeRtT50D2HqvmTzLTw/v4dih/dUDEsqL
36bhwcQZx1lezhP8w8KD2j200Ck19NkIZn0Dgcbd/bGCmcWD2sYPFb2+XJoPRxGZHCo9Lfk9H0ed
dKWWR36rW4DET1uZNGx4Ue3SCZRE/Y4IxQLU29EoW+FdsnV9NOqaPBcpc99l+Ltd0bYc9C3DMISt
pO9hI4tnEvKC6KwIgewv5dTJIay1GuTDdY75nhDY9ACT5Xl0ORKIopzHl58qQw3noxWKJ0T+BnQO
Is6hNAhs8oZRS1AWyeVZfDrfTW9MMx9qWFRukZrIuAxGdILq1yMaZy3D/qYS/gIiQtUQxjUqZDcz
/rw+esJj6ieyxaGfrPmwb57NQICOEMgDMYGq98yABl6HyKnia/fB6ixPmZrB3bBg79+ZwBQq8ZYD
/LiGBGVbynwSYwfx5zoy3K2xXDPzedbjNaWMKRHh+O443puMomNCBTE1QEy/I0P39gfKaoRSR4oa
LXOgyBQIX+G0BoDX571daMkc1QWGCVJgufxuElnljNQP7zUAbvinGF8UgR6/iFBoVaKTwven/KRf
ZCtFtNSh6zKm81yw+AVZ/nourpw896Jlf+O2xO+HF3FduVwYyKs7ifi5wo6l2aZi5npTMxbOpCnz
opOoUn+tJJod3a72eR08kWDr6rRIHC5fSeFCHzxsxq2Nflg59V1jASX/awBWV+xUKxlgU/aYIAat
ZGJqD030XWMQfdtwvUHTii6nCJQha/R6KN0pQ241spzkzh//8sUD0TCucMCPBC/64PncCQk8Fp+c
0bJectD1Kno8FN3DTF2K/iQGET3x+9mJPGYngnK6ZsrRsA1sPGEfkfNGD64XbO2DHRxWOmHI4vnf
hmMcFlyf+GyiYtlf4Z4U3cseHHIakbB0KCbg4vPKlR4NU8HxFyiP/KMfMAhEqk6oqnaZ9t06/mZn
CXviS320wzqiPfaCh4zvSmwa2/FTPC75Co65pinZNcY4FLc3ySUQw8RG2kWzhY2NAEcAXbrMHXLf
6+6NNxRvai/cbOydfqHrodRJJuP8LSETtQp82/q507s9pSINIG3zVHN1ciSeQyJplk4gKy5Kv9Ou
rPuVIW6f1LiLRNP6fGpVT18RWubZk/EXZQuAKTzWi9GqsuHMvj6sipUICWkrp0sFrtTNnUNs4Qwi
HwANeud3pJPnHo9vrG7UlD4FLsS6gKSAS18y8QXRbiI15KglBj1XiTLo1WAjPCtdmna06yvKth7L
6mk2YdxADb2ezMxobmGXWuWfPw+eG4tc16JWyKVaTLFAUroyyLiZKKMRold/K8OWsPVPx4sTTh5b
GADbdWPmMF+qe3gDHdIy+l85gucvIn/KmpMEf4uNiFd/PNFEi9xwbvG6TDiqLP7OdHqSfblw8cMn
zVSYsCAAQj+eqfp9Ehb5O6cxmnUuOWcVRy8suwZWryRAevau7Qg41cFBi/GM0kcHrSOVIUKUxIsN
hAY6ERbxnqArCAt/da0ur4UqQZSvNMA1qvZrsn3Fl6XfXsnu40AeKbp2l/VDJ4JK76MQJyVIbkQy
U1At+z3UqF/koN9owyJmpqa/XYTNIdxI5h8seXicEa6PWetZh/rQzWZ5dY+Z3YFMb5O18l5djiO4
RIpNSTwBUV1mzuoCUN/KWQQfFRQDnp06Vix1QAxaxsi0XLP7bGbxcx5A4Aw+7pubCRAp1rUR36mI
l4OulgLl15p9/Swe7S04cpye0g38H7Xs1PDkM1M/qro52u5YlquphQVDjAfSiHtlMfD0DHXCsk7S
UVIiH4rkX6kftlLF/O8EDgBLWuW9IleZe3kq62APpapWv5W1KCcC7rEG9UKKR1X5Jf/LQ6iz8lcz
ILyID+piAmTSU7Gy16hjpI+s5gqUywOmheY0X97jEQR+5FQiV3MgGSI02JtKLXFJn2PSfZVRnI42
/G6E9Eiz99uGq4nmYu4SqSP7MxJdDoaO75ofjMTHkiTZonISIeELHRgc2KXkTgaZzJuJnZcYHIPZ
DLH78DeEReIHZW4DNpaAyxVVFVUQjIb9SkAEl7p4GyUeRZiyMtDXFgqYWvtTCuJwTPXCH6PKeMrS
fbBxF4fo1sip4R/Q/PtDbJZ7r5tgow8DRXCMGKsVWHjFDUY2Wy+VG3M2Kt6q0SxxubwrlBkYmWHE
+y0U1MvtsKhAEcAYn24IQCct9U+2bQHjoO0wRVOM+gTYnqc4UFVfA3/viTKsPTB8yE5u+KAz6Hzb
eEwu3erqDElZNP6cboqc11RqlxXng19fRbUtfgoW5Fcjt66SnfXhcpA3M8nBCxtQ/FihmXu7Gucz
jm3zmV3Fy30wIYxQSmcpmXHaGUOkpAf9Fj15v48bidi9rQVtOheK2UWkEshTpC3cjuLICUGX5+Iw
DLKBiJHJaqOw31XTMgx/mmWW3sR+szqU/68TeFQPzDVP/oO3Yu0v+NCMspXI7Fj5xhmvI83F+EFC
opP/b/yFNW2lQ2GsghEjcFg3f+VPKgLIdRQW6GOEHAc77QuMF+fi5hdrd588/5XU/XBaHwxDQe3X
YaUhsvaondM5C812yMgrYCgAQTc3qzrZoS44zKmPfnJIQSxc5+SVOcSnZM7pcuMi4OzgHA/o2/8e
riBnbjQjT0YVByXbUmBm9oGvuYSOwOUOyLC8eIhLO+0O3dV5jISC5Dg6i2o6sxHGFZRnsxu5PHKG
0hqZLcXl7LcbDp4XVkentrVr5TCs3zFdVa/7kvsZjseAEfamEFkuyM5m+AWIVPGvFc3twOPnnqCb
FrO2uFn9b1JIPoZWyitQheJYbJFp15JeNq+tW3AJTW1v66V1qOtzWLYIWytuweFH3U7bND/NLPRG
6e8Lnk/yZsJNQr/QIA4cbvuCyR5KVJWGnhLzpbmSpfjyRDb8dpyZppIoUC7QsMrHLaZwFbmiFdL8
iwzH4kPCheSoEyPzaN7mcl6LvghicBS21UiyI97yuNtTpnIs8PH6JSEkHtf7ZwpFaxvDm42XCPml
AfTvGxZvWnRAVQ620ELg1uDUB4GSq/v7mrrVuXqT9wRUqZaq6qYmZkQWi6AiRgVrtXAx6Xmc6jez
JuzSrLs5zOtkjoGAcm/bq98BFilNgLOFGd2RQzZdDLLyLwetIINWmH5ju9u+8JrzBdyuBHhEvGpC
2/sQUYn4XjxNnAl+84lmTNSzdmFMvyIuNbuHW847FUuQafjUqUS/RgvEwDegoia8jH7Xr+sVGMqr
dUnqhuyV2Fj53K2Xx5Rb6upuUdHwzoSS1aW9M0N373nZX0b4mU4HqZLvGddxBwW8VwFQGZdD04lH
sL5ABN3orP1lbmHSpdoFR8nx12FZTALeTehG37M2o/jKicxqWk0E14aEs1qsknX+gfthA6tmxog5
ZlVUHVI//DwZXSeNWXQmxDowTekAJ8DzzhajjC51GwtYKhnZ+ilFfoChXX6BjY5SHE/Bb8tPlyhQ
g9WkVQSZAtywLSKIHwvd4pFyh2iKzHxkH9mi5xS0WCN6frAm00fwU4ULlPqWpw7OHtiPIks/owVH
0xGKPg/b8EAM1qgPBdpLq/OcZ8ZfIpivp1BV+pMg9UOYdOSxIMMMvRHCc6FA9zXQNtKbeuY+1AvT
1yY2BqlKO9A47a4Boh3jAqlPPjCab2ztgAQ1t9dwskrRIYHIxaJHtWYbpqfrPFmjV2g1tkqZUyow
USlCjFJBrlaArLyvdEtEY5ml4M5SEMOt6uYj4gZg4FGKmXENqclxD15RDiL7SayX/4actpu/zIeI
ImFPWO2mIs6z5UI2xooPdnDWqKpcKUSpysCm5/io1G+i1uB/Jz8SpWetSNXdoomiSZSQdRUb3m/h
taBjZFH1r3m4h/Jjg7WfS76Qs+CmR1HoDTagM9vFWKIZE3jifaCMWUzMCu1zziV4+30Emd4H1kPV
bSn2x6NPeRd5sIX7Lh2pKk/LYDOMF7JVN5xDgPnjfdJ1ZiXxy584knRKY7z8Ilj13W3Piol+oOAW
CxRQDu7nfohsadH7RaKgrIE38a4DaHhEY2Ethv4xfhHGdJOdISy+mC75gaodx9hfgP+XDeKYnYOZ
bU4aiklX21OGzLk4mrnWz0jot+z7YQ38hNHFOQUv6imJomqnUnijRSU6I7w0qZjVBlIlgeap3Hal
gtfNEbwP0c1wUuzboWd69ZfzLF15eX+j5mtDUk1I/wU2Y60RXgMINSXHe+5eL/us/GTltaforobT
G/Bxd4SCw+FcE7lOYLBD4uqOp41+ife54dp3/ksWz6w46TaGgcuJLAx2Jni1uaxGKxZha5kmInpQ
4U1A5dJQe6ZqHkTZm/OEoOW0nmr+UJr+PpspJcgmi/W31m8nKxSwZSC30grbU4hRR70ilzRfYSGJ
/G5iXU/GGqU0L8hxrQTEBf/+fRpyZS8wjQLNwi0m1uO1Hb9wQDdpAG+S7bAkH9S3ZHlhH32vLJWX
1no0pnW61uKnflcxs2ww1ACu0CHs/D1hyMyH9y+sfqzi1C//CjDuzaklH7LR9aZJ8E0I2hfQQ0pC
9UXWRLZ7CdZjbzqKFp+SgXNw12eaBtomAVeegwL/Wo08VkzhiVokae1Xhtxgq3DmPFcPvgzEJ4rI
cA6ncobGWewNZSd9Iz9ASndZr0yO7Lq+pkHzGfDhxaGaz9BkauGxaEqdn54PqlWCzJYmWDVa1WLa
q6RApSPHfOckr4o+0J7Dxxs4jw+struXZdWbk2LLwpcV17K9hT3aZdARDk0c80stGHg94ob+AtnQ
Xfy0xkT1SB5awGH7z2iHoebp3vjeItyHALRdj8fu3S6foKxClYlx6ZIRuaUjgic4ctTMFRY6hFyO
g74/cUmP9gyg4uy8XeJNTjLO/9TbGyW/AnTT42/tnEdG7hUHJT26nMyADWBsHQX8FY71yrsQIjJU
wgQIGCFzoJG7NXXafH7sfC6hqhPhCBE5+4ev1gDNHAkPNTE2rhwhnuRmixhZOdI5IPzY1o/amb0L
RanHObW8qjpiXphT51tYJ7tSFZk0cYL6jc7vwMNq/hwMDapQ2NoVpYAenCoe1HLWyeaBpWzD3+dY
ZzOO1QOzFq/nv+tzgq/ObenP9IOMG049i1f1lzy+JRM8Vc73RaJGXCuEr1w12zuUbafDlL/VMkd/
yyuZX4FdyV8Xbz/EFN5nKGIYkkPuBAFqM/xX8WyytEm3JidLNliRK/z7WKQUiYi5S17lRYH8uTPH
n7q0bgU96fmsVRIOOIVGrPBC8Zts/Ry6ItZlXMdRa0lmpX8ELR6DENbasfWwbK916g/B7U6w6IKb
p8x7AgW+CXQkxoYCebKM7DQNzEekWtWrDmDoMQTNK/ura2BxPIx8jEkt/JfmYM71dvgbifsncnUP
O3GfF8ZRsHQ8gjeHedESD5g8rr2lQX3T4JiDuHpuOB9oCOosdjVEbJT2g/zYIjT1oMo85saPXU0j
gk5+C3uT28e6S8NQqjpdkYOPd6D8qUa2ui4e2zelQrA83akv3EY7ll3AbzElQkzsWdCRoZG1nggm
BfrGxks1Slm0lRMAuZpej3a1Xr5t5Bxhf2FSPu2XH7ToMrl3BuvmX/Q0jr402ELyhRsr2IYzQXD7
tlqpoLLtR5/hoV5fPxQT3TU8XluL3TmxrKToKDkeaxhglrPmwwSydjpVQbF1PWfNpKLINiucsp+z
C3Qh+M+5+fPYtQ8UfgirQ6W35SoMTY21ivFPcP+b3/QYVhdEEQhR75P/DvNusQqvdyPKgP1mnhmF
QcwTLEoD6gWSnJ2BttVB6z8Db8Hdy1AUVuOVpt40B+j/7QP7fBmgl+IokyqS5wahUojwrBbb8gHW
Dm/ZJEWMBq4FkdWEacKAm/XGHgFChwu7GHs+zP2/kzS95J1XIbId2A0YMENr7lYhoIAjK+l+FFf3
dXSLCOwF5khIoqeaHBV62oFzpRQA97M33ngYqXLmR0HcE12/0KNySeC4+A027fC8ch1vr77pWtuJ
yciUEz89wuCkCrP3q0UC1mRaSI+TLeAja39LbANGtT+B+kcUocP1V6ygstw8HLjfmis8aqVEx1uD
TfKcsOZAOJ0BQKkBa68WujNLIb2FrzoBFgOEPsKDnarbWkt5cLJQgs5NfBJPh1/4152iFCtQSLB/
J460GoJoHvvZSPr+8hNbG1cj+Vx0qw+4ayX1HN8S7VbG51zB38AsgSyc/temR2Qdk7yBL0Q1HW1h
M5MozJKLKvahrGAMqJq4XCYxx5fGTMG/bBA/2vzDaKjI4RqF0bRt3a+prRohr9Rg/7SKsX8XyyqO
I1/jQYk/lVXYShrd/TcGjzkH1OUP/M6OirIDovsgIgu7jfFNxBQFQs9mSmuEIAex1acV+oo+8ZIe
KBdIZAI08IOpJ91vAKdBiLP7lih7+dikEJBT//JWCBUb/fGnfGQ0N+PZ22dnUfu4E5OT5JKVGaap
Ty0Zb+kRe4XIoAlGbD9i+dGbYKaIkA7NNmharzOUUlIgIVPZv1ZLr6W31988lCvmAn/YXaWN4t4I
kjpgL1c3d+dYGEu5ANfp9+6gPrDfmKvR83nkabhgC0kwB2XPZxiRH+3O7FQtcd8J46GTYr9u+zfL
TEo86VJyBxPPgxbCX7vvyWr7N2WOjB9ixQOTFMB8JV1/1ZWZ+T9hwSxPSYBOs34mXmmba7s40Ra+
RFnHqm94N7bVIUrXn9HbiO0LtPiYGJmzxQZkZOyybmFrRzdE5b94TK/Gz2XifJ8GFQIA+ILlHCaz
T6aLw8JxBVdkNHA2BlgJW1dqETeZ1QRNRXAirvsr8yKS6l8XsT4q892/f0AnGC3q6iBUyasYswuq
omOxTEjXvBcNq5hGitkKQxbazAFgLCW7EEHnqBSVb0XFybj9rdJoyZjpP2tYSmuM7wz3VYOibpKB
lLzG+2m5EIJPbwyN8bKwbm9x4xJYF8yRDUuqG5OOIKBVzLmIlS3oaVo9llgqA5XMNgdP6DM4/tix
lp9pi/Kz7be+tr7CDI2RJSRD5DNOaw+MBy2TlfnD07lc2fMjCjajtTMla78jb2sAoDZcNb/0oqZa
LzStqUV4sklGutLSBCiaD/3Ox0Uq25mEo/LHaiYIp7AAv8I5DAbn91nb8AYoTOPaM8mtGAt/Nhiu
ZC1Yw+WyXfAufY81erf156olVSkOaAGeZUtTCMK4dsQQPSb0LSaujbvZi7/y3rPVLjhAXiuosZQJ
wKWVS48M0VWp63UuqofCAPTE9zWfuhusr0oBVa+2qYriW5Kxv9WqUc1kfbyXykDk6hh0tHYi1wFt
GybD/R0ZRzCy8nrelRAYucq1+IeQLMavPhHvdZQLdZdf7Kd+s3VG6St4pRaqaNAI3zQFwK234GiO
kxLsasAuVA5qrQgDJhlu8JbQLIY0+n1ivl5cjU/qZZyzLJJZ3NI7zCgzJ8S9rOcm2oJI58EeMaZ7
dc3rUpwtgDosv0wXTlHx+9ugBT07NbcQa81CEP3N3ATVwoug+GDMY7ERi1PazPM7NFxmh/JCuNCr
5P5JCziGN1ijxnaGyrAIEguO3YdcgMlgM7gUDs5pHH3N27s6eyItZulIa9uJagiOSEkx0G4sUn+f
peLymqkXB6/6GahiVo8sSfDl2x1MV8kR+lWlijQUZ36KEaLO1S8Udkn9eWKOWZuMVvG4zNBwLhAM
XyG6iQG7y2kL5e29PtX03lR/Kp7pcv41dbGrERP9/ifneCfNiB19yi39txwuLrX7if2LPWlJboix
lqR+iH7rDELzV23gL3rx6BTcHx2suUU28dbMJSqBB57rL9Q5h0KjY00rVUBeHoZf5dQXCfsH+CKp
W7ObT1v8kWTT+cq5Uo3OZeoffOHNYKFpye5jN3n85NGCHfqS4CFLE2/T0+G3wmq9qF+vaobwPg7u
b2c8hltQIcppPE/ihjnRIbhi8dQ7aKYUpiBtt5ptIE8JgbtCARORdXSvnS+x5BlFLWbp6AAh3uPE
u5ts75wt3e5utm6fGoymEMbjUuVb5Z+GziwKBZUvmpCd7IaMJRH/E6LsfXcc+msaH+XEihXoL7Ks
ynBodEJDSv4eaR2/Fq69uKSKWXrkjmiJyWIVT8SjNh8L7zHPhDhSZ+CKZvBWS5/fzY80EVhjaI3x
PfwBEyxilIgchMClTqIZOwE0e+QVP8JxabLgZ8gtdXa1cY1AFu+cnxEy+RaOTZqQCLPWhopITpqw
NVpQQsQDVI+hFT55hUbRBO8IVj0BacwlKIq0SnvN4Fbx3Gp/dtJ1v+3NpEYpCO6D7lT/9XP0il0C
TVphHb5AMeZLI8J++xQkiCABG4hsl80JM9+/E92pXEvGLdjKmCBW1Bwl/GTJ8td9BE72LLdUssTw
SqYwfF2QzjVM0V4k9d2EyU+23yKDERp3vke2ALJh1WN6HeDy7LTgpuC8czKkXx/JviCJjSFxnrQH
hNi6FCiahn80WDqg0Jw1Jt+UZrDlxqQM1aMFVuNA23FZLmJ1U4S+HGIhxbZkspE8mrQkX2soNcP7
T/HpIZvYlV8Xekr7w0knezYH7q+XgUcBGuEWgzgo25NICcu8+A1/dQEdhiWXmdlHNz3KwVFS9oZq
RUZZbaIlAxKoSj6nwuLxYrx0VgJz8Lm/gLTna2fct92Q4gNb1ajNvl4QDuTgpLdL6a1XQEn2RlmP
NqSn2I6WUjcKmHVdXoaZfXhE1zh+lIgaBGW8IsQPevUjDkVrEqPGX2oSo1tCfYPqYtewUZ5yZwwJ
+Oe/sQNzq0F4gKw3q6u++bCixoCLnN2V6s1vN/kW4qVIHYuhiNsHq56Yn1ThdT7OZ2XfJfGXtyas
XOEcAiXTRTObFzaqwwFJXei9Pd/wCNA1Cdb5wkmGzuJE0/4CW45Yh75Y+bOfWxXLMoOsezJ/3nsQ
a5iHu2qnrVXkpw1aiEkZquY805zWlsi3mFC3t40PC7nLw4WDCcJFxxQQU4jhZ4UZ8Jy/jG8FQGNv
PCgJlEGVqbFFKJgM7/fA+eEotA9JKinEQWIFRIyrUolr0BQWfQ6JdG5VjTh5VvTcWeCpiDeRDWRG
V146SAJU/7m26xyF0zP62BaDcJMGZ5ngSMY7SOOh/pt3amG8cIX6WxfvsAgx93yMLZ+0FVKsZ5AZ
ysKS68/1VnGOw+LqOGPd4QzQdG4clO6h9e7WDQmadk8zldXd3YEPtCjPBllq2VSmp4iwVhj5bHJA
JwjIR510EEXxLHCwYx6OpD17VMNiTuKKctlcELSqHC1pDPGwzqMi+iRbOPOBOjZkxx83oR7jruEp
SC/Iiq8HIv+1oYOThsO3AeNeNCeGuDQX3007K0Gx7hqbjbX6oZQRwmUxHDsyFlijib/qsNQ13f/D
S91yuaXCTeiWCDXbvZWh+43PS52zZmy+2E143e5jezNNVp/uTDoWX1xI9udoHXC9f5ObEtYodnZF
xIAvPLDK47j6nX42BJEWILWbR9G8Q3JpBcxw+Se+VnLXEML3T1swur6sLi7bmJx/irohvoCfOkBw
ItNJUG1SLsIx1/HblbxBJ6Q9cG4siwhbsHj3atf/YkmBDcy8TbNXa0FK2TqqpSVpuU9c++5qJmG9
WiHycpTK/+c6Kymj4PCrkQmpmWUYtBBa/CFqwLtHYhJwTB1S3ljOJqXmXKFjTcasHd6cZZ7jN4RZ
scxIYt1H5O69RcZoRD0yReeyuVsS1lr3QUhrJ6Jnhea+qZh0DIa5Otki/F0AjNiJ4NCV33GLiMPc
gMHGGMjRAtHcUOjo4ORvgeIp6s1EzbWKJOvk7VhfAeUADaCzzdTYiwvL36NrNju5xvp4nA1HJRhH
6Q1uA0RU/saSQ1TJ9eAq41CxjEQYd8enmi0zZkA49BWfKQQUzmJKMSnbvwlba/+Z8HD4aTzcMkAt
zugkwXnPbkqMziQNpJWFHP/qGklAuwad0qhPf5J2xREHTB9EnlTzFVtv5QtNdsbBY+yiaEKBF2nk
glrV/EOnOidr/SrSXYtLAqOqHvOg7IGrkKbDFbV01gcT81dI32Xz/vZ2Tw79xp+SBWnzRkraavrH
YMegGGI6mrKyJ0eWgQUhMhV2C9DrriecxQ5zpnzqqF1lv6iFp7sX0HEeTTcxm5MUggdqfmlYHIzl
FwSGrScSzDe2Wytm6wPlfTaRVQ8VZ9B1g+EMSsQ+SKtLBB79BzVI7/FghMFtBvbJoAXJ7SKZUtwG
kQCcD/wyMT/RVYZRilXwdbxZ0Ltiru7n5o8s3HRUgF/Bh4IbaM+jA5broscQECSbgpeKblrjTMOE
ARXfuk5P05LWxcsw8S3wcjrwYkpFsri1Ci1NP+AOpsqrbAmezLT8kcztWb12jjmWPIpY6MxhcP1Q
RtgAgQJyKJ7Sl+zjRc0r78OMoYhMhDtX88QePBsBE8hXEfTch2x3ZVLJ5O/iIb5zHfe9LJNdh9k7
4izCQXa7W0aD9BOsS6WPy2BnoeouOj4cwT2cUUsn3JLD/TfT1gxwO6qgNM5XgipWN7pz4jBnLTeb
RcOciP2cHNMy66Wky0zJS/HacITOsSkaBh1uEowOzvDhZbBrhcdVlf4XO28+xL0MAuuRMUmRYr+K
EoA1WmdW0wW5LrAts3YTAilyNv+rBW2EDEDRCLJNe7H7WvUmXipSJnIYt4BUU0W4HiGMrf1XorcY
J8y8qriwdeD2/xCPfxcJAq9aN852QMgZYpGouYOxdscnpgIeGy7+z/jScQvQHIT5VgTNV+EK3nId
PUU22uN2tNvjjzr5eWfyqO676zspYChHFo8E4uTW4SRNx9P4QoP88BO6iEKKSxxM2Yoix69Kj9Al
Mrq9e7otm7ulv2pmWe4xFfwgBA0hJx257TI/xN6My+0EVepz76dZ6Xky5sFTckqoLXutc5uK5A/v
sByBrtPAKNGP5awlZiWRFTrPlFTjzCVBdGtXWK/LR+WfZSK+Z7Val1EgrlaUoBhMMtDf9B+DynoC
JVGGyvxdi1OQAL1ck8D2j4BchOfiLF8YeKwSVDMTFmMSANdLWqc5T7zeebRYldPdnLEiyCDjJ09n
qmF+dT350W+dxVz3t6mPBWy39VAtb9FLY0JuQNUs/MSCSq7v3wNxpfK2PYmVDUz3VVKvbK6mFEAb
TqS2AyH6KHySZbRYwK0QeYJAcMEaSmrxHspLiLqLxy9EdnBTxQPs8rwFsuR57oVeI6uLDg30doID
eh5PICfPk4vV7Vk9eoyDR8pQowN/TySmver58cBOEvj1c5911VPG6/lbKb0ZXyMPIIWzjIL0Ln8r
tDJkgTLhhHyVuf3LnqL9lcBDTD8lFcU71X/eDAmGu14jOtuSZLhTmCsijuemmI7THZrxEtFUM3q8
Z20VFNtz2TqjkCG/RsXqGpCmENkiqYWvf890SBklxLAw2vNCE9a3SlsB7xro5c8Djji+CCrU2p1a
SCAelO+T48PQDjCZddLePkiYzyP90R70V74NZalmuMCwfFiOSUAKl7u/VZ0OJPnZU+QmVj0KZKpL
y6AGR9U0sgWOQ/M8BrzChh02pzBPhhJ9EVGH/aj1e2oUyQoVBV1rlH4Fb8qzqZaJedGMtPoOqdal
1QVtxih88go4aaqk4V913+o1CySPuLIs3l2/f096Cp5jXWjr3pLfS92sVUjpmPsJqY7cKmjg9n0O
OJ8qyfWOF6qsn/ldWMC0bZGcF+XKSNDPrMWkNpPG5Z9lkVbEa7H/xZJkRMne0IDPHY12zF0ACIJ4
BIFXHVhZpIRVbYE1R3SNT4FaPVL5SwREjgVNIhCXZaFS+OupgwPjOX+l4BiHIks1v3SC/UXJ0Aa/
vRa+3q3P3vNr+GzwsFKDufhpiB3f0ngq+gDQovhSqWpueWW5Tf5pGLmxRFgxoSpe3t2EcAiGL0I4
a7PZrsxYNYh6o6tPWapr/e/s9zq8W44U3VyY9CeKU+GM0yx4Xj05DJxH0HG0ll4/9cWqyUZw0lCk
Ye1kMsjjigt3oD5XYJaSWFrdbu7voM91LmKaYCgeDiCdlMouAbFQDyzOKZEZ0a+5JODAz+eb5SAz
F3hxJtP8YMC/oYVYq3w7N/x+hb9TScZjcc7HOd6sa2mTJRoBEZxUfeW0RoReG4paz20xdE1N/N6q
1pG49CLcWzdR9ujpKY7hi89OkSG3EgjsG6ukIS0E2CbTEaMRYfQzypxlNUI7U6EXpbmEz0CJSXAH
WnfPm1CG5MUE3Aqo1FsB6iE+Y5oBRhpO4fSDxdxH4LKtSI7TzuiqGG1k2Ugbf6h/P9XHqsHq3A3a
m/sNKWCrcD4TRKwvDIWZfg5bDhwV9dQZvhzI2aR2K6HBAT+xEzpoiNiu9UTbYs/EWqd4e48QH7q9
9pGBanAG8fpvl1AFt1uvZ7c6neAaCzZJqsjBh1y22lPis7WHjyszv7sR/U9m9BBMRnOGRNKHttmL
Nylt/8otT4UCqunSL+PsGcDtmQEYE0MOOxh2vMGZRJntQePyIc/uDbwZfN7Y3dmghu/xY6362OQf
Bs2pHXoOjVh6nyPhOkbfR2nEq9BRWH0KfUfuue6PpEc6ZKmu0N88WZQUSw04htTX8Bs6v54/LAU0
f9hEJSjvniAJm9l6LjqIQTG2FXb3kubuPGlI1b5iaQF+AojRhD+2mqy0hv7sV5MyeseloB4hW6ml
3gm2ZWZ9JugBivJhpl7KQxMIxaRBBJf9UR6KrZen5qljz9d6Y4fHYCEDH/N9+cp8wB/ug0Nxw60D
ZWfocIsLll2kyAbx/q6qaeNON3ds/uHcARamk6FoLNf9I/H+A14lTmd3BqHWqHrDsvuegcrDjins
mEjkQPecfaobFRFGoYAB24vvyHAiEdWozTVH3OqSRmRAjvOJMd1HsVjl6xVvnd5N/NQIg6zARnaR
ecBbuNKfUvwCrwjVt5BMoEpFDKzglYPqrgGjvnjKnOiHnoiv+cr/SXVAukRf+A6ZEhZCCGJJo0aE
X+iEcF71lWS77f/V9cukTgRlKAXPiB7YZrhSgzFhMiEpUiPwPHo4t4g69gPFr35qQPXndI20oe6t
LHF+lB/OMsmXsu+W+JcZ8msZPwCffPT8W0zTNwjvvWgYC0tz5y15OQ6JL/QsDsygTeQ67+XpdbOw
cxghX7YP1A+qGCM6V+81QULsXP6wd0koexTvEDLx4dqEVrhJd4jcL35pjj3it0Lj0ofgxxnRgiYu
pMLZ4WsbrpLXi/X3b6UOy/y3dax6r44r7L3jbbzfk/rRzgVVMzs5M46MFeutS0wd4SizPuVaZhmb
XEP5zrLD4j28YRqPN7gl5OolWmnwBEpi96JzBwhc9FmZIPo637oO/iOvftdOxqU3RHBCxNXNIlKQ
pd/L3Xw69oG8Lr5B/8uauk3KvhITeO8tGPm67DDzSxyVsCwS9B1eGP+K05gzaT6tBy1a5UBbH3Kw
ooHlnGbbB+CdNZH52tVImaBGPblPo/N17KOuyGhN/dSUr5WTPYaPMbiNBlssYNVf8W9AmC9C7qjQ
s688uodk5qsU4xecX+aDqekEaPriU6ED6IhxIh9xP9YB+IwZB3zFaHtTNVTnhrhZ1dn4avwTHqC6
rbe6Uj8AeGgCZX0yEPu1bkQMBq3HIw0+g/6iE4FC2JPlLM1BbUWUwQWeCsAughqYWpbwAqYVS+p1
f4yRrgnXeuhAmhlLIsm7QXZYX0cZN+km/4h/CYfG8ujgX/ovKbWJlIh+8WjRA043mDDGqRHvnZJR
VPp49C5fPTnuOWtjSahb/JSb+ToMd7klNnWgM7mYuYrVj8Qeue/j0Hlg0ZCSJziznTxfkVvziXSn
yA0Fidc+x3fwrJ7cyB1xfLzPv7xGv0eqU6MzpoZygliECJlW/a3a8GZbaXXatLUhBMQ1/Yl//59n
9GZ1R9wR7IQBzcBvwJqJKfJ/S/0HLN1jzyToTzNXA6qCviU+mQdhZMSknD9r3XWaEPl7hhtXz5s1
KTZrBBuwjhss57+23DOp38DTplgEAARj8Xhn/KvOe5Pi40y3G3mcwMmGazIkxaK4/KNmaJHyzkqp
ZBJbmKOzPJRTFjgoUki3n15E8AcYVSK5rfndLYnhW/CBRIq18dq08P5NCWRzNDOBMThrwPIx9IT/
SBw1itAvZKekudd9alQw2QDb9jdylMAFA0NJdi8FN6MjiZmyH81Kj0/qhGuSKfdUCySDBcN5z89o
l46HcLKq17SCY6FvCXFJISowIEDIFovKeB98gaMHMlZlzQl0kVRKmx6Sk1jDilbxs/uEamWZiA6f
EwGkxZIxuBpKXGWHjnH9ijgib7Sa2NQ8WX+YvkDisfrXafkThu5vDIzIsuJG2waxNlxgYc1LhSl7
WNFigchB1l/GPtwnrc8+eH0mDHHyPaL50qf61aHb0v7a1LUn4PJyNMybrRJiRjZJYKTCjlDzzQo5
SULJtST5fqdv08KDwBOv3zoS8vpim4YOVHVKNWurUi6LbXBzGsGOktKFFG4D4wXNyCd0u7PZIWTv
Try2G4PpFlgTKh6o7KT/8RHs6YH0jw1C4VUF+BZNVikbCbmo20vApjt4SMzgd5/q9qtYUMz4dyeq
vI7kiilSgeY/BDEtnucbs5fd04EdRAbZtboX29QFX90n/d2hOouwo/XUHN9PvlnvURA60+33r58S
XIc4wskbXfFN/uAIl3ApOAwAggPp/mLmuhzr53xCq6u5cFfXOl4VD4WX9qpe2OEMEzaLuiQXNQNh
upBXap/cdIiKZS5gyP6Jdyy4c47Q352Octjkph8mydb9eRcvVrQfI3SDHDE8xIXXWxoz1Qo7WHL+
BGiN1PQqWJ9mKZJz0XCdOHU7uxtQPEKnmG6InZeNK8V2co8DHxZWzsfZV6gK+ZY1nfKMTg3gblcb
2X2x7eXu3zrk+ZFgrFhDIQy+l3ajjMgbCRsgMgbVjE94M9luLisX577bEwR8+OwggvoMkEp1PdTt
yTvVSTZsG0SPl8XgdO75gecmDbhRgvlV0ZddeM4T/hi6v/ytRTrBW5/DtDoHJGGH7zllmw2rpOWi
ovY6ZMQht7PdmZWGyDrYL8RWNch1Mh6TY6eJC36OdCTOmfErO3Y6UiskFBh6BZegZPAouAUa8n6p
B1t/BBffRpDdanAbB0PFXtgzBXSkh1pGJ1+F1/TYnOWq8zLuckAi0yOSXtVj+N/Ey2WC3YuB9t9u
7GoQA0ZQJ1LkJb/aB2WFHefDQd9DUhAxd6x1NoBPhDDVgdgEIJZ1nADeDywNsY8EF5Nk0woUYxat
gyHmgiGlIRzqeXsmSA+bq+UHrkLfC+evtXCSrgXg58B19HPf60YiuCJ1IL/BHcU5AQFAoW0PS1QT
JNmDJb8lKhj9hEqnX6zKpqMDq14fu0Yoqsz+NOgfnFoKePV7nqeCJHzXh+M9qoJJR4ykL8bGsA4X
Wx9zDaDWgraNrnKFXc3cikO/OxYjRpvb9/brSlQAra/+V34hJbDlv+4ZXObwoJ6uFhRWtOXKX7HH
diOoVTSpKWmOuyEipVgwF3HH7tbzxRcDacEqj+uhKNppHCx94zC94zStr6gsU1ZLkOQSnrEycGV4
9ZVsCrBBvSKFey8DPUWOkgt1l691dgnSe7PODtsvofMShnMMJKrGmEDSIKo6cG9UKwrzaQ+NYURM
qf8o+TIZ7GCE2knqTVoxA+o7394dD1oEja446WUpYw5RslCuqw9TX9FkJKdQA8t2X30CM5bGgujL
FsQM+as6WVASYvXDky6liSkDaaq77PtFzg8R2s2ii3FTFzeRpiH/jFgkYjbbYynYwBxwhhP8DRAR
EWUKd9MDS3KKIlLojf7ZL4eID7MtPmu0e7OQuGup2ywFxBtWZnRD5HfUr9zzGqUbTrXH6Sl1gDeS
aoVkCETeQfZJqVhVASJVpYnXvVElXCn8eg0qKkt/kVwHkEpwJjPhaP2OFZzCqJsCtxaUqFQoB6pt
yvQ3M43u5itcxn7GvKAD4LC9GLQam7l9ZzwcPUey68rGcLhqJSTIGmLg7hm+N+5YbtN5aMgeQqTT
dP/PSJlB1ILNHo2lJWVWBN3JHNpArXUvBGDP69PHDmzChnO4zvs7gB2wcTsaOW1qT8uvHDK8VqbJ
Xy6fPhgmbtHyDBefrvvQ6a/8M8T+PhCJXy6q44lPCndeoVCdlrCanMTuXLoWKsEB0NB1V1PMVLtx
xLK9B5rTb90QWsFPmDsYzkYX6zMn6DSMlsOhaiHjzAxPaLMp5i9yEVRvWWPALce6Ld9W8rvPN7kL
+BGg6CTCQ87ilxIL7p0ayyLuX1RtpYlVXG8hXLuGB+GuLJ7SDz/Aqff6cb8+dLyZE0jBpPrczLsP
rFJclkX15/O26hPbcLLUnRBn3Hxo2oPCIZ8O/HORxU/41OPfnUz7TDZ7Bq0cI5LLPsLwGgHoHtAA
B1ZCA3BMrf70R7IVEWlZWq//N3To7dWFP9BVM9j83lXvZuX4WAtk5nwwQtPtfaxKOsB3nU+2upzT
VnHt3NcpdGE6UlNTFFQKF2jJ3VQteBhwJVFrVkM4qiAxucogZRA8Jm2kiu92Z1VqBxz/CSMmh20+
V7PGBc3Vb+9IQbKi7TRwE7k8q5XFMMoPDF0po76ecrrQ+YNEKErP+stkGdFmPrqyGRqh24vwYjvE
Mx+awSjvlpKzaEm9S/vmtzlzwQZnG42agsIxCV11Nv/o4AdGb4DBVVtExmXSw2jL+ilkcV7SLHH0
e9vRsDHxeLKWW3lxYJSB/3V8yXOlayE/yfU8Cwh+KKJ3smtBcvM3gicIYJvI3jZqGryn3NHOqOF8
YYqsnVzwCldjyryOkAXJmv1MyAI0uo+VbqAcdxm1quUJSkXC6nk96ir2X+yoKxPXAVE5jwXheNP3
zeCApNwDx49b7pCtq8ipe8UAMHSxrHfEq8AGCuy6cqaJRs52tNZxk7S+NQeItzFG2olr3pz3nsUm
TvX/z/C9bzpYCPJCgxJWxuuzuqJcudLZyZp7KUzAA7b41p3y19YQkjLHD7hLO9SosIHWAMBy5blb
r4EtBJg0WQ223fZTbJEW3FT6dL1b2GZUorMpvP1jNYf4HTGknVgbWcYsVDl+hr47dvL//Pmr4T5s
mlY1/DBgnRipuc4Xnp7HRCRrSlEIrxnjF70nSnOeqIh1L9/dJBWRQrHdF4Jpj6GEg8bZTbAgM7xK
JMshgvzGDjvCHrINGT/CEDxwEMEfrXZifZg6gPcIUeo+7BT4lm0xEWHgj9IVUHUpnNItyy+YSCxS
kdgaqTs2DjovMwEWVtgSs2I8jx7UDv8xtMJQaJRFvQ9KI0PXcXxjvRuJfHwGvfgJh2RXJGVULRHt
JbMmYlurLr8ivM54VHP17eVlhPYiaYk9SuDYG36nM6Hpe7xAiNHuR2yABPjceBccl+BiaVe5dlxq
uBTHVZcHv4A66o+mxs/EmqwLye+CdzBPsUo/1jW+aMWFg6tMTq2OxCCMtdA7G0hSbHL7oX2lIrk2
cQB8Z0mj6mILEipZjuQ9AkbQ0+ROh4bj4md2Yon/a07XNhrjIDUJCKg+Cl6FoWm1i0wyrdprA/Bw
M6b19VRu61A4SZmR0IFqy04vg01ybzzlW0pTuTelzZoVHDirQCeMFNUXLgcUe0L64+A81/WOa1YI
vd5fJKkqP16PgTOMjtE/AIovP+zWa7o/YKPt+1ArSmYLMmjjlA6NVK51bDgkmq6onKGTB0nsDams
IFiM4ownoVWwazmQNJgiJ//1va80lAfRwrzf77DIO/0DptXVk8F26vNKnqRUJW1KpcsbmCW9kpAe
F7ACGrOBz1lf6DWleFUZwVyg8BZIVKNnvnX3Ba3CQVr0t+lZa5GTeAHrbQ1crLsCSr7fyj2wpyL3
92wqURVjDUAAYGZt91xC1ve3FBs7801DlWruxSOPlK4Aix+ExpQaJEDPChxQp74WCXut45bS+viU
uo4779zYv3TcBSjc9KIPKpWQ4DXjGRYpOf9uKppXeIttUBttSP1wJrKFF++Dy6NAVe3zm15ZJvfM
NDYCITC4b9Y3WsXTshKq8NVJNoapEDC2kofylKT6Ju4YXYBIxMt72xyXFrLFKss2Y0+5ly9bJ/3F
AZ5fo7K7TO8nRbtHhHVWl6VNpAv9lZ4JmKHrdj1FEuMsMvJc8Q4xTS9XxApdCYyX3fSbDk/FxbwB
3E9ZjG7JQzijyyxjsYHpdBqodEqj24wtixEoERyfIJhVmcwIdZkXSbYEx0Bu8kph++Ni8i8KMRth
oGBWbQOhwzkJGiy5JU4gwXA1aiOjqbEVYAcDFp55x+WfXZmzJqnXGZFVdpJNrb4Qc/Fkj3WwFOFF
u1lkWS94iWNmA1e+HP8T/BpjY59w8li5I/mpGCHuVY1gFAEf1wJx1H1/FI/IwOeNKuWe8v4Fsk+q
GBHQC65xAdUd/gJKD8gN97JBf6//20O4PD4f+/x4MkVln7gyUpdqO1Bffhsr6IpUYoosIxDBdr1x
v7OCXKg5zxOrF11vwl3oMfr9jBH4DuIp7WY6BYpCtNBV9uaGj2gvAgvFkSSsBexgXpNHHiFReinB
5gtbB/wLy6xGqXDRt+rexFt14zyBGpf1B1EM3raxK2MiwCmrVCPaCjJrSBUS+lasO1cEMxYYCA7A
lUXii4Yxc9tfAu6Qsqn/edUINtFXekcLzr9LPTMH5sSbG6hLUk6EtOUr6skOfvJ5oR0oPSjHUBDr
jnhpDr4se9/Y9wi4GoRrGazwPLF0ocnbnJEKFoKU7swnK4FbXyznZV0uIMOskgj+88ZFET+tVXk1
64tBXqcUl213yUMWlEWpYAUsJ/TRfWELxXP/qbGgvNHMWwOJrGtzGWHcCwLC5YEGVxlf/x8d+m0j
xOYW1Aw8XlTGt3HO+gYTbx0l1uVYFpO5BZvorR0eC7u2Ux89SwhUxbjR1/OLJ1YkFBmh+npV597+
xHPFlhj2YH/x7COVqbVM5ZAsJrzAO684VVhxwJ8BAbinQmzgHmfHlUVo2wUdS2HK99E+1Ze8FFR1
RkoE6/N4xuw42Iiu8iDzoshyHUfTr7dMWcCZNy/C9j8eMcEVUeLZEZbnfKxtyELRE4aqT9B4zi0e
03RFbBp9VyragAK9zTs/vVrZaPP/GBgYuVnVKAeKUgUrr5+Fs/wKRffHk0mdsWGrdT65aFwTjY57
m8gofZIBH/L5NSYcSjBOT7SjHN+R2mwkvx1C1wMJBcqlUH2mCYeMB/LBIFCmLjJHzEUd9onh4X+9
b8EnPcnOm27WTdwQSTb9gGUvsPZBbdIDbn3YCOZQvUhcOJ8O0s63ucBmzo9fNTCcfargp1HLKRwW
LdA54lAze7etW5X478Clk1QI7JXcZXLxP2Pa84uaJ8+81IXHzTb53sEKq8ZWw4eHnocSK0fyVbdJ
Z2Pb4E6X1RkmTU/yl0DHmwO/UT1vhT/RRdqX2U6wQjRUkI3LH5E4Pr6386+HzufsrGedF8zksmmY
RmJ3P5hR8c6AGtiQk4bO7SVdyMWNCMqBl7/Gv2peP63mo8iDaaiQ7ZnxzHeGHT6oM2BhzT+HPjeO
hi5Siftd9qQwrhulK6jAaEhyDw/DEfae224NuFGR7m2Q+1DcFyUoDu+dYj2tk355cb1JVDjStbTS
3oiNtRm3dGO33rH0OiM1BEOm2usu305K7Tihhwqf+yesJ8YjKTLCliNKTmwSDqV/MLfzai0ah735
dni6qyEGLeubDmXq4JCMWZnzaJejDzDCXmoNhNQr4JtVaRo50rfNVW9bk+DsdN5QSJJmgBFTkKxr
zzfs7SPCa8R96B+y44OmHV3/kGFrQ81Iy92NdNJcJ/XdpBPziJHd3x38/0K6SWFU3sWz8y6SmPMs
GilXemGsUpx5jannH2DPSYzTjpC6fzu8ZXWByYxz+5DiDSIASKIBYegs/J5Lp+MiHd3FJ0irB/Tk
9sLOBwolAy6qRrwJIFjpRwbkwAFyxaMmCJj/mhpHuhP89OTJSrXkdPY7YPORdW9kto+9GkKdeCQE
Kxu1kUMHo5zeigLZ4y1yo02k4/htI5f56fubqoJ1Sze8cxjDsiRZc84HnXijuIMJlKDIwrp0vLGz
0HIaIKz8xXB+2q1+1AxfUmc/VW8AF3CrAfHSy2a337yVtBYutpifSbe2aTWwx1VrVj/ZWfIh9Uxx
rwbgwPJn2CPNUP9lbjYXpUo6eUrWFWS05acVcLs14oagRj2X8QtPEX3stuvl6VpSZ2GzTlBugA45
fk3GcY95yTABsr3Dk2vKZ4PFeiZbTkouRbhY/Gs+FD9khSLXvFH2dfnGbqOg+0Q4+XXtF5Rabi1A
2qbJFvVsKyIENrToB6vcEKYmjoRH4fcSJ9BqiyD7/b9A5SN+P+1+58ba6Rwi8eUQQYghbTL8ttGf
TsWPNHhpd78hF5oaeRK1XagBVk97fn4I++CiRT+w/vruUOiFaXzYxg2hUyENiPuTARY+ZM4NK2If
hFIGiJJpaXx5h8xBTfRVKZgk6bJ/c4X5PZ+1Ggu82yW4u2oVL0n+B+/PDnPcQ9wNZfhC6bIXf5Ba
TrUqPAbFNHOWV74pmfqOlhH7RxmGEhbNykgFixvzBhWYUpX8jUflvkkV+zgjlHpCGdlLkYs9Uh9Q
10sbxS3TxcRTe/FiFRXa+hnpRZL+LMr1n4WNbcH/4FbbO61sq09vV5QuXDUqpBDN0YBmZgQp3o+9
CZpB77C5bEqXwcJdO7wMWjwyzJl09rYbnhaOWH+rKoxyGeHFJRbTZCWXf1ZzNyJf4W2ehcsb2oG6
6cs8VbG23YGloON5KUkYDsOgd3vSxr+0Ryc2P3/qxzgncfgPDLAKc6f2RziRolvPu2XpIkFL5d+6
0KAlVn5yqzC8UsOuinDyVHh00/ScIrlcobYOo/oHu8fNXcDb5+CV9W7lv/WzXYTe4wkUZua2oE+y
hthADevSga70QYmCPfs4RP9hrP7rFm3rN+whviCbAyJ88cKEhKvF2JXnftY61XPpeH2+ZTLcn03H
5EgrKAfXlGArt4pua6Soo8yESpDMbMeyfBesACoOBObrd+5Bta9k2jO+Gsic0iHNz73JDK9Dmcd2
7ziiMcGSAiImVjz+xL+jHNUaxsf5iaRU37NAQXZwkjaUPOBo4vpWF6Sh7SUrGM+iGqZm71nRmwWQ
30Wne2gVXZ/rQKXycolgtqR+uVjYijzYfGNilfxw39fFxXq2DciQJsUvQZh4rZ58EBL6mPFU9TRK
1t8Zen7AcPeIYjR+PLiZkTVZspDw4prdsSJO3SfToHIreCGTLGc+BRlcQJE6s8wT4BvGs7NcS5KE
2y1wjqkfyUVhxVKYaWBj+6hFQ4sLn/iVwod/CmyWZDmgZX/PK1mnCmecAT9P3rRBMxl1+fUaQbty
zE0o/OcOw9GA8MBCMrTvLTkoJv0Y+0bnCmGTne92a9FlyJ72OnVVkYp1JzjGlre18ueZev6S/bTo
fpNhziFs/ju1DbOQhD9rmqeDOnDcvtpDo37bZ3xr/ZcR9FG9GqDH9iXidICvb1UkmzPT1kVOfh6U
cnmckLDDI2DDSNwjPkAZASatYSJ7VAmVPbh4ZcqO0Kw0eY2N5vTFFymOru91+C6pDyv50wEbN9AC
rMX2KOaJ3ATvXp78sGrPqhw3yORhWHMoLL7glOH9dT6k0xYj1TVi2R6DJnwzckuvGOmoUUgakp93
dRcMLNfFAzqjpnplhvNNYLbrwPSX8AURrNdLFU9Ba4asWHg6Tg1TJKAL0i7jpzpbmlwnutv0ldej
t5GZWhnOk/Xk7kbPCieFml5zXpDwObOb8J3yUxbw2qNP+I/vudzfm/+SKaSQm6h1mIo7/dKh+wGI
lO0N/jYb/8Gr/liy220EJigN4RBEDuz19TqYZhIwdEs+2L7CoKcVLQqkRnUJ3Z1ChWNl1HQEdeZ2
VJfKJkJAFGiP/VcTuw0VoH1PDV5mmlMU27heKRrniAHb31hvcpOQqQC6diCeghh8poqlLndpI/pd
BuXcCq8Uj6d6Im6oxyhNS4J83ixkCwNFcRlHWHuEIIzVSVsX9Cry7kkIRq+y4Wp3Ihy2OkueAJpt
P/MxQujceE03q1HxKHDiHUPhQakxYHQiUU+BXOdvjgYyPjtq+6B3Ddcuna+06jscg23wMcSM9Cgv
FhSJjTRE0tgtOJ87uvLobMVdjzgam/VcHgjj9pJNY5pPRpp+SzpEsbXzsjbHBU711zNYsaAoHB/w
/SbqlfPzmiqMbenFRftyLbJ9/iwPoDnfILdx5KrpTlIJffQVW1MxGNP/VR7r3xdaAPVFDzt5+qNU
BXxCf4ECxwltoM4ocadxLIT1rrbckWrjmbvpyz2NTvlEKaWmWXM6wioPY6aWaOcZcOV2Guacv8NU
5qwhCoG4AheCa24wSCZSqtSI04Y/g78I5/neqNtUuuvjWz9RadaN5E53UlUcdjtTxGDrEEVCpGxj
+gRIjUWdFbCsXKqiTKeJdXR/eEgql4A68DfZ051uq4yTrOP7Yxm2LSpNKiWgrBNkeyvZhg2PqF7d
v07BEbis7Qv042a8PK7bDsUXZMf6Q0eZ4viEZzn29yISjwbzLXON0OsJreLjUxYczTY7bRute0gT
uawsN9LLaXYSHsJcFqdFIaLbd/nI8KtwTJcVwRF62JsjMG9skOemc+W9RyAb6c3j9FK2oV7NbJnl
xMis/sK05MyaiLreUHmrcHSroIfaMXvIGIBpUGiqaOdrgipvnaGE+By9PIB5TQaSvZGY9LuUHjjU
3q1dwQ+D4+COc8IJbiqpN+lKCP839VszH3U87BL/sVb/hoPAbxyhpQpVn7Nf1JmHPQ+J64xljrBK
klA1Q0kY4FQy5aJi6g4F+AS5vlrSjjvkBDaFlhSWeeFAaq0yjuAHPHNf3hwfA0sMEfgtyVryCiXt
KlzaB5DWjuEvbnPRRIU1Pg85A/3z3LWptV9tuEhTGG6FUWtQ2DQuz0WCzrRHkoDOTAMhnAgqTHZ1
U4Z+eEWt1h9n5jnWkMng72fr+CGJgz33tCoHJPfiOE1mhiSogjsft6wif9oU2LuIO26o1XF2+Jru
HWvJ9h10jaQX4Cqrxha0gOLYMvLPJmlaoRkhQvrJa2VJRXsaREKmH8iy7I/iQCQ7is92FD06HhvP
UFi4STd+wpTOfFy6RB9s0m8CFkPQVCla/VQV16H9ifrPPnViVTX4p+Nyrx4pZFzPeHHrbarUBWSm
szEwfVpJStAKOILPRoaLHzpMurO1wKdV/uafOy3PwmvIzG9432WxEfQDa6n2NcBliKlug3AHr50n
V/T9IF8euMBGJOx5s8Pv0XkyopWdkkAtGO4kYWfoRlx39xnD+bJk0cKaId1lHZ0stvVE5Ym5iWhv
fd0qQjlRImSOjxrRBuycF25XeewC1IpuLPcIYItEgzjhjB/cje+iotioCQD8EzyUanPgwyAMWERa
lRY86A8ZjcybZKLcqARqKzyX6hfIhgoDeeSjtBFxIRmwinLu4GpG2M5fuq0+u06fypKS5JS27TX1
mFGYRsvyEl/nUIh8J5UHQgFfn6eVzhm8ufU6mYiDd22yyeWs/d/ECu+rB+dghDVrO6iv54FDhDkJ
oBs66UTLVLC5dXWmJulEaMgrUF0QDHLA3Wo84TdMQuL1bUBxu0r3mNOqdsFGNDKu8/v0gK5e3b2y
bm0xFxJstkKlYtCZMTQza+wwbtJc2YJo8r/ait7cVOc/shKWjnRIGb3YyuzZrySoBQA53ZFQU1MP
o7IFrcjSN6dPzOzRV5IrpV6tVZfZokomr3gGaObXgVmP3G2D4Ie1oGqpBbp3LcxjBtxfawyRh4tc
RtP2KrGyrTOFHyfx6f82Zw0mmkP5n6ObbgkyegSNKrupYk60lV+bDKdbC3a8YPYxra5d0+qBAj9B
EhU2ItZGcrshl0PQWP+i4A3neKkY+v6+lr+mzL0t5mTDtk/+PWEpdI3XrIbMqjdGsUuZJqCLKA9m
P2BujS/jttobddgaklIr7uUr9ndM8DpRYTSzAyDjw+iyE7YX5s4nPKniXBlnnRu27I1c4InxhGcx
kuRYSCr2cClUIXgk0sK0qlvam+tRt0AO6ZDK3dCXU22TJvUdRJ3o51UO6WlGx4Y+DBUWHaWENNH4
nUaNEzd08n7+9nEdcG+cW5oH10miizi50qkcTSLOQAgyBKMHqqYBwkpgVr3WP0bHDpM7nLzSDzPB
8GPBfprusN2X0KnZwiHQezJZFJrzDPXh5EzbR4JdEL2s0eQ54W4pWRnxy20cagKAO90tHlop3aqI
i5EL5dFvv73tqMl45quUrLo/rmdH4DkOW3LQAcPXzJ+Jgn8Vw9IIgLXLiLF0zpBVsesvQAohG7zB
i+8sl7B+7ZOx0R/oAYpxWEXnnu9ZchlFBsfms7vNCfFE1Umd47lhiAkPVIJrR6azhmu3OaWnoE7N
GAwjq+sKL+TR+kmdLu+BwOQa95N5ZxwoQ0JSk2G+KmgnUAihXBQHRS2Xk/P4da/2F5LMRyVL3gfc
1/7LAhqoAUXaLs0/NJoMEXKzjXAee52EeNwWVKuOk+2X1BEvJzElOftL/9eFuHG/sBszR/U0pkM9
GOVCg1kw2jLgTpS5O5n0aHKawLC42eQfw63p4svHVVm9WMHEVni0+UeSM9Jv858gcA+7LVz3kDuh
d+42s4MQK183i+dki9JMEgUtz8cNiCn9ikS60bpIed/Eqk7vyTaSSNhrre786mjr4PIeihDuXS+b
unm0+wbEAddJZhDPQOiN2LuQ99kIyexTO0D0MfLpuQ5q85dFLDbG2UJk+J9qf/ZVdMz4CrWMpUCe
Z35pR7LI52s0aXXSZ0J66Vk+MchI2vDMzZxxkq8KGQyClPSFD8slpeRFh0KABM3N3iCfS9xaghjh
/fThWxomL8JarqtyWcI2KbIa8JwaWe+OiTAe5P4qvZI+g86SR1JQdQZZ7z7R3k28BgtHIO2j4OlZ
GTidenXpeKTLTd05rtK04CAy2fAeikvWw+EEuxlKTt8j+vA2EZbHzxlQTHEG+w7DlTvBzuIucfZG
AsxnUKRc7sSqJlpvowmggjntJlBcfvby6O1kMYQbcZHl/AdTQkzPoUmMBOz+mBJ31Yh+iqJkoyPv
Y5VegIB+14v8TpwggjVPcAQGFxekT+0v35dCatlTayMKF2px9+0S80n/0pr/5PdjrKcyjEGnnXcz
IGgnMQJcfce7dubkQU65w53WXV8+jmt9csrXH5+vJqbglOGgQ0EF06sV83r2XtNLgulJyVfJIjnh
x1w0ufYeKTkM6cNNAs3ICbmoOQknHEalUYbU75NbkFLyOKOEqkK15joGTA7bgieIRbebL0rBAR4g
1SIAWdJylXTTj4nhcDgvVZx5XKoG1waJBXSRhuIBWcQ6jrPrAFd1ykzBfspoBHyZ6H0z1POjNLBt
locqGYfsUezIOTbXnl3swKH1XnP4ZCdByqvw/bnbLb/ZzxWwTNXz/KL9ZiKQddwI4lCfpbqa7Pis
/5U3kQy/lC2iL1gRyGGHlJDS2quphhWsHX2Cjvn2+90LEasqE9OJw1kexx8cbNHtb2zKoraDPcK1
rqYo1sW5vVauCW2jjWDW0r8LvU0NcE/0iqONP3SpF6wv1jTedtccitfD7f1UDqRQ+qbiEJMWIG/3
OyY57aFjXIGkpIXii7Na/OmG3umfYg5SAQ0XEzaIe8OJ5X5Egg2yOCOaE5iOzmVykx84DVd9Gv9B
i2ESYLU2i1dVkhOMeJXR69xCU3NTn9vSFTRU4/9P/DX6CrMkJDoDI0xRVCntJMN27Iqvx+1qaVlo
MNpBoRaUWVQvjUJ+8/8Cs5f68VArDUEnNjGAcMOHEixneWh34rLw+cuSBM7iClGnV+5B0yPPTnlM
JpKmmpyKot/SAcex7q7uFF670ay6P9HXN8n3n5s93RJMgiavkuL8qzrkPEB14w8tDWuZe1hZd0mb
ZTM18V38Ym45bVYtoRM5IRW0FJCKRvKtXj8YH54dYsmRllbo64rAJ2Hv2UPSMv+GE0WYu6G5/a4N
z3RWKVuAP2PXVee8UuA9vPQADVJi7wt6eYj9Ir5DB8Wu2Yzn2h302mxFcfnendX1rVaWNO+Y/s7C
+ZUGMnjBAwoHIY3or+Y22VEjrNx80/NVFL4neRlx4qn5ryr6PPT0MoC+6XQDG79OX47oqCEmRXpR
DqMfgD2Xxd2JUXLIRX3n7IlnjG+z58LSQ9ydNdGPLp0D1TMMmPN0xwlF7omWQ9JD3Dt0UmFGt5jk
0MSfD4F70OuSW1wiqyYDkXiCk1S/DqvSptYWqQ+1pHqVZ/lluO/JmLsRcLXCW+ISo4tV30mU/ZsZ
lxBvGjlKMb3YQC0JLiz+mb3atYwsPBGZXP0GHxieTorua3cVlDC7NEYMMLkQuk5uo5YuKg/bXxyp
BbF7/l5M7618aRIrVCmeSos4oq3W4Qlf268tFe1NdJkR9/dAmKw+TBi5D00nTG8yK7uHfLX1LCaf
IiQjQFMeXdRHq7k+DW7sCFBtMMOymi7uQIqEvak/xMrxCeyS6ouY8TpWuhuR9kZF/jaKgScEwTDj
whDVlSrVOJZw6WTqO3ch44k61t78TRnVat6WUG3AnhgMnEPQqt26Hg7wZhp4ci3+bXKjPQFz9jWk
QawmWEeXWc4oZMByE5FNl6uFf8nz7lz9mBydDNUSUbUB5KGXb/IBpViHBydaaPzSOJbaeY463e2L
Q1vZk8wFAjtp7ALGKeJJqcnlj0nrGYHT3HniRYWYTXSg428tnuimSyyLxjVQrXOU0HfWUnXXD22z
wgCM4txFTPs+R0v1GyKZbZt0xD42Ja9SU/eKHRW6SafTGXsHtH14ZbKzxTIsO8Vh8piDwLFOUzvC
insoCkjLFds75DKgkWm5kk9lwIPXAPA151BVgqOMlq6pWauH0rpTZZw/pWpqesd8QhZ5K5/LpxqX
dadT5avkc7rrUJrf8riO6wnIEVbCSheeXcmzG5GU4DAqLTlXhn05Vusm5w3PF2IEM2gXT8HQRWFN
SBUdBFGzn9TiwnuxVRdzIf4adW9ZA5Nn6cWJns6gJf6XBI3hG/NM91pZ0W6tSGVlOMnSKYuRzv/4
RyaIFgKK5LBqdVpWxNBAADWLXDeHz3QwoFtstOXJVRinHxhz2aQ6eY6iYkR6qYmaNOwQxI+hmWuN
RODhB2Bcs66RJTbu1fBlYWM1gb6YwmAgDDmHe2yVGedj0zBWFoHWjFs/iq/qoxCKlOvRaYZeXbS9
dsjZd2mp7iYvjztsz5Hb0wpm4inarcAWUNffhb0zZivwJFdwDOJCX7aXXiCGtGZXlYir0VgNjZoo
Y1uSkGD6zIRQbBzABvts/cMbI8x3J1W5VRvOuILnhwWVKJ5+1/9pEc9qZh7/BvXkzBw+zCvrkTAV
z4aONtCYBNSTYut0Sm4RmJWcOzlHHLtp7LApecCZYLrmNZdVmBHT8fmt5++gx6vyQspW6Ja2wAOj
sOFgOeBaos+aWYMCS/aUtHclvamXvQ9tySvXHL9WEjuKIKKxDip5wux4LuvRbi1LRWk2+fI2PuuX
4MkfeMCz9ICuYqmD87T+cfYRh6QpxIXroTC7e6J8MbMjg9k0jqCc5p34pTsCF0sbbYmy80QZVyIk
Ts2SNSSUzLoSUr/5pvtr4p+Yk6Z0hIyiRe2ciNQDWGgNMQg3FlQuOx+myIf41NGWJSIvBHdDudH7
dQkecGG4+nOvN9cOphh3Jj1RUkvsZ8wScMuPurFUjWDIXuLZLTUySVEmGgGxpB6W7YXMBBN8ID9p
P2EQdPFmywI14UruqD3AnGVtu5oALM5NdzlVD3qOf8wTiVKjx32dBNrmAgJUkYIhgvLQ4lpn/IL5
JpuxYCgPm6hRIpm6Y9RDTYaBWxhxqnj1RZ2iDGMF665b8wLhbh+Jbsk5sk1Nddwox4Zs9No8QFmk
GKYs7H1cDCoj97RA/gGoA2w5SYszt3mriVIUMFIbwSFGwyLVgMyzt+GcbsGcaU1RjMg/98AvuKQF
BB+reoc1uTiREZpiiDBj0J7U+jWq6tkS0JyFyHEn7KGgQ8POTbrzO3Gr8/R0+m8Yjq8S4rzUwiTq
+IiHlxOm7XlNnKwLVYxamg5pQ46YmRRU4QkIV19nIcC8jynMtY23XZ/aZV+eB+mJ/Zi/Seh3/q0e
u77rCbQvvN8gvdp3VMV4Oe0rm0n87+aPEFs3IxicPYYOBo/of8kgSOtab54iwZjfJVzeUAfEUek+
ZPph7p+zNFQFErgeEwH8E755K8YcaaY/MPKpEr3EV1ABjTd5vd5bSp7wydK9qgE+d7DGbjlk60B1
trmLZzsOKAD7mP48teMoGPwpCNplsCrC9Y+eDU970MnENnM8FNppWvcA9X8RVePRw9yYs1CKKtqt
650PlBG2TKzMysmKrmE0e4TQmg6thAsYvQ2CYtQKqPpRQpPb6hyXBO/cvPvsHpFmYaYUjtyZJ/lQ
sfI9c8N+kOU43jt+d6yxVc+MUqr0a512GNqNgXffg/pw0PSgHDBlFzn/qoyzJWutcUZiAO2RZ+wP
xpyk3O2BjfLwJiXJG01QfCk2Mw7TzzzxzOtIcJqq5mnWytOlEoRHgKl77hCEe9NQ9VFVM47Z8x9/
bfUZT7uOYUrQFHpl0PFio4RNzMKSvVqdsWdgEIYZx7SGcaop3fmdjXxSuBeEykmRkXQGBl+sPrVs
oy48HXe1HMtPAcPq20lcg/DT4pM13gaPng2es6QlIz776ihToCAvi21HsUhd9RRpmgWQytEjQGfP
T/cwqqgHHgIWptT7L0K+kSfLM1p3Dt2q9uZYtycVV/1WiwGn4jTMdqk1sjMSeSZibNM8M1tKHHjM
dfsHbwcJFtLqk566ZDabaDCVvE3lR+l6Ti3AJpq4UoszgiQQZK7NN2ZipVLrwwpQ/YGOc8Rz1pIO
+8/dByhO760XYa2XhZUvXDpChEKgGfi8+xqxSDtWsmhiMAYN1him3fWAH2oSwwub19Qlqi829qGl
btRnP/MU/ASFIWOY5IRVXFRdR5J5T4yIDeR8lleHqwsZ2ItVyL2CipqBZfsfPFpYFNSbiZ1I3iG1
s4l6r4Dv0GNm9IwDaZXTn09DCDVagRn5ViZpNqUUQ9+gVixkMX758mc4IbgL4ImJMdV4MzxU5OTL
lWRSLFT/ya5Vy/bzSL9wUnevSb62ta/r3fzg8sdlGDuO3k87WJADUlYN7im+s7nL2gRIm+rZ92ei
BtgiQbbTHqG4wWEZk1v8Eg5CS7+I9fSNWsg4nWXFDEUXdIKzW2VVLTCOsPCoN2P0W7hYZRe8V+cu
qmb2KOJAMFGlT7FnvvcWMLMScaQt7KaxXwqb+PjHUaG6vx7YHebAwcjchA6ob+9qTSROluv4OIjh
WvtiOk/h050WM0bB/Zj6fpzSuBm+4tnxc3gL4093YVHDzuO1OEmsjBCGs4W0ymj2Vi4Gn0Ev5HMw
4lDWSHnr/NTSuFQJsR3/8b0wOybMdGiMAFOkCk3IUxM1ZzXX8k/7CeOKmTAS+LwLkYbCfPpqvcDQ
MOpPTj8qlWYwKg4Gt1K6DmkPu25eL0XA+zCWTjsTI8NGGG11zC3lBQK/qhGvC/6tHoBF8DkKFl+N
nITuwTHc8ey5TsiBCZVm3Sq1dkGOBZdh2isusJXtr+kxSJSG9Op3qqd4BrgeynI05h9A4bmrzJWt
OZtSeo8uDYPIuYkcRayeEFw6oGhUMztyIY/AiVU8wtlSS2ZHkuzYSJBXzOsAUVdwGbpQeXCFQAOD
I/NL4jEZplDwqUGnTgwCNEILS959ozmAEBPA5gzWKOGeLyDfVS7J0V6cf4VLToK5JJqfURTBrT8/
bgT2Yw2Wr+hGaj4KWzcs9AFbBobjixl4kaN8bFfr3XEIHAFzn39Rr1Q75pvOLT5/+iWhcI/9SKLt
lcjHFzhWDjGNtGe/U/6+nM7/4ZezVr8Y7vC+57rcF33tlMA9JseHyqB1hZo1CGmWWyyFBGztLvVS
g27dYPkHDmi6BS+W+XvHoOkQBDXIUXGLvmnJdqVSj5fahtd6Tyl2U2M526yVzcJ97CzvY+xK9h2m
jifWr6kHqqoSzlTckTk3me24GMuKSGLyiV501xSgsijwXOWJakmxmFx0hnjC++8WG9UOmw6KvlqO
VhaWRKxmNkO6IL+byAXlRuc8AsWL2hY4FH3QD1KBw/pscHZoQltx27qYNAX5AMwaJv6CMruEAHuX
abW+664WFoKEslSCMdUlwXogvDJg7qsFOBhi/hGVRHyez9SaY/1ysMz+oTu2v0p4lruDEGGW5wNg
VS8ZT0JPn4p+AtSCDWFt6t9IQ10L6Ppl/klQugc+qwcszqrec52SlnnA5N88IFhsl4CgMl0kBm/M
5gZTmoXZ6fSw7pWselOk1DuqORmvCA/ikiZ/1+UlEXbNvoropF0nDg+9J6EtxvQ5NlSM4FrBivg9
KxpbLJl/pREPRUuKdE38A1DHmoElrsJxNw0sz2OD0FnVvlVexEFkkUSQ7HQ0QDo02HMammiuGQNS
PkFXCakES9Cd3kD0r/n25znEKXUuqnxciRvDmV3/0LXS9C1nVq+BTvuU9REz+IXFtb11Rq4hu4HF
JKpppluKfCqYpppHZiGEw0A/hZ1yy9pgkyfd2RZnNUtzGCghxhjvXWE0m0bTwtLRGuoxHu1oUUIr
AMME8C9Yund23XGHkgLGLKsVP+B5JrMo0Q7UXrpQ7kkhUpiDMc7nuu6YdHvL6rOHefxnW1/hrKYr
80iMJsx0H07RqtgSUtqj2zUlT/pRjn7PQCQHYuLeoPb44DfNwdsrq0b4qXrjZDf8NJCcpnC69ovY
wKpDJDRIp43erHhvWW3GC1X1w39x12lmGF7pAx7x01B0WdY9lnBmBbbVje5e19zkiw+s/WODypWr
+YslUPJLitpZ47YsfISjJkOy1hd3noHNHPPFVYVwe8MCmyNKikHRfCW+s5fQ+EA35L/qCTAoB9+Z
w7tN/pNq3cwNXpV0thKpgb5AcjEl/B/HxSfz9vHMCce5f9b10zaMVu8YlQik2VTPWUo5L/2OleUd
TsJyhR95RfCv3K/Ize0L8j3ai3niZj05oCHffxVE8o/ney8WMJ4ZxEdNXtqenHHtE4KfWWORX9q7
wTSfaxfXoLOy1MYjRcc/Y7aGcx+6oRbcE0oma+EauAQeeuYEKiETE9K+y/uT2PNBEM+1AcfneKkh
KZ+PAe0xQ4/e+4xnVWGsKgdFaZBBv/iRQJYFWat36JKK30gclB/3S1/opgPn2KFTDyv3DIC2dZGc
yLkM1eg08pormE34+ohhMeCueipX73qo6VVk1fHc6ovbYC//hx7ZQ6UJ7kulKhAeQ56/glwk7FnV
b8ZD8aQIP/p+v2xcg9b5odQPcyi6rMrnnQBzTqU6j3uK6tNTBwSvJrh7s8o/Gh9ZxwXvyOj8xd4f
xj18b6IExsxql80Iv3lnc3ZcNNfn0/IMEAmhNvhsrcH0gDGsxj5FxEASMUHNl5jBSusrwYCulKCb
WA0CaESm5LUzadtaAvZjyUsoWCGrLDxnXhDuj0cXXrDkeNa5WGqKcmkWfi4882DAJYtPfqFQe265
/kj+mq3B/ZIhyH6FCJMDmRBcjg+iBOuMRD5nFZtMKadciPVmOdeFexCxfHCF6wZek5PkXDkBV5Gm
ET0LdSwWT1DfRr0tCMFqdbNaoYdVlK1kDuFNisRCKspUmPWy8+rDn9GYZZcuQcepx0GXDAHKzHTu
UqCVe1TpOSIuayNgg0DCh3RoVz1QEeE+MgW5p0PineUArlw2T5QzWXw0/vXFFuTALNdR06hX5REK
Bdlrm1+rUDm4jGYy0P02kN0UlnfhNmTFwmdnbAqefn+jmGDdR5KeFYcjMPZs2W7VZT1HHEERkQvp
8CTBMwG2Ojo7Kcb01pY3xAoPwV02h3GNVaRZ+B2A3UnPOjJ23xFeI9EZ1Jx9C5bZHRmuH6toWX2f
2eoeXRMWMJ6XDTiOZLap4d3hbW2EKkzQGNX4v4AxIaf8OI50kXvcoMNjAv7P0v8thpqJXJAT7qKV
/xvxgzwnawQ8IK3GgfDVHSo2i9NiQfqUM+PR3Ia3WwvU2myR3QMB0MlNrvQ9Ixd7vspjHBeVYEOf
LQOdUqLDDWfqepDfmbsHuZHdbs/guybMYRJ3tIYN8eQ7dkECz4YXCUPlP/af0pY89pHNMVn+tMm8
cJuxlG8p7dtZZZIskMFG5rAw1cu18sj2/B6W+AEnw9DgQG5YMElMmDW1ulSviA/Nf0tfRPb6y69V
daHrCgkImbVErD8HviFXrVCm+F70mE/BB0mFD8zyzEwycAhSXCgEZjsoqOnEPAuQfe2bEYvXH96T
jIwnGZuQvRxmmFc0VarT179T8wceoJVJ92iYB82Rn8zWO4McN7sxbqatCCeS4NJHX944vZGjiq5w
7GD3WC5xdeSr7YLXASW4kz1kSb0LrYwFY0B9Qq56hqi63MFGYt1W8aiiiF90/DvY/KO0TyRynGJJ
/gznXl/9saVnwB+32YX6oiLirQDIF5tZ0dcgu8KWkLNbIR5A6z1NAacNr4CgfXmqI4Znle4HOyga
jhrKh3Q+obCEInGVPXaeDmVCEXrRsfgWkouhtWHGPtbISUwwjx/kuPYwU3PUEah0Jdz//Xqvf5L7
7ribBgg3tbBYhkCkfBf7vlmUSkqV3NF61hn6muupB1XoptX1maKlE5jLOn770WYGK73t2bEnuIdN
8hsV85hXYsO3x8ARuNA9c8PdzOfH8L20iMlb4MuGXm+LcI2OYX3pQVdRPxDqLK5OCxDp5Nr2Fl6x
r1MJ84TmoCCrYXhESIr/f3P/OVYwmnv9GxHEsae//3F7t8jHB176u90Qs3EoUSOOgWJzpVgdFGQA
x1ahA3kB+C4I+SXdioeHNimLtftie5DQO+MwVOGoxC4mlkZ5DxEFevO4j5/G3BXHAlpD4ZMjIkzM
fx8+/X2LSfxhL9mdZuFLaXU8L0SgBNqHZDQvtaGjggma2gTjjJi+L5b+/IA3pwVxl17rTdV+slj1
XpkzuGG0icX3yqyMFl2DGJJSkTSXH2+Hnb3QOH/13lpmtWxfyLDjhlpSR768lsxBODINfB0JxOik
wh3jA2a2uLkNkylVS9xyux7Uq3uG642wzOAld0V9qS2wzfVvKmo8Y6rktPaIVyWMarXGjc1iP+mc
YkZKGm9dl218CBJzl2fUYFh27ccPLoRVGVu8IV4SLzWBaq0M/pU03BRZBqWjfoJQP8+8PBg9uuFk
c5Nwhj9NyXaNlfar9fyDsQrgfxVd6lrcKkDizBcWrbIrrlQ2kBymBuy069JBq1S/JUiEqpJFw6gp
fsWHZol0xtqioohZQo1QKZZYhMPyKWyE9Q+A+JKVUO1BvVg/IGxGkNxMLkhd5kXY+nWmuYASnfpR
fn9lnCUa6vhXwEEbkAJ7H7RSldIkRp07sh+ZPphqoAdKLGCNlV0cfxNzUxI9scT6lhJYN0q1paf2
DV0brJLyIu66rFCaQYBREcuC4PQYhc40FYI6nKVycL8l2WF7+VRHLrkZm2t36rQgT1dIi6Aza8La
RjPqrsCsVlZY6tJmS7N+Td/6XpSLx94e+4yL+zVSMXt/2c98hZuHHYQEzTkzBOI8ln07kjUDLU42
Bfh0ERkk65YYGK6dVFI4rOwMwm8CMc2ciDLk+/2TXoEqUGFRo/UEW2hYAn2ZYfXPdd+WEHKnxYEf
s++BKNmEZw3WD3TEOoPj5LOWCxjDJMjbFH/oV+lLMgjlH+u0gblwmbh+tvb6m7Y1quXktpxFWf2h
qBVxEdxG5lXc9MQtdyKwgLl4nwm0iLt2j+hqirol/4CAtrS5neJZfxnqj7bQIqKWfEFMHobyX/pz
ZdSkAnh1qrCTdU/HCUXzf8yFyv6+HioNlzPIoHJnnC3hkikv6Ssj4k5C7E6cLv31QZ5BJf9o5KZT
i2PbyDIZcgul2P+gNNpe/R3swsCOMT4F34gb3WdFc0gTraDAHH03sn83M1IaH67Tzn9H1tBenq/Y
/lhC8slUcuPhG8Q29ho1pokPter1V4RIotjSErtphas/lGYXOYHyEbz8GkecM5xqlAS8jC2SoV7P
ygPo88m3ZRLLRqSKhOOob03XoX6d+5/1bRYezMqTwGTksSC/OZiyA3AtfaNDIOUAbbcuNv9xRYhd
GLDmuvzHqqulAby+Nf74pP8FkNO1Fiv4ml91sfRCZsHxtr/C4T8p5LYLh6KWNOjW+w2Z5RZ5xIFY
TbxZrg7GFexWjrrEPVNa+UbJ0VYlKYIm31uIHOf+Qr7r6oSVjtqVKxk/BaKimYI/3DzNMOghY6aq
zPE4jH//idLrLTNiC/CMS9FzbsTWlYzbN+oyKCo5jU1og+Bm71LOH7BWn0n9J6ybEozYgNPiQZq3
oXZJrDaNjXQV0/C9KNgD/of3tW6V/OYQmif4XWcRMYMhlWGDBRzWQzv9GMggYpzNOMI3KWc2VRaj
rZveVwaKQ/CSUQzNE8+Z4D9/JSLix1eVVGj/C1IUTtHNb2ijz8F70z0okfz4tODhzbw72B3VdHQi
KqB+W1zf2P2FSisjXmo1u4roQHvLXg3Z1J/MJZJwZYSd7cWry4AIDU04w5cSKUkVymkVBgzajfAQ
w01zmkXXd85RQzDol6Y23/L/n6guu6EVa3+AOuC10xOgAbo7byE+7Yw9maeltnZlSFWEeO8D3bDt
lq4qAXvfFPc8KU3AZfwnpPI/VpAOIXPc3YYFcNSUpPeoI1UV+ZKjqtpCV/0JhDlOg9Qq9VNru/L0
Y6rxmAFpbFV7c4qiw14dVrfWedPfb6dYzvIos+pPhzjrYhnm8x/Q00jZ8ko3zvu8iM7uxlRSA3og
5d5ouP2ty9bby1eBs54QDwYa9wGYkJ5V4xVw3SPREBCX+HW0Z7xcThIHvFbFjEGv8EcaXDty+5tw
+en3fNzkSyanl5sHQsxoDeWfX/ZEkzxHgKq2LR80MARcwVImFytWPltRhcddgMTRrn0mzB0ZgjL3
TRdO+LMdjVLZAyXuPSXQqzgCzZeeXn7VV6kPNJLaM/Je3bMK5AClU/6U7ijHXOXyQw64Pj2uJMWE
UdOfNUIjgRsMoLQYvGtLUqQ6IKXIOHGWukx/b8Xs+HwbPYQ4G6pQKJ/Mzi4lAvU5of06tqqbOWpZ
7ZNZNaZtO0m7SMrhcGvb9JieotIDTzn7isRV7aL1LlZXE1uWIeE+iqhv0jxFvLoFH/ZPmweAHuMe
lskK2+iLpI+h69xPyF5Hg1qp9pWvZt749WBNv+RjJSvAoKX9M/2z+yO57aDhevJyZMawWfXQbUv/
RKVAr82K8TsppivnEX7sUQ0MIlF8ap7oud/w6VZlXccOxoE2vTsX68hoUThXYfk1uJDeYeaEqXnb
WxW6rz81nPP3ecF/I3iUURZoLytL5nRMZ0ibEJa3qqfgYC3a4U5PFEU2suaC44EsDzD3m2cAvnNr
E9F8JIHA4F56id+1uN04W/UG9wg60U0STrNTt1nhOtLmKGcdfysZmm/o2DFk7eYLsUxsHnekRNwn
IDuhhJ9wteeG+yv9n+AYgpA2dGRIGIihArn0+WeXEvZ7zR+PqL2s6bvpqp442UcuiyvyI7/ra5I7
j3ze0dj7GoVRxKYFcaEZ9KsLgYoH4p3Al9b3oNaQz9jW9SD70/tv3StaxS0kgYhmh5+9rSzUt3jC
3/W91FgEKRNLyzaDl52DSasXNFfHUiYurNKbT7IwzQzB8w2mw1JB+neFsA+B6pBE3sNehbPKBTYn
y6SDunIzKF730hrnkwIsRvTQueLQ2Fb+j5tS28ZufXdmI95RRTAH0qY4ghUB07dD1aHv7By9D8w6
xGXQChRDqpf1Ot/BXO3NIiI6MtzC9omFAN+wbtcJmDF481ioygDM8XvmwiEUzt1zVsBUxEW08pwG
MjVgMKV6ZCElzatiII+/ymOhw4z8QeqbUwJCBZ5NsupYArP/WUssji+INU21I1eDjkh66hMmzHoE
eci0K71H6wGRmMZlk6dtPAw+Gg/HOZOfFJzTjwydy/EWSR+76ouzebttYicR1pxnSb40XBNGaqMS
oqDMEWVFK3S7eFY/u2kDelq2sKyOteP3t8CkOFU3BJCe5r1p3OLQ8fIDehrFVoJxj8baRghbYCPY
8i2GXsSlLzUjvQxk5SFGC25If/VOxzIE3EmBTSW9s6ot02oLJk3bJtYOlKMrREdQsaitDiexMmi5
YhkIHL5cUPQZDbjNKIbeNnel0i2dkd695S3FMpXzqsxRRBn9uWh94bjOcN1hKThDD1gqa2x0pJcl
4Qn23S/MQ7335hKQ+c90BUrATwj/P3rFCxoLp0WpEp8QIqOWtFT0wcYSEljOR0mkDxvesjIRLc4w
WBZ1+qDaC4omL7Y5Z5HccyJ5jbXnQFWI8j0PEAd8vQxpgJKU6hBafx+l5QozXw27FvMloC4h9uuP
hwpmVQZz51+4TpyHAtjh1nfOKxGsNT32tMvy8UatmMm8z3IUTMgNcCzQgfyKGNVcYUZJoup+MJCl
Lep1TTXJYY1BMwczcJ+TdVD/hco/cOuOSFUWd73+slekDXYFSFcDeN2NwnXZLXSnX5Kip0i+DKgg
Qhwld0LTHVpEalNxQgDLUyiYMy03F0LxMPaV3o3AlyZK5CMoDTCmXh8AlDXt0c+nwHzst4R1sEeV
mHt7A+qBHuKQcXndCPLYQXmM86tQzEY+Zz7zMehiV/l4uxPTspPYqD8GhsNzcKJuq5qzOoTv2HPi
W9Ot1RISrUPpHAlNB2BMOmztIlVvcsnxK6TRYOn/+IljORELFzSxXasNumldRE4JEM3GUdtIgTMT
Ns2+E006728gwZFmgcntoY8yMmzEZ+QNRHhpunlt1tF0bpfwoA1/Aa25faYXjqU3VgMok65lyD/r
gZYOl+DJvQpPYq546++dhW/25Wc3bDvTDwnSXul21QueSUUaZjJ9M2GwzKaxKrFmhrpZb++tORLF
5+Rbx7xujqwHpXu6QZ4d8ApS3jYxt6t3UVRMbZfq0pq1MmQSlW1Uq4V/Uhrncy9lELC2gsW6FeCJ
FbWUAyisd8RYyiizp2htpIPmcybSMkjVVLR1+kp3FAR/csbQQuZ+8iXlMnPoobHKiba86M8Rm/Lr
89o6s5ti5kQg2x42TzZ4nSB2bqvtfrnze6qiZ+OyjdfzqD+hbyCfES4FslGVHmFXF90N+NUkeVVJ
Ph2/o0Ee8fDOTO+M8tfvvnDD2CHjKc2OOPjJwj39b9d4rbnxoGaQkwFTBdPjykKnPWkI4iH+Kt+w
kH1s1A/rm1WhXj6fZ0BFDp3pC/9wLnu4FTGHs6A9Sip28LGSjjuTRH3ER7idjcCsf1Mg5vpUPIbW
A4zSNwizIByEDiSQV57Sn7uDRtNjZ9x0hKrDrb8Ys9DU6ooU8tbQzL04l8gtNO51CJaICXiu5DRu
PBboBcRHnvpOkQzJ9fMFfwT7Z23ABwYFE+VcJ2vjVUWBqEQ1D3PAxkWWoCRJZZ7C+JFfR2Zx+SM+
BmuHh8TXUpE/mqFcWIDGWHS+LL1GHWyi3Ke058H+hJhi0PgjhEqxH8I3270L5Oa8njKuXVfF9Zzj
Nd8mwCkefdhpKLAqAeYflqAoKw0t0WZN57mR9++dKqCkzdXHUGbJQIcSu/iZ118ACBTSiiMVnvVR
HcbdHvGETwQdBtFS2vHAWekPWOCxfHg1JNEBM+IurmyefnCsWOhWjGxlIjHzQyfMciRUd+1DSg2A
iyE660sVK6C+GQzrtTnLbi+5GXfOoRvBZtE6S934xH+O64Qnybv6wZNZra8dqKHancpYx0nj+5zv
ORgJo9Zhb+vH7bbKWZjSgqjagikvyl1WpWAYKEJbm9EFJBk1AK3GGFv+lMT+8WWa5mAfNhQ3fV5e
FAy3u9/KB0eFmP9H7Yh+cOtbgjSkBFINTcbbKHgdd1B11YBe2AVttwfySrpIjTMtnPppRwmKi2r+
+9PG3sB1j4hja9jMPwhnckvSvYbSNBUpT1gJAb32WwdrYLrJThwRgyNFqJEVw37Wa22PMwgq4kwj
JYiEqwNl0k7amvI/4B8i4qSnMr/dWSGAWDfje6Qa8lmFYQpso8ZkFyZNBs70LIqBsz7KDKcjjPHP
MK4K09btLT5MvDN1QzhTFceIS5jnTdDeCaQY9pH1HJnHSSFafr+cT8C/JryCW+N+Iyw5sR0PVppl
AsJ4euAyuejPA+b2yT4utyDYl6tM/x1vV8qsU0Hh1Q4mkTN8/18NCroml5D3D3jA03NU3eL9r1w2
4pdnAY3faHs4Jac9orrXLRioCbcmrSM1iuQVn6wlkgKBqPiNAtw5iVyBMudSrogvP89snvK/w7Ap
Lc2E2Tdnnz5ZGGbyW5JcE/ViIwoC0kY5x8HLaPLDX/vUyOtO688HiTChpqvTtEjD7N4nENdXECvY
nF4NuaaMFR5/moPJ0KY15k3ci6jqYv1Fg3za6DCTjCVqlhIsfuLNMyUlE93Namd0mTogMgw0DQpV
P4sZtXWp32VZMTv589BhB8A0yZet/bvJ53SpEOsGDTqNPb2R8slAYrKhaAHJdcRWrd8xUPcNoMIT
aEHvv2zRRSH1fdqFPY3mBUg2W91aC9RpCdNSofRTSYvzr3Q8IyDVicZka+2ZTMeXvK+arBf81EzC
LOdiMz5Zh93YZ9YGkZCx390rJhnqv9BKhBelV5Mq9V4OHhHBUqY1OMKEGy+UtqBra3e4Gq7Ti/g6
XoMgZmzKqvPuDZqY7PDQiurENPsUueU1sCgzAzzXAIvYXYgC+oVbJy61l8BX33X9uquYwU5Fr29i
v4FIMc7oTL6g/o+xOV4hXDQDkgz9Y/yHKn50MVXnjccZFfWO92GGFb+bLG4XtQc7I+6MTGSDUh/+
Z2pvaZ1k1QOSzmryx35QbfOJn6F/VdwHw27lIy4B1th0QQ7MBnZFWKC6g8jd0L540nb3Ljv+wTdd
cI4olFGDQ/M0b4wbrxdAzvF4ShgSYl+zsfi3SXy1oj7JsuswKkOWVlDyv2vPpqJZo6vCYkrswbcF
LEIYsHupssDatQ/Knt6yD6maI2+lr7X0sEITA0X9J0tc4LUUpFLTaI7MI+/B3geDJYy5fSW+yPH5
xnknInmeZt18x6omJwJHJ6PGIRtwHR1vgx6jlw4ZJ3WrfW+CQ2fP6cLpOQzMoz/fh6xKF3kTzP8J
PbZ/B6gwIq51Q570y4IuBqdRpKE6xyGMEsOXyp9yzPWyHquyCvK6BhRZSY3Tix+XMFbx/ceCuN+I
wPYm4A0/GlRqaazWdYoQZw14b2cAvR6Cpn+uRBEDDHjMG9bNWE+y7kUG4Mh9kGaISb/QUbDq/giP
kLtaNZDqR+DdZEh+rI8m3jrWH5GS++RwOxNWDJ4cthH0+vk3mF/V7g6TfaGwMlWk76RLVg4ErgN2
uVoaUhXfR+E3M8TAm8KKBj3lQLqoCSmO2CfIOoOC0uJInpNGFZM5XyLqQkegUT22XMG8/FF1bOBq
xM3O5HKPaynxlLOaWJTE6/xAIkF9FgJNSJ9H8YPRTYGmP0gvkifBlOtzb3emy+ORf8OsN6puA62D
Y27906RHV+UVHsABhz/ja8LGlKqONAsVyugxcS6r8n2ZthhvWuvWpzlGXI1YrM0r/bKGdN05I9AT
PvQZDfXVSpGxTvKELVpQV5bmJ1W+fwo+0zQQq3KMzLp6lo3ukVeeprWsmIkcQaep4s7qqH9/NDVQ
+KmUVIdI0+f43i+0XD9ZxG9ozkje4BBXjoXljm9ULCCarQvvsT18qHpTd9ansv76VpMIKGMoZcgf
/Ddz4V6CEQXKZW2T0mGvQWP7gTg5uwW6LbDlzba3qCZTCbVK3nQY4THjDwIofqcuXX2L7ebWI4yZ
PxbdJEjDTZVyl2lfoqyQZ8vOpHwwqWy4NJ1EUuNqNDaOts/gMGGjDEnMRoGChd0weGA02zI78l6K
W5uuP/pZNsD2lDTT5ojzD0S/2xKmAj323YbZmcNZkMuznHXvQ8qV0XhXdyCBnuY6No7Gmyh48ucQ
kDFbVy96aKWRqpiRlKszfA3KRvtarhn6aufvZme+ahJYhPBqsVoR5zOZ2hGFq0aBdAqn2BqCbUH/
h1NOaSPSryS3YzPJJFPxO0Q4E0Zw5MDDVBx0yXs7iCaKnEO/CrfOY2TmLWGJtmserPn2zcncVVu4
kT4SLZ+qFp4F3JP/Wh2rBPb71+BXKa/fUTun41THPJ6X7247Goa/bwkEP0xat2FqowmwCQ2Ew1bU
G4fm+zs2xuzDHKxUcEmILdi0XnXD7FJJ68bN7kSZyZxdf0s7dYG14d2vWt/3A7Tct0LJk7uypViK
euTKpVpKuF0G8rk3tuP0fsyK/BYdr3T1wlHD8cGczOae43XYpw2LtsycKIkpkaXIhAW1nvhqFOli
vSwuvJ1o5yUu9a+0q3N6ZRIpdNlGGLh8l8JCHomD0KBJZKjBYt959TCqBtaHgsrAhwUzA80ShaSX
lVqwWnhd11P+zVB8A4M+8pm3J9FMnD2XXysf/H4H1AmKlI7jesFeggpL+nKRQ5FaMLEX+yDsXw0I
gPKwdWQ/Tmo8W0zEIlZf8OOnT9qYZLJrNP8EhsjvRmYgX9/18WqMuI1RGvwPGpvcmy/F4ikmfAF5
M2whHQxPTBQN+vI0bqRCsDmJIMrRqno/C4sml70eSMtQffjUUfnVQunWoszpNBpUfJHTalwZ/a6U
ZpWPCwe4yXhACc2bciFhJD+HrdRIPmq7hxP2xD+sBpsUk4okKUKXnAOpFLAXOPODn2vmz+CPHVvy
gn+tTanlVskqcMojTnMYpkR58Ay/53jWsnycB90rQNkVn17lRwsDIS+thI/Vu5rdz24SO5n/9OF7
iEeE/lg3BIxTv54HVsHs+0zLh4EkgCPCQerP1rgeC+ERzFR9K80bHCfMr2H+4ntijYkvX/dER3Bm
HYRKlyAohQNLnZ19wrNCZQdw5vaTuXLwB93kz7VFMB/qoH3nGfn3P72D3Lvz4Tiq/IBAnLThsMrk
1YHQ74WrxiLaXYhCGqF2tg89U1TiG9k6Tpczy8JEam4r4JhhFr78kVE8i6aQgBTdHL0y9gg6mhif
8w4Ed6a1JIwLZDFRhV99zFCUVT7MUElSWdpU1n7xQLHHr+sG0xyQO9DMM1pQDkeEiAf/ovtYkrcx
7gZeUv/aAzzlChxqE3xNsHpuQJH5F/JfW6kysez/L8en6amPrR7HTkndXzfC4SKnEftf57q3ebeu
/OL5f3xTOkdv6vW/esr+b8j/o/RtVRZRJxehRm029qA0+UAOhrNrRPqTc2iISx/4vhCF5FZGBHlA
Ot0dJdM0Lm/bF6f8BPff0TsnhG9QR51I102b5PNnSzzzMPRJZzhQhbBh+zzZx4VadlP5BW4n5YU5
M9Y9Vb7wLg/iDDc2Hi4dqPR97/WSyfHmSidSfsNG1RauOtbCYZVjnAgZYPvF6k3Naxts0kTO3bKY
WEoQHbUo7WhPr/+AxGdg59pjbzKMaRz6+z99sYF7661fCS0i0Mp3MqI3GXf+NkGG0hYar0Pw795P
OmnkIhll9P4cZRmAVKu7FNR8XxVQ1ygBKocsxuAOspLYhMr2ZSHZ/reBZC+AbtKngvRFy+Fj338Q
MBDwGG3XBwkK0SyvpxVGq7nigQv70bCJUWsm+YlHuQ/PIDJhsiaWezcLoIGbXZUDirqkO2HJ3e3n
g+MvqB9DL6x9Dkc5HzoKJBbOnqbWax3kDSmIa+U48BM8gJcmtyQp/g6QG1pA98QdkjmGLafasprJ
LwyuLcy5NxS1/uaUIN3VpUFD9suw8609epkfQFcHBRXfeXBA1hFq4ZySYeuAU4l+4Gssp0If+wQz
v7umrDU1rpApd3dsx9XnRH+5j4YYOB42mBm1Hh1Ui+ayikV/FsVNnLRvtHbygW/vulOayDCImdrj
ck/5iSW78KDhtTtQlBtKbF0hkaxJsqSYC0rs0kXCiHjB88UOreTZZ+7umy9h9k38SJCewbVREBYn
1i2Gd7afoBhHW8n7a2Kw14b42jqvoQyqtFdVEg03D9P93D5mWQuxklKnyrRcKskM9f0J7IJfVHUb
Bz4II3wnvPFcWh/hSn7rJmZDk3caBAa0YQ7al0FE23OgOp32CLw52ATMdzRkJFsbF+sZ00BOVMZj
8rjcsRQexk1DQYiwkI0ZwIBEFEAj1WEfNhWobQVuLzUFhNkS+tbqpdDZeeI5criBPssHyeneOtME
TBBj3k8iIHtOViH5vqtr3nWa/NOn+zCcJXqe9hKKmJEU7B5/bsgaTVfK8l2QbJmWD6yUelSxHMcJ
TErd5/xMUGFsaitbsAQkZCbvuChvHm+Pxaf1OWAJcRNyZeb3iSnvjogoGZuUlEfRKkjePu8pcx+i
69nGYXQgQ8V72CnYu+RtsPggnJo2p6US/5INT6Do+r5BN8QZsZXEmf51z6cnzfj4hyc4ifpuLXmp
v49c+DezR6H11aWTEN5bEvMYFAmMi5RRFFTB5jOUz8Xt6rFtkv8simOHVVyhe/CplfkeSsKtn8rJ
+hQjIm7XYvC44hklVe3yG5uVEX5CvQAdZWd13tKwb2pcWwivYahLohk49+AEIH1hA2ToKtwFAswH
gbz1V7aDE5rSXf03608NJxoy+LRn0/uZHqPywVwiUdTF7tcSukLyO2WF2AfeZ7hscf2HnZLQ5oY7
YBzAzN2GZ5Y0p9uzyOP5pRbymalbug9Tg8rjDf15eXJQl1Yj2SI0b5zCJyu9cxDyjaNYr1x9He8a
BNp0RI9V7rPOZNhqCZNnVTy43tUNgLjoa5RLRBcpcTKPutD/2sEH9D3vrVr7/B/RZ/9VaRL8iZCY
17fsj7iGFflYNrlh9MwvO0qIsE//i50sgcMbBwyLD/aLGRrrBt5My2ztZBiHL7LZW15/+mBxw212
/8LHIm9ZviYpZIBmq334jFjgNvDWy4s07K36ag4mF/meJeAodgcZuv4t5a+yoIVkk03KCSWUOeX3
ZNCZGcE1vPkGeOG3ODyRfIxfArCmEWYyg4RbI1lEjt0n9wta7i16L4ZMl/QQNk8YUyfFi0aDm/1y
y3l7ZA/mWeskxayiFuXjtk6m6Pu2ekch9TCEpIoOVXloNemYuiHFOTjJcy+iCdIJ6RLDKxc3Th0p
kaNFz1hdB6UnZ52qdcxfCyprLh1RbsM/k8txvweNhRxNLAhgo8uSuB4d0W1xbZXqPgbAVnrYqEHx
lroXeQST4WXZw9FrMaiL+uy42elRKbqJw/bRfpFNtRt1HGmF67tzYLNPQJ3zfPLWX50o0FKqcK88
YEujkZnUQ4qmwFP6uUjwt4O+kGU4U5KVhC/XRMDY+b2PREA0NtqJAOjzqj0LnYyvmQlK4p5TTdg7
0KHaLfAo/aDkwyNLxXIL8rTfQjplIt8zwPG1g9mdpFNhROZ/+SZsfGE/GZceBZjbbgeypH+NaTHK
fJd1pIL0v+cbt2KgUZMWImAGAb43xoXCgaPZdZ/f6p4UMLP1B6nS/WYZf8zml08PFxJGfujogtes
k8ukgMIuP3mH2jUNvE7h9EXwmmaMLsqgXABxnWrahHTW3GKUX9iaDI+yAW/MpOYpKNMEZGqiTvcQ
719tfOzKMRXJDqnrW1xcsZvwQuBV4+/kL/dy9+FSC0PC1M1NoWC5sXRh+6geKwRPjHkBMYcb5DhH
t4Ryh7KdOJDk4X986V4WeHR/tDLyvW4aEyloeoI2uFFmUCp+/ZF7h2KJgx3ObQgG+53hZ3LHH8S2
JY+9N4ZomL9itWX5d0xxgBmsW/AXwGmw7GG1BgJRIAas/JQ+774XgZFgPG7e41yzfe9P2VQsoY54
LwHw+6vFIMzx+k5BvjE+peh0LYYa8J5WEVv7SJI6fbQip4FwFeCN7H0PNYnjsoxGQYtp3zW7h83S
PuHn2EQj702/T1fXlXPtn8MnTWGYkE86+BwFfMa2GsW1/f0UpnKyoQMQOZ2B+fY5qGHRp7hEbGmo
sEvU+YiIqfw8v6MHk7hDeW6GyiSbES/ekkPnGoSx2FPtjuOEGgpSbhwrgR1+rV9y5D2OK2U1OLYt
t9PivsfOgFXj+M6v3mYFyI+DH72rxue5NLcuvvkQR8332zGiwjbjHjg9zRldjj7YVUFPb16a8WyJ
e5qJMGI4Ed2me/929KFBap4Pl/VjbgldcQ00XJsBQvubNmkHGOu3LYQfMhpbWsi5ZRd8V+bvDPsG
+dc6PkCZ5njQt0uSjRVrT9sL2JafBE2Wn8vrVsfCr+nDZxi2xwB9FbrsxqOFFtPMblMfm9zohQpi
DU9LL3CSy5eAf8Xst1yOYKy6DfwU4asRVIxwW6hQk3uvix9ebKIMUhr5i7wROtQHsQpu1hHYM3km
NGztmHwVn6DG6wRHWK1SjwG83eDQvpWfYZtnZaXCvKb7WivvQgm9iKGYnELtka91KXG2XTawbkZC
51RcbE44nQyoF0uPgww0Pf87AHfrPUqOYI0l3BbL9WRKLYNXkXYUY22i0cExMvJuYbVc+humjUIA
PxHDNk+Svtj3E0gJmfQtUd56sOgdTHqMCq8eatXPtQwuTaeYyC8RUp/zSsnW5YHAr1r4+O7i/pz8
oe4+sNDppvArHQQdtn0jFvd5iWCCfoago3C5EzXdeQYfm2L0bj5bhiErte8GWlA0wKZYOtNogJ9R
joICQqs9IcbuDz7t8YVaDSDttIojaq0D62fr21T9tYjYZNPxxSPd6LdUL8qfXK28fhLvfVuvB97U
yKdabjY43LfmKR0UDlCqV4QpkJouTmkzSQUDhQyV/IUgTUDHDuFeS+qgnbYwkMdo17mlq4SsH4TB
yBG75aJBhz/G3WInjV/IMZ6rcw8r8YVknZjw0iPBrHBrRPEwz2d4BJz6N/2MKQkVJ0TjrWLgXnct
CXaEonmZmAOVP/FuWg8ma99HQ8lA0/EoHtbXLsfWRTulDzKFd+6hNRcPFitXveOky8opSOxoZ3PG
ADgM/4QDui+YCq93yb8RGBYmEb+K/2TRu+LlrtmWkJkQLv76sUWrCdyysY7720MnXu3oa3cqL14w
RS5ugPX2ZMilT6QIBCE1fbprQQhbRRtiATjz0b11SSf6rg+zFfxt2lH+AZGkJKlW5HZb30f/hdOh
raAz4Xif5g0uWAXuEnbc4jOschohzSMVq0y5VE6E17N3nyYy/fzIERe3u7AsSqIrI7+Fr1SS+WA3
nKIlofGxbW6M2NozbA+DO6HFULslVcyFwBz+H2LYEwkTs2riKvMpVlRlKP3qB60JgOVp4cnIXsH4
IQ90YHPb0i+AlIyqFhxnAR0TL9qEDPXNiucHDK8d8VnCFFtywQnd8hw13eREIUYV0ufogRX1Njgt
xa2UP8JUQdh3AWZtK7I4Ui769oY1NUWwKsE3MfGlK6EEAxghNI//tk1hOFWHfk8Xx9ogEANXjis0
TrR2t5i797Db/W9VmwsLhYKngG/8rH3uYgMF/tFZ/Rr8MtWLi2MUfUNvAR5Bk78WshZPYu4/nmQT
RGcJB5VVqNdFcBDgrnrr0Q783o93fVZkrY7EPFOsVeIRxV2nFRmVyofF/4rZGk8PnysAgStye1jA
Gn0AfrhkcOnKpTf1ZOQe+5Rq0xEr9pZSzuCLM7dI5mtfXAYJAc4j/iV5Wf5gPPcZ9qYg7JCJ8NaH
xGKpDQ93cqoMg6fY8NuLikLlubMh33R3HUl6xz84hCOnMrsdCeDH0e17hi1CRV++yoBaxoJjW4tz
DPeNSVlPbVEfZc6p9mxYoJh/nqXmgDh/TsriPyyrafPEDqQtQG87qeoYhufNs3+THgQDhB/h2JiJ
7uuD1Rw1LrQpZ44i/Q5z+wIppDmVUbgWnUyXKfXTShiAggUv8TMQcu8wJq4LVHKpRL/rDNTx9Ij7
v1juvvcc8J1euehq3wNocT96BrAzzLCG3UdIMmZQhDImUYogwtUCFw1uCdauasWdeavmcLYglLI4
ZguQNAlgTOhm938YIYsveRAf2bBrFiCZPcmMFD128s9vmdZG5f1xn0FcFfn9hMmOoLdZHUTU1KD4
S1qvtDyDun+DiYvhhP0qUWhew9s0BW878fhX0LrVGW+RsngXarZX9Kxq0UcEurcu6JyeE6w+XHX2
nQoCHJGWChhlJSTIDxol1+owEtfJ+iw3AJSrAvXVEpUK+6NnPQ19iJnmRmJ+7pczEJhrrhiTf+Ue
0rys+z9Rb0Hn1jlJAR1pTAJxsMpHs3640f8zaM7n2FQX7FSaZoJnsxJVt+cUErQcW69J40Y/5Krg
2NQX4yQhfFCqlnOJHScARo254+cfy3l/vcYU869s8DxgJdeCDg9sGBicvwm/u1p8+ib/6U6ka5MP
Pqe5W/F69zCBbeKRtJuS9XJI+FjqXtpeEmOdrbK+lrX0h/kIM/WEeoHN+PIdyf/8i6MJWsXUNvoW
S3OEkGpj4GhP6n4y45bd2UFS/KCY3ETsUSzoyyxP1USORu6CEWYdDV4MQuooi3rrqNbbWhID9uRj
S17g+Z0e3mDZAh4EnaKrdKjO7qd67wgkfMTWet25hGd8hjAsLieT1DuIB7HS2gVoIfOHAWWff5g/
nQBF0HXNLLQI4gxQvgNNVn0X0k6/Bz01AduiKjubHHEVui5cqKMmUwkq4Sb960J+CbHvuQaoTWUH
RmN1z+Y19eOnxr9ylKIeoVsO/reYZwF3BSn1l1zR4iGpzlZXtBr161+cSXOJK1x8OpvoObFQsJHZ
cO854JwRuKUjKglIwtP32z0CVF8k6P6wMD7qZ8B2Fx2QEC46KhqtBbaDWe7o697J41vbwqT5ccjj
yhqUZClgxX9cBt0rlkG8mTLdJ3KWcuNkp466z8yU9ZwA6OT2LhUP8+01V8CtH/FU4fgb1q+J7QBx
aAzAdPkczrpZtWHNhSvx4IEV+rHlQ0Af5ZlcK0weJ5uK7+JljMMj5OxuNBkuBdJGPSgKlWTtWZHW
ug79XWJYTsH2DxA7C4ZhJMhsZtefdPsOaAXrDf1k7/o4GSdmNcxHepMS7eSRH94RZT23cQSbMzTA
+VSUqNvIrKClE81+ETtp4IR833c60F5QPeX1aYrNXQAweZY0mqxRMVJbfLda+e4neLdT2kkLEURc
BG5Hus68wdGL7aa0ZFriGXFt9JlZi00ZRlpmi70jDLQs2DA0a9QiFY3s+4ge0pd2AakxexCZBVRN
DEGRk6SWToETq8FO2KeR2SdjtIuf3OsmCttO7BrNru16O7pncH35CagyOm+TbSxE+K4rdqKZScgi
PMDtvmqHA3xEZfKIDz0i3C6V2/qTzFVBJWxEiQ6ACIuniY3xyy4/uReFTfB0Dxge/PCEZfqCNjgz
XHjdVYxVf6gWKyq6w6L0XUOsCtZ94zNwMYKphRSe8kdjQ7rKt1OhogoqYThWdB5+jJUeoxytBoMa
L+cVBQFlo8k4eih0DQT4BlDfPlDw9TV+eyNbNcMCy/xs+cDBVk1+RRA+0FuJPCCV5sOm7lDSYvH3
A1GK9N2tS4Pnq51FH2cggF9PFNNEN+ImEfqubHVHVaxpxyQL1a5VGUUIVA0P8bdGbCi2Rg8l0UBi
KHTexkxZiYMnMOYUwmyJBpsfeCrCMkjL9gAi8jCuGm3rGRRdJ5mESpBYMajayoujsTV/TXL5ioTv
TPmVNlCrhDjSwSU7AS8GyZpXh9J1H6IaoUNkWkknAalY7CkecAZrgGc/i7++q7nQK466zWAW8sil
xBiSzJdnvIgHEaUCIs/DIY9boP/7XmNToxW/9wErp4XDzN6NN7xWjDp4ci3hzTEzOLWX3RWrtT4d
vczGd5CUesKEi8R/euf+srK8naeHWe/LroV/XdzxLb/6Q8eUFzYMgV249lbgjpzQAkT28Xb/4zhB
W6xBtr13/tVLLoW782kuqNrMJxIsZZurj4+8qctFuRKszDRPw/+Yx/N5wkmiJcB3kBelpBbrU2TL
mcvCAtL6BFMiSVG8C12Wkq7oQnq7mv88/fCnU6kKlbyAFCZ3Dg7yDk/YRBnYxDEj5kOycB74OBWp
fT1bZ53GEPoNJe/O0RV5mHbGAsxK8UrlEAXUv70JvEh4J/JquynQar4ARbTtipMpyX0AIx3AZ/Gz
6vAFIsfkyoezuPSqnDYCxi2FZD1vT2EeOfDQy255dUb0ILTYZp+u5mhqIUdlLB8LcWLwrXoNqTbJ
4jJoHbpBZLqf+ggH/cqEp0xMis+ayIhD+H0NzvyNl8NlOs/n+u0mm5gH7E8gIYn6FJzLE+L6E1Ku
9Qu/GvkO5qZoyrEewGKhySK3wolnTaRS+M4Em1FxazFEM9JIFHpgdEAHdfdaF68wSXYOXcTBgDvN
8ZZ20UHjIzSACUbC9ugaUl10zz4fWYjN5O8Xwm33eLWA6Oe/s16Ahu/4ynhIwTvwErJ2N3pZUGE+
S3T97xDKZUvhA6uud1r/bYDjXaO8DkO6Qv6HQIm6YcdBCPXLTrkugLFORT9psEJFSuMOVJXmWKnD
DDsHbWvpY2nk/zwMtin62SkVn4HUNlfXdFSKeuALvACwVv7VP7ZyPpZKom6lbM3xyd5LNLyP8eDD
SvMeENJK84t0Y0+Jyns5n0xgTtgGN+SEosLyR7F5sz9CaZUYBqy3U71/slm86lceZ3cYNGUtPNmB
Qsz1WZTc3Y7I6D8gTVggCukujXgrizorUvinNjbmLKuYw5sDZ+t1vx9uZDy5wIg2dkV3JX+dZiEI
+8AXtUoj+NYMDMiH7Mforg2pk2B5rHbdVwBRHedTHS+VI6UErx0GX6TgmQDqA9PvEJoWNhgtcwgZ
2h8hBfombfC55yeqaXhkfoktCcZAChoRFfxPH98ebDLe/+8yx+PuLWQLBnn9xcsn2N+2NyJZADUr
1hk7k3Zv3NmiUqIE/kpqMa04cEB43OOb9ioYRfDVa58Ti25s7pvG6OhaYBK4cCDqIbAIa77n2JWw
06KEgxGo+FwOPnvOXUH+NKxZKB6FkhMD1Rgl8/U7YGdOu4Z9SBZGX4TwBmkc9pwm5Z4OBVycyFTu
dnTveAGRcYKrBGwRAOtObKCnNQwWS4sVsyGndz9ziLpCqZKXzeT7ZJ9yzt8c4NQYwm9r2cJjW6lC
yFbs67ZgmpqaBp2R5OzOmvyOPuDni0eo0bVDnvh8XduK0AK5ESuR9VOFOXsLQA029W2X8XT7po7k
F7UEsZJKIZNKisy7J2Uq5QJcSRYMpbaZ6ZXA3+dqRAfASagdAqb1Gt1OHd5xOD9VNWDTsROoAUDj
e6MIg0tflCn/2dYYhJqCGE4TNiaZCRcJuQR3LIIV7vcNh4Z2AZf35DBg26ii/hoYdRkuF8eDEbQL
21Tfb+NDBU2JwCRSuU47vI5aMZxB3MAETwtbgLBn8VqDp4CMCnDuFFOB8XIgb0LTKP2Rp3z4/1/q
vXavjIaenv852WUSUTCxRarkX3ipRM9DqEZ9KF0LiAst+dPU6VtjRa9uj65HpE8oZ2QDKFAdltb5
2GO5eq6RQ/bGT12S9qZOrc4Te0HBpRjzHxxlu2+E/Klc9hyLkwCwQXfHQ7JL8tmLR3XV0+8UINwf
hBK+offpaLqqSId07Exdvnu1ywU/KVvAiU7NlRxk6Tg0YRQK9gTPSDfd3CPbWIsrwc88WMMqDznS
ZPCjYctAKP0O8JNg3hthlKegr+eXcYfE3M8Wq119v8bXh6dDECekdMGN+7V3euz/keqQBjny0Dzw
ZlZPO+M6F5mxUIZvvCek1C5cAjRSt2jBW+8D1deZNG0QKAf353+BSelBv07SL33qPY+CGYgY98LQ
dczezIQe2bgQa9jwOR0MP2uy4HXKIC5j/QruGomrMb4NnChNK9Pnus9Hppy0d2KXC2QQmaFEKEb/
Z4qNmshogmJhJSkLJctVnazaGKtV7P92YUAy5rXcIGS4isRFtEczQ4GWViuVqIBb21AFRxYfdgYq
srMcY2YrHJZ6ToDoGpei7UqJsccL0gM6v8vDdAj6k7exVRdr663eVxfNqJNXk3YrrnQbSI3V6PAl
dxVMPkQWbvdEED6EQ0itPes6LzjpvjvoTaUuBQ/JJSMTq2RxvUjiFKdXAr4ouN7eRb784Tk4ME+/
hlrs3h+I1PaHMQA1CT4wKHqdIJpXUmTqdcshsjjCBE9QJlp/kpuwR/U4hlCiM0LLKgW1WgvXyBUs
Q14Qkrn6MINuNQIpTvOW8jfoK9fcnik2nmgWLZ4PlS2zE1WgnCZKE0ORDVETtIkq9hMHMxu9rdla
2DQ3+uytJNnGSG0sljTi9Sx/7hGJ5isWlh+zgDXif/kDQHxbfn24Q3EPodWPKm8NrLF404MWCJQr
Af+UmOuDTMDzEe8D7pVBcftSolGNG6IgHb7oyFOvMwpPrB94XnICbSp56hN9GZ7N7tqVebIORfI2
e1pDMV58et0vdN4ZSuet/2yY7xcxwbU39IJDuAiQfaUKKrG5lWAmW92yAuz27NN+R8Nnbdv/PjQ6
E5toIukKOG9FCyINl67c1ZNXlYhIwndi9NyT9yvt090lPHGhmeke9fOYufcnaUS2r/kR3jI09c9q
QizylLORq7nsgYZL3cfjxKPfsC271cIHUpNsk0SqIbshP0Dwa7CSf5HozhkSTm5K66ev6mxuJaZK
xkL1RXTerfcvDa+b95r18x0PfoEbWU7bj95I8ynRIx3CNEUsJef+j5GEeoA7gMIInDvWvIdthEME
HbMy1G9qSkBm4E3L5j/esiFqFMCcj8ush0DeGB9GGfV5xeraCNbMLlLcXir6+1F9/SjbIyVqi+3Y
YuShkPz5cYCKjtjho8VRa31IKuOlV3R8ByPYBBwv9ja/slPfHRPwjCEMxuQkOmQoIAUQMLPl9vqG
/O81xSsg7haD7LFJXcWhRI2PnGJFHc93sNAOQ5sgakFJ4Cq1SYzaETap1slLkO1JgOLY7olAtsxA
QR042ElJVxEjN6HEtMvEz0loA0OtDXs8IPpUgr8rMuJxVXlI8BYmk4QgPFWmimQZtsKBsqnJzLLR
tzxGbK0v0pxsVDvpRttaWTNRUdMS/hywiN9N/OL6P/Os9PUPLzFfaeZEsAyDuh0G0ANw84+CNqlE
tTkkUW6ybMfeCnbJPXRKbPvI1cuZn5zNWXMnawAMCdqumHs8oJQ90hyC/l+gbashcFZyA3elyh7g
7SbQHGX1ULLMCMXH5Pu+MNvJb8tstauOcVvsv+rG2QdHCr46AYiFzvZPpijfH/pxasArjxhlkmoE
QQZKAnTic+PhJC3F5egoivjPc2tilMkfLJtJUqbxxvAR3q70TBHDyZ9TvUqmBdkfZ8FPLeUwwqQh
FoG06t3pPABOMNYJvpAi7aY1bBBkqD/glr5hLQ59wBHXFXyaa5l4B5x/KCKLOVI7wVds6MjEosx0
LKwe6blO0J0Kn4DbFLRvv/7CK9PE5BsKDVX8EcvE1aoDxf+hO/mQfIq2B5PjqWiJbfLR5sm10/pW
bLyiQjKs7A2JBmsp6SQoc+qtjtzpmFL4Qer2aWlBsAAcxs4HLM2JgQAM6Hwt4ut9qLMMP11FB7oh
jx7hI3Re0+ltidiTUZimQU35bN/Lb1s0W8NRR06AdV3bwNKOT6rz4pY2ewJzNBidEOx9vtcdHHS9
5brYyqnwJPHRYRDiMin2ecdObOaqYtBPCiyG0v+DIU6tMG/IVk68iFCUMWj6angcvKvznmF/0X7u
bH3jMxyLCUxBQvzRR98hwqluMr16FYQTeRb3WZH8Ai0BWPeTcRCimws1x2EQLsyaARnZr053M8Bw
FbWWAMjZi8WEr/zY8lolZyyLPxFZyUfTd/kcnctxvUvo6IXR2lz7XWUilPduYOoti/xZQQCbnbLe
uguorVEilMwqyAz5ivtTiAdjHfkIEDFKTJnGsVVolfcqRKZV7J6cmZ3dcmw+9+hHuCE5y7eKx3Zm
DdtBlChzfwG/5cEybrEvt2oAKdCzEzJtWoQfd/lNXYweQwMmbLtAwI9FKNToKJb9fRvTdZteVf+c
a0Ypw9IDdnBfEo0v1UnhNNZcSeLv9XrTzb8TTYjg3wMb7f2Gmj1cJOel/b7pdTdhZAFJZPmW5Dg4
D49lirMThGuj9ME3MzmQk/4xz0QMjT7cVPvD7KYrzCzGDfi0TkQaV2VrHrAtvlr1xoyqbXkgBjFQ
I1Fd0Hkc0Lq3+reSAgM8UZBTU/Io6ouCVLczE25gqUSJNwMHespX4+w6RoZyrcNu6M7jRBRv+72k
k+0wzPzHhkjzPQ/W2UioApMEqsp6NqR+0e6MwbJzbGX+Wl4K6Idca7n3uSebH/tTkB5IWLtUnL9k
OE1ThV046Bvg37Ksem13LRnmZln901dbiWL5MmFFQPvB81+mBnsAThpATwSvdwKgTbrrABkC0veY
UHetciyhdB+7Ctupg6ByKbbjXGD7bmgByrQUJ11Ft27Il4bMHf4TirmwYqXgXL1xEakxkpkqFcmP
K54zC07BsmQq+zdW9+azTAAWgV7PxdbmJwxkH0n8nXCu4zkAC27PI1n7UeGVcIGjR0ZtGati/0bV
orWsjB4PG+LYBVYhcmN2OB4u0+AFtLo6Qpz4y3R+ZjR+EIUlqElKojs5rT9YFSdNqkmAStoYTYpp
5KWQjWLPsL2GHboiECbib+2+bqCed9QC9QT4AOIEUzHb0odwb1/Lh7El8bs9+OF9usNrv1sTQ70b
Uc4UWuPWc/Iqg7P/RuMBaQVIc07MNLHPi42NyPkWswWpyy1QCagWa5qaVwxTN3lYarb8fD9cdwI1
gc/b358BvfQXiCHcM6A3pTDFSmbukIzhqVpgjy+ljjcL8BRg6xvFTIzrdOGMrRy6VOPapJomCz5c
NtfjqzF9rbc3YWfbgKYvwmMx24S8e4Vq7v/IXMMEjrulseT/Usy7X+L2OPhQAkKQZQZ/7qCWV2un
hoPNb0b789GR8XXOyiLXu5tA66PZSXEU5ojXJ0XpP5yvmtqGTRHNfjrR8wUgtzN0RI8UqE2QyUpw
rnJ75a8bNKLiGFcG8M5ZBWvq9G2up56RWTRudxEjxvW+shO5sy/3d5jYgk6xujReQIushkuaM0kH
X8MhoOCzWLBOumCfGS9WPSqNonnGFYK3lad5OM5V/i/0IKDoPITT3KstVK4TLOdBS3Eo6ikJPdJw
/qmnExaQ+u3X1KmyV5KBa4wD0UvS1Xpwb33Jr6i94zB3EMLHxrWqV6JWusyC9FiSYH/ifa8Se/Uq
xevxABbaIYuhnlYsEXGmGOFvbbHGGiJxeD8vXW7knglenqTCPHfobrj807LMvVHtvjfbvibZ+/Zu
Dv0N9xkkDdObheua9ZXZXGmVZon+Iie92ryc1TDiAbl0KSC7nj7z8wBLTJwAwr6yQBhlP6pdSZnK
rUef3GxA8HJETWjAivAzSAwLGuNekv7gsuxvMOgomjlTh98TfliM54jrvVVVaaqJckAawQ/wTFFs
9Eh/u0KL34mRpfzF4TCmram1WcoZtKRzNoe2SdJsG3OETZVPDC2x0wi1UulJnUgeUaMO6QwwCbZt
Y0e0Z9884bAair4568Exm5Ir4jTudZ4WRCHG0KRImSDJh7L7srcVyP/kH3U7gAiJKG441tzpRTnH
oLaxSnKr1guXcEI/55311CwqfNif/wqUIwXNlp8J/5WVBijEqp5vzu224he/Ob9Akt+jTBgEsrEr
2LLAqOOHPuF1Umq0BIKfUqB+AcITTMvJpSJ5+6jbiihPZQ0nQhlglMUL7bwALTJrXjGalRGs84n7
wvrTBcfkhkeiDYZId92mK5iAzvHjAlBePKBG6UL7uSvce+e7c9ydW/1e5pW+TfmzlUpl6xB9Qvwb
KFm/+t0mXC1Idm5T2STjzjtlG2BjE1GWdoGYVXiAduJjZCJLlMG/09Z3UbE0yY72LGUITN0TRun7
tblQVV6Z+WjdshS4RnbK13PW47VHOJkg3yIEDMHczXEMQnCyd4YC747mVDwnZAR30pd14BIR/xKX
zHyhKC79e+AMX66dUpYcQ/LzerGsGc2o51ffzRsNhkNv6JmuJBCD1AIvr45T3t6mpoN5VP/JDN5Z
gflAXBo6bUSVOUL7Fc8qsQWNpU9XR5OJPfZeSPFX3kUGZmySDRKVq4Ym5/1oB79D/hqs4gk5Iiib
ZVWeg/SL+rzPr5PdvM4JQBwHesPSNDi6WriIXh15PYJAbqWOZZL8BZihmoE2sS/+vouic7UomXPR
QPh+VI+kIM1QJ3swDUSrT3jtgZggwaoM7Er5icvNxIwwogiB6xS/jIkw5mhP7gO6RuTqdDIozGog
nWVETEYSuvOGNlDQzypdY38hrYq4dWqt0PVTMdzFsjpjKfmu8lsZU+TsyVQcFygwiZY0JllqCKTJ
Ad2owdleyTg2ja/L/70zKJtXop3ChI4HCzDcn1Mt961y9V+M8JxdyVjRfxc/UClAG4X3eOa+Outd
+dvmOBrNuzZknHdFiOO1JHMYdrvI5jO4c+5VCfaqwz+AxD+S0eKim8yDjzfQTaULsLMVx3q25/TR
F1sMIiyRPlfjNmAbq0Bzky8ODz28FUaIhLE3iuAMyAhAFDk63y26kIJD9RRtApkmxaD+IovgLf4r
rQsrDq/Dq9Qqw5XthT+LXp62rpE9KtmCLnNg+euNcS0nGfHLFpT6HpV9YVV1nd5MfSwLYORUENOm
XZXfhDaNppiKVCzaJjR1nZrF8ZPVFAo67iqSQcnk1uApMI3LP+cLsiPo7PAwbiIqyS8SDspWNBTr
CPpMryf6XGZWzz+MvKA0VNNlWrH5BCfhbf+eARwztDMyuFMHkmtDppzVT7gt2pxp1LHVKaJB7WKv
SVWaZqeSHOH0yFdn5WbHiijTudQ3yaaYtK1Ojr7VH9J5AXmCKfZwvY5lT0ao/HfSHtz9XdZRawWv
83CqxFMZR42N6ZwDlHmjFyk3Nbe22dxA601IllcnbhF70SMGGZJWg1Rsu4cJhu6lez743MHPyC+d
GqZ5UCoD7yxUka38yEVhLdY7PddK5WYiIBdLrXtOamouzJw8QeSEHIpAhtSKdcsqkkqw64EotwEU
wcNASKS3XXhn7rVFKWUe+axbBHmRrAxSR9eflxCjoW4K4cCI2rhygcJxYFQNxOUWvc8G4gMhHiRw
RpSh5shJPU+Ri6ahYGsYVEPgTLHbZ3NvnFRf0B4UWBfHL6ZHn5YvDDjU2food7czBd0EW8ANmr/F
alsBn35XQ49vF8MR0E1o/JFbQi7RTdhZNUDBskX7eCagWKb60Plo2sXzxd4ew01w8yri36ivRIIg
YeLCFtXSmwkFHPK2TUJj+4xFnG8KGNchezr/1Vm751KKY+NS8cG3wUfZWoWIYbgZqavqmUwPsUcc
x2g3LZD6GQeiKovQHsZTnMliB+K73T1n6trUCR4mz7t0cr1cXZ1+OR67lP1jD595J22NFID229B3
TwWOcf0c4q2dwvaMaYHHEjUV2WXwAUAvVOIXaWZH3FxRkh4uwl7hYiEacRltxeNbl6KlYIjelo6p
dw4XRKQCbvKCir2BVQ4fr6uaBDA4SMHkoNOJKAiJSQweyCAxCl4EpPEPtpe14BbuFbwIXXa3W5fA
S5yXTwZDNMFSljfuHEYUzBiUTfF7nuS+mudxXHxBZ/azOWKtECZiY/rSIc1fQcz6r36sL0SSAU4T
Fu2WptVap5hx5ovN6yk/mt37918mbHzA86UDX405UcVAsTfChubCyFL7EVZs/1ecXlexfkaRKGQK
vi4P4lnVNlsKCPtDhwlVVVAxUEPasqMLbRfcQU75I6QsM/fsi74x7386kNVIdaPaOY8e9KTm1VmX
KGnAi6ZjzCeTPTvsyJTjN7Go4jmMThl5Li7N79rynW3YkT6+AHoVesxaiLHp/ugMtlBm2dgqSf3K
F4sn7ptLpdZZACcjrd5tOlC7xzmajWgRr5OTtEx50vKx+6UjUbHJILLrjA6sL+NVMtwGLYOrGZ+S
FxXaVFQ4Akwt0HvDvmfXz/M3jQAmTETLk2+zSTL9hSB+NNs3nqHIpoYqYhq/0R330NLZCeNSGjXo
xlsTSqJ+BInGxqJvTdmNyo6sKflmkb79dqSJOMPhB6xbZnqNCM/pBDlEgZAwxt/2cXawuIoJ1nK/
ShroF6GJpdWTPOVJhyFa5chx0uGciNgk1o9Mfn5O00dO/+d7sVcgr6MQt9CEprftcEOJ4Q4jcR11
uKRytYYbvebzDzsQOHSzXTjnJWqSqKw0cmmDWhCsZIzKYVjlsPU7WilLfDGpQapnZgEUf4Qnv4/k
iAPagsRjOt7pL5dE4k0BAB1Mf8uQhY21/dNYHkl4Tj9+M4H03iL4g7Z30ORFSx3BSjQAKU91wIzL
0y+5+cEfiJs2ssUgQy/ik+TME92lKAXUotfnxUBsoe8NUHuK+mLEGN1zUn/gup5RxysXaiponqw0
bwYzK1+ee2kwaFEld7gRYMb79koZA66VImd5f7NKBAavVYfxmvf4Cj8b9lXXXjT5fYcEw/xkFDI/
IjuLx12dTZl78V1PcYzQSn7QDmMlUoiZrBgOJQzr8VxWASdKwQ8W/sQTK04aO/4sTgNhHZZvG1nQ
m+VVMxeuPAVrBxjiEQsmXVzTNZK01kr4SCB7QC3MhL5KvhwjkM3phSO5QIIS1kVKs1rUx2NeP8pO
Png5gm8wwkPEM5oIgUf3iEtMWdUd/kaysfGSsF7a4HSddxqLeMWjNWhx8/uwG9ETyb7Z9kvRS0R6
82PLuHp6ri3RWquQZoBoH0quaD6dtn0vKamggzG3WatmXUnZdMwUP6Vyeel6QvuX5BmAkMks1HGM
fQB1BrYd7Taw7Z96R710IqzKwO4/baOhKWLZLDfIFsVts/EYYa3GXTz68T1i7ORZqmBdIzJcM7UB
E6SZBLwFkvJ1A+7RjZlcBDXWdDpwUPmFU6axVClqOH0gWsdU82cbOl5j7t0sOSQMWML2bs+1Cuai
GHK1porqLOJMV4ruUXPKdF3m26jaBQksO1QP9LaHJFRud5kqM2MM6hUq6b3RuDHjGTl2BB3+kYGM
4jmSXA0irsFZiH17AjsqrV6F305L+ZuoYJ6RRLFaVm312DsRnStjs1dGav3epGRCXOw1CMxjp1ui
ykqNAo9vNWvny4NXBf6Nen2ptnWO6AUKoDIoikfEr1g2kOPi1oF+aKdz6rpRczY6INBM56aknan0
DsEK3BgUTZd8rf6pJrwBE27aboy2H/B0nsJkMRIseIMQNJpkhseUGevDpGWkXJx9y9kNtodofP4q
3PgwkulsR+j9g1ZkjL8b6vHuG63YDiEpaJBrWEkbK+5kT0N+IgmlVhliLdfISLH6xYS5dS9D40Xe
oVFDm3nrQOt2giKE8LIqvsqM4MSAXx5KPc56k6nYe41uVPN3OxfYdo+HvpacO/a2JtY9/+kQIz18
pmk2tUzSgq7vGozmqSX1HOn7Mjja6nk4PMgMPc+cdx2nahvfXA74cbtOO/Jb+/oM9JieIfedbcXd
0OcWVSsXlhHRKTIzUmkq5DYn7XxXXmvoQvFCTkr0+ERZSXXbhfqA1rDz2pvvcBH3jcrjkNkBfuTY
npKp/M2UCF6gNmDZ6Rpr5yWMNrbKKbTPYZDkb+6ZMXH+tmDixmxR5Hia6cccXe4M2O2Ph5TAdkvc
s7qoSGEezMaRBovEXf+/GMG8iabcL8BffERH/cckif2RuQLdESydWb2nR6CYTGv80Tclz5+r3aC3
66mcbyKfJkWnRgA6fKwTi1uWkTmd957gua89nHxkvOcp8BB1LgO/77w9hpeQmvIt6XnRefXUcAwu
lBmzLszXHxZQURTlnbgX8W/wIJ9/XemcVYYOoxMOmHT6SZVPUe7lcc59TJnWMkqR9t/mcs9C0puF
g6jANFBpmlKCDbY7w2kLF7uQTYtoRXWtY4VvwIXbtkd6zoDcgPh+sb1JNrx5sLGNfh+CTUbWWgvG
RVAZLWM6DHP9a+bi8/GzW55jjxXi+rtDNT386OuF27BA+QTCYEbkrWAjiQpUh+q6An5MPfel1CCT
YmIwtSq1JiHpEN0feDQYKx3wjFfpWJuewV5w0Ly5eQ4FIzu4sSCfIb/997aeXMotIOXJgZzm+vgL
2tWNFPBQX4htC8jAYw+DlYIp9FdQ0j1oV6U5wMpMK7YR2GGhqpovYQYnN76vhdkihTmXUVCLDFyH
m/ku2NwF2yyD0SsID6okh2nO1B2M3RNFOEdZKMfEY8HqvostZ80s055ENFFRmTlZohhLjyuCwfRT
M6zpF9KWdp8K5F8Ev/gXIhDiaOn3PdZvK1WOrOgLTlnM9rlds4yhG4PuqEvcPXyu7hlvUxgMU7+D
TVS/GVUw11FE1/IiP/gx5FOG3qzaQyy/9Clpug/bQyU57cnFVlRbGApx3e4Z3n08rRFALr6B7qtW
xfrlEhr6iYKgtoWi0gFNM+3wTxYAwaU9xTgoPNIV+i5AjpmdGYqLXuCyTemEsgi8z8OrasR4vo3J
1kkMkodOnALpEot0DSLNr85DsEFcXnXiceWsGXohxs88HdN1BqnK58KCyEBrac+wfe73+SaNYaFN
TwVPLQiBwFpgD0x0yjauglfrjAuNxHkiVFZvNCtWfFXTyP7Bvpnfubwc0fcqeDMy4skBWHlr5Cw5
LM1/QEXmgVJMv/e77gca+Z+TvAwJxnPJ4IHZH9Oa+iZtRrUwvfk9aAG0qjqrWIcCLz+PTE3OR8Bv
WhTMwbs9Jfl1WRGMcN9vTmcKFtQhQZ8I35D7ozeHIOAC1UsOxfJccKDY5k+cyMWNkYW3l1i8pYHM
jjb2hhPhSC3Xv1hh/R969Fzji++yGQEHFAZfPUft5r195MxX47664H1NxjJ8yQKk6il6PyQKW55j
aHnM8wYOHZdkFpfCz25YDHkkBzPpJNfEWolnwa2vWVtG7D5ZffJtrqznBsnK45QYCd42eoVxAFv7
kCjWrSlf/oooA5bZBzwS1iFVba1hXkdoxdFoSGIot1Y7QuV7PAnHGu5iQcfe3nDJCc/NqhpYGsNY
rqK72trSRSkrU0HSAWZzFc4AsiLRhsXKvRW2U69dI4G0I0hDC6vxlm/zcjz8xYQ40MCA/SOb1zp1
qDw8kjq4SLjZ0vZG9WpTHYweBQdUeOneTcGYTSGGsCK9IOT1wdPfNj6Vsg6UJH8bO4VNhvnxQiYa
Rb5Pwa6AeFC+SyS5EHh2oYIyw5+yuGYQq5igfLhQ+6Tv5S/QoH5btyoPedcak8y2G/8l5NOnmaDi
wL95OX5SFBYb06EQPOCqiVJ6mXfUct9DTCEtWe5FQ4HUuGQ1bakMRoVcQpPSie/stT7b0QU1Chqq
8Deq3h5/Jp7ZGVvEtfp6p2bwBoGcW7BWvQISyNh6m0KpqRf0Ksgp2VLyn+XCRT7RSIt0nGDurmNQ
qPe+mg2yEIQr2HfZ9+Z98WB52kJGk7NjwxhOpy446ad5DcWyIC3V2F/zHxJLdoc21UxVI6WI18OV
ZNfrV8R27jxu7ksSN1x8IXTIC0DYFwKDGsQ+D2JIHF69ej249nnCxfcAqW1/uNZSFXyZimLYbKiR
DIMRbe1ye5Q0o+p1tCQiy18ew97MrEkbz0SYigPqa6q2sNFfdfwflxxQoRim2wiiSYAssdXhTIOG
IC4Ozjnc4hPcQmMugJ8qrOFMX2hIkFCogRqfzjZM8bWHhms66E5sBtNVvyL479b8p5EzMCB+T0eW
HWZwo6mHjLJ4pHT1wtNi7iS0HOI/lGzt0q8LssxrUfnVITxNoaPSwNwezU4sDONU7KpSwYNT8iCr
WNNvPVNbTm0lfYK2xHcuSF0d1gvGBsc11wx9y0LyWtEt1V6OeZluElR8SSLe9dUGOXbA7znULJy4
P+4djmmri8PbYq8ouJVE9Gu9KF+4o0Y5sI1taK10PFuWTF7vl+RvgMr3O5L8PgCYgJ0YUVXuz7rk
EutsGI+tSMliX5qHhkfe+ItO1ChPuzTXscftTs4n8PB3XrFsyvH3pO5KJSCS+CfIrFDqMiQ0JmvH
YvagKpjMclzRkCIQNKg10VmBfidF74ugtmDqWXWzEMvgH/yVZvUGtoAyKIfgQGMMcSNzcGdwYTGp
ukLVfsRjzDGAYnYHeBrmTfFQ4thqW911Rmt7ckv+epcvjwNy299nSLKZzJHjPX19RCuLiNP1tvDK
QNchf7HxjYPqfFp0JOok+MEKukzmikz5405dnbdCot7QJt7PG/qN8qajIh3Y4Ie2D/EdSMnVg8pD
HfJSx5Qya9iwBvmqmBov64DTDFU5+E8Op8mX7Qm7oDRotKYAAUUw7SNBe2S3d1gtpZaYxNSw+/sx
Tc4kFzW7WNkIuf/wK/a34YCOQDP5hICf06IUKe+z1pN85AqeLcMazUBGzjPDOFgp0n+dM/tLZS5F
pAVMSy+Roj9fkDQMi3dvlWhBTolsm4XR5rCYr50rlXdoCec2Mod00GGP8Zz+FchEuFa3Yttfkf5w
USIBXuAszF0vUjArOPjKbPPxLvM6aCIem06MKqES+7E+O4uJrv/TlX6BDGuSk4iNtqVJvFnDNK77
RfJSQwSfO6+Tb2eQugTMS1yw0qDPucUjZslVwE/XBxoh/fPBTpLjbWmOSOzzQ98WChXIH+IttaTC
W+ra7J08J8IE8Hu+KzlQzbqQUdXhC6Cn+59pa7YHz9SGCvKpZ/eqWsqaKBzE3mxgI488pQEFiHQk
iCU7j1opV5Z5Bev3aI6Q68Zo58+dXlNMBAjWY83/kYqyUjj0/jn3uv8Ky8mw2Mdrv4NhYz2TINNh
QA0nZK0hqam5wDZeqEiKzzKc4tQ8BigGNNVogDvpVxeXn7mjqg3wZVO4zZ6eEdp72JeYExfWGEg4
CR2Fvz0heTgb7PpqpqZ685rUQqrZBNYVbnWsQneXw1j7SJlFumN0Ra0iqp8S1y+yxkoJwGubppJu
ke35QbFKBzqo2SfmGUWonrAcXs/lIqGPCLXjjQayZ8wHE1dWmgvvtMYGXkvhOnwFku4mrGpGB89d
Ejy719KCBhI/zDR+dl7csLElSkEqU44RXobQb+ShKJigSewqXRCEJXzIEeyyw7KWpObcr12hFWx8
dJ0TVOGbOuKLDDJIbxmkYWlfdwxubmTgGA19BNtN+enGeoiJFTgBf57o2DndjF7eSTyXjy982E8q
IuKzJgkvSizl/6GIxAuAgrtjyb6a8YCae0MSVaH/2/1X43MhXSJt9K4wDMcOOWqIsUEBcMJMv+fa
8o/i+nhMYP2Pl3wloqj/79OgaqDmPLIAJyBsAhQ9NBH3LJN+Vuzuq4qw/VHxsGkS0X2H9ZAkyH44
oVvuYFHP8gGAgc2ZzaVJEuyXEdMiAm/M8fpGNkYqyrZLQk0MciyF+LLHEKVcuj9Ozflb1r17Ts+s
874vuWt8jvjWYA+mnJaSMqvRhAItTISEZlmHuGa3WXy2AxvzkYTYTpFhuD1GND6Yq/fAnWw8b31B
7nkfAQpJWktJLB6Y1p4mtsDmIfvTU0wO73a+eLH6Qnr5byykdOk04vwz1AnveshOjvmx+8TB8jhv
vEqdtejf3Cky535UgplCS1vxKurEhjiKqbjm2K+jzb/8v8GFyvJGPfL2bTFjGk8gin1HqHvCoMaP
0mr+4Ynoo34o1PednPENlNTVoshoar/r77JrgGIa+NOgsotPJkeNOZ/8u0m4n5pem+aWMQ+Mif0n
PSapYZ5mnes1PUsSOrW4k90+DWwGxLNZidO0kfPQyHsBEn4g8h8CINR2vi1jUi4qU9Aii8pHjXbf
o8OBomkja3BnB68iuZsMiFH3X9xMtLez8TypOIQwTAPBWJDYTzf8xn9s4sGZqumUiCRVPOPg2rTr
Mkas3y5VMj8ZYrAb86gu+lYt++PvRgA77TvAleOVHNZpmIB8oC6jMlbKcifAc7vYzxwP87iH7bW3
MJgdz+kxkNW/bA1PzMbKuM/fVfj/Vrt2uhhO7QAZylgQjOjFQ3HUOcb/JxWTZvcZuXjFwiKt7Sgh
Hdqiu4B91VfDTvdek6+UwfIXZwR2Xq9b6LK3SiO9G5g33bEwz0JJ3Gu/DujVEnmdh1AJ749yiqet
b3Hg/1rsvTkpqhlIUjIxxOyXdWsptStc/Cj0BC0srkPPAhIM4nTqWu0xtWyHYF+VGuCy/616vB68
wdaW5ByVVXCe+Rj/htiTZmOkl2G/wxhU7K6aC8vsWacWvVOOW4gxZDtA7P0Fr1VbJ1TPNTMwnA3Q
uWBxtcWxwOxp6iaeog7fHqm2VNg9qwZlmBAhQcmJvvsd98LQIi2LgQ+va6/PYELHGPqvCDOR5Odu
xT/egLpfjHSTGDJTnBYgeeZ1Ni03l8eiSIDH+jkmk+I37aJ8ghfRpmmMC8B2DCNiWUGJ4yCexerq
c+JWdbR9VEq4nB5+PIZE3Nbk9x8r2l6kFRekLU75bGVV65faYTBJBRrsr5WQ1axmT9VJmCmTb+gc
ePIaaTkG0v/01rCe9HRZcH1h9DfmBqQZCydmY4iUyY6/60nVfcA7Zeqifk8dJFNgn7m9c1PEs325
3hObG0hSrP9jYtRjm7IyTPXr77MhlBtLCUESdoDb04dc467zdIc7hnJHxaYaYxD8LK7C4DRv1jzL
LUlivgZaAdSg+70UbHjdFZ0HcGKdZHS3xrqO2PeFcIARW+i+JERFhYhDlfgmwWez1Lcv0BBhOqBs
XS+qMuDyMQbe9p0ZPFsFFj/xBcL6VSb1fBp8wURz1MSZdbDGIOBzKEXIzFp2GAFbOnPs++jVSgH1
eoMjsqvIMK1f6opIUO9i6s3V2SS/av0YnI6NA0TZOJS9oopUPCK3W6LiYQJs9ZgINdz6q9O67n2d
DJfw6EHi2YWjtBu5MSNlPch+x7mso5PCq3GIsBSjyt6gluG4m9OLlpimMPAdQFYtU3uNsZizSfme
Aw+rODpovOsHlWhCGQiVItjMrsI1RVyyqM+NhGmfLjNYCkyx8Q5DqwMk+JSU0Cnp65C06yxo5qWR
0G9iWiVIi/rnJRQIGZwPZoBEES9TXHenJGE/h5ivD/0616A9ftqMb1Qk3QRPLGg9WfTOCKMKusnI
eUbc+c8YPLe0nXcgzVpRO0UAeoggS85Oxj2NUQUTQ7Qhd3Qc7+OyptvA879Om8QHj+dcgwQQdQgJ
tw5Q7X3T/dy52lLI4Gw0BAhhS6vU1gKxk9qtTMm5Ccmo369SdX9xNX/Ep8CSxpQHitQ3TGHpzuh1
I879rPL2N5M1nghcz+lKgWbNSi6xyEfCQDC5rHhp8GVt77NxV8/D7Sm1SLnx/X673nBI+NYLqAM+
/2y5vgMQW4xQxRLMAiCiXWqr2ok4IPd0gKG35+PwmZCg9AF/S1Yidj4+5LV0rQHDQ0YQ2kAhXOo+
NehGk022uKqMU5NHdquhI5ElJzCTS645QYzOCdx5AugmbVMISbnqtmXkFlv1KkhZHkfQAx95pmQd
Sy9cyXGOTfpXkGZFxMwC3gnGNeoeQrcMyeESqnJn9MzSJgn7BdV7pCT3Ty3jB45Zc8vF955EvMUB
fu7kg73d/P76M4BLO/YiI9/vwO25/C0m7HpTzJ4zru4rh6cqhYUtpSQFb8BP5ZrcOdRy7WHMzmiA
i2c8vmrR5Of5z26x6rbKp0p6M0T+aYcq9Fi2OSdCLRPijiX97iSJqUiJIK+wK7pd7EQoARHe+ZKx
xUDVnakyOMHtzn6mTjkkSmYGmMwqFmLBxhAwOUIYFXnDuPr3FPwLip7/xeG0BYXfkQqqjbjLs7Ca
dWTfZqZFack5N6wa6AHFcrokxj4xfZ7wZu65KvS0m2zhNxypxUzsQuJ/FscRikPrRjpaNtn6t1Sm
yeor0z2iT/Qp41BAuwnWRdEK1PF8434La70dn4a+4CJ/JheRYL6L4mbzXtAJ3WHNxiYjp0QV4AxM
jMDeu8m2DK3jW/XNs6uHbiz7PQlWYGDNbyygwHHi6zJ2NHL+0Url1XVHxd+fvQ25lyNT0ibZtXL8
JsK05403TtzYjMqdb/AYz8kt5a/z/Xz+u68gdMFvc7sKXxtDWvBH9H8yP8ClLe76RRfbh6mhA5Zv
7/IgTzJqUU2/neL4iZAcBZ1L0kLPQthC9QRxvLRjTE1puNXDuFtTbrQArbnkoqP9rQOhfcAph7aN
YniInjaLnxE1La8AxirwLAqNHZGfPiS2WIbOE20OcwLLlXufiHd7V+tP+8Na5JNwT1HdJW1Cw9V4
kpmrriUIculla2jpeb22qv1nhNt+d6GyrEl/50gDjAO/2YSEa9G2kh8ybjBt/Bp0PC5TLGEYbUPt
DJ1FVskfW1W+EX17/WrrlofC6CKGilvTGULh59kqD8vgIWh/imuBZbTvbZvQEkimWvaiJU4e0xSG
pzFVJApGWS3GNIPp7q/YJ3cRx/L7ODuk9kj6VuW/7yZVJQ22lejUqJBWeAnF7B+lNB+Pk1RlAIpD
IzlKJQwmn6T04p1td5fGsvgx7+iFHKzjlP8yvzhxUrAMFZcaJY4IofobNdagTVeN1klpo81e75P2
hglSMjTjn8dDMZ4CxazGhrqyhXjg4b79p4P1Sm9BHnnO7EX5HFA99wEuvhneZevHDd1vaHHPEPdn
q1th5IRjKPVgOtrtx04Xvkt454wLYu6IJ5s+Y6Jz/Rw6Zcg7JFOgljXXOEQZB3ITU5dhgGotzl9i
IkrcJzXfUk0gCTeczhBKn9mqVgjz5xF5X2fYBWSisk7Zl4KITEvXUErVRcHSd+iAxl1XBWpMfgDJ
UOEqN3cB7sOAe8CuvrHKdElebSfSjjxOxEyar17/biMuDtwJeZ32BK/oqw6pz2hQy/s+j/wMty1w
iEn+q6d9ihGj1QQKo9UyWzoaEz4r+2MFAF0nSr604nqujf8cfLkN69JJGozuimhWlLd6ppXKElVu
j6OvS25afsywcAM7/y46SsdKmvfgDfWF8hho1Ag1QNH4IXm95Vlk82MDD6W1ItsCkFvVOBg1wuf/
V6Tjt716Nt06AS5ENXBe2gsa4CS7CnZCdktrumdIfR4dSopGt2FeL9u1oKZTM0xO+zpH4mAHckA3
fRCWaolZ4gY4ezhpIolBtqMBZxpot0JxSR9MvbBIY4wW3HD403gn1wjG4AUHIIikbM18A00wPPjF
P2pEMYGw34rAne9bQP/Q0cj3V4wi+Agc2lMww3TpcYN+orrYFB0hI9SOm4+vo/t4c2Fg7LyAJ2sK
ENY9wqsy4dvnoAxqTbhjTJ+/KByJjrsP4VQc/iGTnedSm/0sDWXxwUtHmI7PLaHJMhnUxwXMpPCp
sr8GwULMq/lr2WWmRFDAKjMxEEonvlSoO9gq7tPLKo2El1dwLQuFxrDQyECFo8S+EZ9bF70Ek8t4
CPEeoOeiv9iKMhklUSAqRdhPguW5okW6o0ZqC2AVEsYqmd1akAEbxWO7wjIN8RjHI6JOJ6xN+VH8
ZTwUHNB2VjColYE5e4sEXbaM3YQheN8lug9YxypVi3xvEL+qHb8oV+f7Pzz6VtUk1W07vIy7eMXu
JaTr6+Y0lMMhcmAmBoaqTMyx0g1MenF9xl4CBJm7F1LyNaQHZeZrTZnbPMnqD3upeENFxxNnJfnI
zcM+0QYVMwh+nSh5u0EelxG4eG5yhIwA6+GjkjGb/hWtYoHsX9TI98FIUNAaMIVD51giQryEkQUM
ZBHKeVGocOhxDfznYn73/Z5+UdV08PVj5e3pYxB90VA7LdAdnStvUiio8vwM00WON6mxs5grbBMz
akZQFpJhnXhwdt5HW+PKpcamKfVgg0W6PEfUVKvTRjpQNchcf+uuZp4HasSShg44wDI9HLhZyEqW
mZq1jMPlZQH2SL5BBWRPTsIlbxVriseH3ifee36X0ckVEhwpTUiVfjjWx9JMpRcm8cAITvRV+iIn
awGkxrmWgnaBhoI2uE7DSBENHTyR51ycGYdakiS/3PWsABxJg2QliTZ+loADwgEr22mA9KT2I08w
9OjJhjGOMPKrl68QuK6t9dbad42hJUYbhqGBV9+MZke9CH9XdC4pvLjZ1+Rdua5x7ZBsQfx7yO2D
xnBJcS9qtbfq3V+up7DIVX83dsK65xVcHxeVBO2B7D1b3bwo4mrMb03cmlMPQlKeRlm1/YDr+QAK
0iufmT4TSTDj9lLL2/3TIUuZqAFBBZGyAAzcgXyKS9WF/ARzvVlorfMMIirKsTmTggFDNyPMkwtw
BrWlILcFrRHWRO6yejjAlyCz/85SdHDJwqD/xTnpGjebHnxxI71Qg2dw/2bJT+n9NQYCOFSnTJow
jEPOrDGRokEKjFEh1y98cvxvGW7BLemW40SJMqrL8WonMwD4J0TNZFUKg35XO986zvoct2RKvYq9
/jwcdTII2rJO/ScvB10qMGaM/HkFGN1c4FqQ7aQmKpc6Be6rIACiBqeY81HgpZS3szI5eLkfaePv
drmuHC9QH885YU1XVENZ+y5IFpq0w4QH7hh91KEV26HjXaXKF6J4ghM8/Bb1bMJIIoAAGPHN0Rka
m8ItDRPwXnhLkjbO2+q4pHqBJ951jql0d9psNOtnX5sqes96hBxqeKTMoYyMSMswJ75pBaksuKmy
FqzFJEFJoZHkj8ky7yZZXRDrnKp5G4fwQSrJ8fpiRG/LmNrvSyN9B7UJiwtrHlPXxEr1hCpF7wIA
Pjj3IbWDTLDp7biUE81daD4bf0/U6xt65K7i6OW6bK6gmVIEnV+WFfUa0VdMxfqfO/kiDku8TSZ2
edrtLjUl1Sry4Xw/H3Z/n3ZRUkjso4vvIHd4/MYTfJNmHsa4UZMFKa3BwqfxLe2UN76KDp5xXVoK
420euiTR1Gaz2E3RaDu8uKEV5r/IL1iGpb7orRojj5L6PbZE89kP+GYSWgzhvitev0Ug/SdRyuGl
VZ16N/7AzYTh8VVEg/fBU5L5IwQpCzBi7Ccgbslvg1rdMu5xEhsLipjVVJhAGt/05CMTFOdb715u
Ph3KLFvk9kZq9/PE7WB5hz9tIcRA62zfj2FyKhzOvkNNLtoEf2K0deUqZV8e7S0kBiC/hDQDMzLg
pcuxGfC+ebXKKHuCX7lJVSoJJT9uH+9BeflxV58GB4boVEMpc4sCsiQ2SHZk7yqCuqIFTx1rw9h5
J3Q55TVQ4CllN9etsPQX84q7c+1iz46U5N4ol6f594W40DQjQCU0OQyuU7uMW8KgbH2x+Jp2butM
MysCkk6yFGsWj6ehyXgpxB66SKVUia8X7YYVVBVe50t62Bogzt+t5rf2CmoX8Woo99/E2C00OjFt
3PWQQ7K37XUBpyZiapL2LsJ6iSDm/YZhGQhrmW/EDQ+d/2CLshRl+s03UJa8pFBwywA7yYElblrt
KQ9B/zjmhJvnPX5PVDH1TK+bUDpail8SdW7Z0AElc8vgTvfhCoUtOzqaKPUPnHKw54aOAcUS+RFI
+gMIOGv4BCMiGKlrajHLQRl9bRGbif+xSZ0vwZo5dwEO1HEqFKA10SEAGmi9lcPdmMqKRiqUw8PS
PvCqkhNCyEsMhY2hoaSXk2i14O1SKUFqNvuduYV8vyHIPE/jTPtl1/3V9iektyjU+UDGHl2Lz2vy
b/MF6zO7s3+qc4B/LN2OEOel4GikYZXuTqElGEBDsVblTBt8Ot4EKLdmDrzNuNzNA2IDN8f4WMgg
TM38vb8t6C2x/dKM82ADqgu2aWUYUudm30r3n/F7W8WPYm8vZC8YMul0NJc8VPGDoC/fBIEK0vcE
z/+5Pxv6ffP0ZPop/8FJzsVAH9S8Qt4PkTXghti6F8/p/VkXSEV5gwUSIaum2mdtSYSV97flqeeu
ZxyZkO8GYGyzloynnWSZFQaRWJavJswcZf9WxhpWu5fzuqeFNzdHUGlVJ5GDMq9DgeQEuVASPCdh
6J7ueUDnB5t+V2rL47RCD2E1UJYfpN9a5RgQZulYXDf8/Gevm1gwqpvSM5Nl9fQZkFhbFg7jkiPL
VOghqMubzUvjMXubtQhxsPr0yGwzW00+tqdzkoR9D5xy7b7tvNGnBgaeC3GbPyL6FI3voyTI6Z2V
gAWTrJ69dh1SA/2vDxMuPJdDuOJBz+98bFQmhrJkB/lmAENumglUSNTwux7lxKohQGhjqSIJBBUY
hkBOJkTUEPqyovj7gX5JMqQE0pkK0iXcRuC1nG5pVkbcPJuvjWsuA6E8NODQSp/rvfy9A76fKdk2
Dp3Bb/LRX82+ywtyKKueaM36pbOUnu7yypUlO6Zyd2IeQ5OMyGoFr+yAdjzz6N1jkdicaWNIRChn
Q7dX+Ttse3LFEV9JSMdgGdhfu6y1mWEYjZlwD7mNoRRVtylJx8dC2n7gSzstPn7MdaGXoURnSvTF
DeVm45bwIurw8C62adAB5I7M6OxvnJiHm4QsbTcK6xqxgOqXIsf62xnfqdCsw9kpTwqSytraWWKK
3EKe5dvuIsiQC3NznrbjYZzVs/e4nOEC1dV7jPyePWIKigzhHb6S++nPGbVO/oqHPxrh9n1tI28F
wNgQDZIVo8MICyRs/y6jTTnQ2wkVylhGVMH4orpPRLA1ZNh6zv4DgsqM6TzMNnNT7lKSwR4QcM9v
nrvXZoqFj4gvIV7ePBv8EmG2MCRH0f35mceOjgQJQ6w9tM0MgGirMhxhJ1Zfxyd0XHl6wieXPjbw
mUczCiqIGyC0vOiLEOsSJuDFqeDR1iOwedvG1HpMbcST4zOmckeZOjVk7OHumnI1/ffHIRqSCAxe
qJs30fSHzclJuCUDuy2os/LhSM0Nerljt+F42h3H2S4rXJCell5eHBtF+raerf+F8iaTtntFWpD7
XznlFb66Bpwsk9ufC2T/baQ8emI+mVhABpZgdt0wdhkKmGiAsi4GhxiomBzZc+OHQzNotRihjoSw
QTBpgnGICLCsFBi47sPCGBkLxepv9BIXPQcZ0dnwSIZU+5Ji6DrWGTvwwl+InxM5OBI71NFN38Ve
99r6YzxvG1jH4NTQPdxqgWK+wxXEB9NWD52cx8DPa7QTkAS5XoOrwu6P9N/w2p553OMhs/rihcxm
nCvcMwEq+Dj/W1o53M6En2wpQPR7PXQ0n+5Q14vuOGCQqmMR9ceWmpQfc5wvjRk0NoNGXPqmrnP2
FvBn1LVDbUgry4ifewlZRSP4PW54w0Qrg7rGnv0PVW9k5Bkx1++VZ9ICFfCVQIwUTSCnley3/09M
mzcHa8X4cj4FKAJUKGsa8shvX3dyk6KIgB6yORog+O5OUKF8XqH019y/cH23lp2461LCBZMA7rc+
j72PXARxnoQttl/V4HpOxstlg45pO+oCWzLhT7HwmLzqw+rpRvszYxgM86xPsMLhi4RBHeEw8Xu3
Z8h9Oiju1IkRswZziufkvmoCVheJk/oJtu51woaDbKr0wc44Y46elrvBimk4+tPfJtHD2Yz1ChtT
+RxLiX9SUtd20MkFBXlZTxF+bIQTVtkl9WvepGPQyzrOuV20DZU/M8dy2faxDv0YsV9E8A9aN4HU
9fotCNAktjIBD3m0DnsNCXxKiV/JQMxH9X3eDe676nR5355/153FHf73wptSL9trvh6x5HAV+dr3
Ylk5tqvyEwQSu5KxA1LJNQ9Raf1y9gL868tFnDR+6bcH3NtINYdPl/7x5yfPtpUmaqOjdsljct4f
c3gtTkfLtELtUpLfkqj0Qkr2LSpaLT/hUqh+bNqY//FVjssxdJteQQUIEbCA4ygdlnCdKxJUd3HC
+afzYmaTWXqFQMmUKLA6nxj9xT4w7c+gblVPqA54IF4ipVeMiunfMjo3A17P1qcwCnaZFwCjxJ2B
3MdO+t4tM8vIT+BqoFg5YECduIFTxXTvWGRWTV2m8ksPZE4NVd/EYivhRpjkksjdaoA5RCBt9TmT
j9b8bIFWLHziIlUvEDLTyxzS6iSgS7nl4HLEPElsg5zyyDCbI5iT0wa+VBXWGyWcJ5WkcZL9PNok
Ei4mIm4LWyImu2U13pxEgSI94Gq4FIpdFbqZWRmS9/duRSair0KwNiwS7QBRmTSukEha+dKtF6yd
ycKd7I3paSKNxQcDuomGY4ThSdS8TrNz9jAsUbJYqaQMBQRU84XvjENU6LiOiIdloBhM10mzfAKA
4xupAPku41JgXn+vNdRVrZ/EueFWKmskdoSivSxxxmacMRyiIPBQTIRIiNFD4Ri6y/GbgY/eeg6X
xNnOpVOw76JHcKA4XTgDIzr+QItWZqcCY9RwurMngKmaHppNBS0Gv3DTbUCeYAbBg+XaG3zNo4/F
oYtq8XrVO9bg6D6xjx2cKkWdS7FkRIOgjT+NNBGTYJD6lh8nWt7cwWFiE/iCNeBWzxwbHd83W0Bz
t3Uof9TOtDvWoOgLGH9wGO5lZx22xFkJAbT2M0MlzpY3wVXoLXJmn8EB5PP9b+rpB2BIjza5uo0U
Pb3nPXvjmOYfQwjmdrM9OU1cKpGg5Jg52teGAwopxXLGHUAPwZwSOmRRgt7XbqJOhXHXEd8YbM93
GRiimOg2/gjK75rZPSl7ak3q97le+nppKTFEoFFYqQcEKheWr+Gd3IpTmJRa3NeXNhHsHcWBtCFi
fa1O4BHReJz3dtwym8reBebq3k/6MyCGkLycsYEx5g3FKBjWm8dI55zEEh1YTaUZHt2SwM5VViJi
4x3YJL3MpIhhPn6ofGFc4vu5zVKtCNRxGdzq4fEw4J5qRiV+2WjHsNOlPNxr3eqLFLgeADkjcCWo
qBxNlMFpCkNf3b91QDXkqoIwDBePODC3mJCdK0C/u/1QGYs+/fj6AA7JzrLg6NrxyiJvnouz2SnE
XFGVVJH3UhOiA3+6gvGrLCFDsDCG7f6NeYQbLrI/o2/Z5491FVcr8M6GQhyxjRIuzlLfLkvCQ5vd
eYMQB3aUeUjGiy4l0vvRqka5mLudlZcjV7Vijsetkye2ashSvCqXRwayN+VyMpa9bNDX0LweL7Ry
S5imS3IK4+8AiEf2/wpKB6Yoe+K8GGvujA0CS26g9a8NjoOUiS54mPWVfuoGExarkwZXN96vh/14
N42lWT70/DX/v+oAuX11itnXVN5wm6XkSeEIgMQyBP9UYXAu9/z8FSKp6083/UhzGLSjt+53Pzg2
x1b8zWPwoSknHJtZ1TZ4Eg5XRcWzciYpDnEri8NALuOUCC7G8h9iYgGvkeGkOqzVaqluVgOP5cND
76B1bOEQuOu0H7DJp5CFI/gINDdaHqj34NKy5AK9aPwIa5U7tbyUQzKG7eqJfdo+IT5xqBqWlOud
GF8M9tGZ69UG+lQtoiKigZWMOVqWtCXC1ylRXI6UfGsQ1I7WN246iWhX4P5APZyzp2uGeWvCph8k
I42D/vphwQ26n9ooEyDy9T2+kVsXgNXaQePfBmNEB38lGHJmwB8Im/5JNojFEMcb6e/4DPAWdlwq
5SZ6+vlB4SVfYkU6O8o9wX3d/UGjr3txY/8giUs6duYng/nWQCH4TfqYDtJ8TO/DDNfKgjdrXMzE
TMRID0B+lE42rAF7Aw+20aXyfK0qtDbMZF+bg+IzZiS/mbwhBbTkwcxpeyCyrBf7FSTRPE/GAnHU
xIx6Ej2L82PJlHGeLv2Am/RFugZAWl3LBCs6R/srfluBqCIRDa9d5yZsghTr5qBPnRjKonb2uQ/h
4uCL1FZZrR9qXQFC8KwqD2raHbLaz3MS+002OPlWKVDwQZhCrxbM0cs2BKK7WhL3jz/TV7GY3lZe
GLD/xwNckq33ezIVUa6slg56Lpk3qS1dT/Ma5QRclS0OHb9aNkEd9LipHQvLaCUMr6SiWg41O3NN
XGfIVB7nvDta+OjMdXPZi9nc0F45t74zi7MOUc69zSjdTIDtXALujSSX/wHf17ba7hdV3SCIalKc
DyG/mFRjXBOc3GlBWuyr6oL8aV3yf65r06ZMjHZavQqGArOloHJfgVpNbgDQjfc7KC93KZxeDVk/
ES5mn1nxxZa90eHLynBh2f2ieFJkxlHxodn7/0vSr4TRY4xxsLLQtStnC58lUIfYCXlZeqcB1R7N
E9DMggEcZ6TUMgT0FWRb9eqluqzqVmb4nXbvdo6vym7RMmeN5QhRAXe4JcnLyYSyHDUw7EmMCFgc
2OZM8Y7v5yLiGzrIIMrQdwtwyXXd9G9SysbTZ5kaFMSCweBzem9nZ5+ptL86SJwB3HuVk9wVRggU
GQo+mIo4m3QSh28QaYNrxiPtQhDO6SKtwnPgat9USLIaZqoVW2QtPUQDCA8TYqByd3n7z+hPfSeW
mG6c52hKTZIOzX2/Ji0LZp970o2g1CLi7Zcmeaffq6rOgo/1Mg7cMx38bAfwY1i+fTBxx0IkfWi+
5t5YqnDWhKfxgJubDns2Q+nkLxUCH+BTfZhNbBEBeILMj+zKs3f/uRYIX562/iv3IMX2/p9eg9eD
pQ+xOxq6Xp0vV/4WWEDCtI+/keothbtj58pA2dbhIaE3hob2F4lcbUoB57mVNu5qweXu2f17oQ45
vrZlPjrCm1yCYhOzVTuuMOkCn2m43QhLZpV5tBdPkL80iclt1eSHUG5RUgtafeUviE+1LpOx2w74
G+ttHMIOzMzrU0dhtf+qZEs8VRRVzD5TKyku4c4RMwPeIFgA8rVDKI/FssgQw6Of7Zu9qxOfh5Jg
+GzXa2v2GqwMQJCxv/eicWRw9mGL3i9tsKsjwfhzZaTAlU2hPWXlstD8XUekojb9Kprx1l7Us+YA
0f7WVZL6BfGi5Bd4Hds/IuY43r5nhbAB9BRNmoIa58jxjoMloc2lyalW8zRi1aLtZRZHfFlNvrAD
RJBKGnK9Bo+W7cbf1Bj3k3IhhxOcmrBRrXp0aZ7xF89A1vWDsa5kQMREnSawlJL0Jc6zQ9hHp0yQ
5Kr1CCmtv3Cv7tpu+rw0qygKkEMGRASdoiv6WgmVXYhe7rfezfeUFbZYI8FNrRAca3G+fuxJrzQY
I9Mnogn4hF0QMi6B9PQO8NDTRWRIHjlxgwg2twbMCFGzv+yGHG3QO0Nv8e0vUyK9zGDpyXa5GAps
l2E0F5JmhPk/iHdMyc4mkmD/R3t4ma1jq759UyYUJNqhStNGHjd7yFxxy7M1sMb9RVaJEUAMPwhB
cqBVIPUbXDYL/UZNMd+EZSjcptLWr2Q1Yg4u9XMuUQK+51SG9Cg+OLtWDT1v9qr587BuzXONAmNS
oKRRKdwCNGkhbyamxojsqEfFjKqcoTV3xzxgW+cYkJ1oiAQZ9wrzfQ2x5u2xAihGWdGiAD531LcH
O6gEcbGuGqKlnPj38k3JWsMCD2Ueauv560Jzy7UIyzZgygS+zQWac25WRYH3dIB8+A2t3Dm1RyYD
rwgOCvPg+cc45n0IBLcu/m5ym6SuyxerfmM7qch7gemWyxmsQBsXlsSn7DYwP01dZjEFYQfQ92RL
qbIjpzl/MNbi1+jDsl3JWTdGWls6du1uvf/a+59/cyu+SfXRUIRi2rCeXbuz32JmiQtZfxt990Hv
trKWoVNb7zQrwx8InE+14XmyluDTmMskxjqXbgdY2mwaus9VphvTqxSnCdf89iJIxq31kfaxvwP4
KTKDSxkEH2VqxxzCbjChmjCI34HnRk5fSbn+s8pCcV1lBClG4Hy4KMbP5f2NS7IXMewePC3IMNJ8
Al8frc1blyYA1OgDWTwdLB4qjFOxdYHbeEw0BCSDE4ehMYBpKcwbA5+d0AleyHpLX9S/M3me6z69
Wgv6YguRcorwGUyp3Nw4C0Y7PAUEC2aLYqqNmEl7AEAKEMDCuY4sYe4AhjwOTeu3X05uumg30Mvh
gBVjAPGA8vJbLBVoQpGlqJh3K3qUKZLMmnZqgbYVaZhBn4NIJEJ5g7raPaK94kEGhS5X1Kec/RrD
0pxHRyhFB7EgexQPdFZTqH4CjeMfpP97J3LMKaDZJfdr78bJ2hC8wapLfb3qyEx9+oh6ysubC4h5
/YPMkLFGxd1utFIRFs3qICm5kMS+f/3FKZnjWb0iBjxFgjYxIRGxy0dwXdbKSjxxuXITCvzSSvkO
Udx2S1/Z7EGUjC1ZEcoyjEqTnfG8/qkVpHjYLTQ3T3t6Z5rYSmGrazzv5LN4H5pZzk0WvmCYaN5Z
dyQgDjt8VWX0qd9Gqjlzb3V+lnDrN8mjONqX/tzZZIiu0rRv/2BdjNTa9gnAb9ul+7GFhlAIDynD
H5o249ktn0SeQfhWjh21HjduZasQmsB4kVAEyZkfTWB8lyzbRdW/ztiAJpG7LOlNbYoPupmAd7tp
pVCnCXHCVYHRt8cp2iUFziV0d/h/IPTJww+7OXRrsR0gtWL97ZTewsbF9CEmuCgE+MlLoVTorozz
pegJ8AnP0Vlx8QEM/Mj4Ee9SsMt4tikkRZcyyL+7eH+jaBdli0t9YA3Sln6Kq3XaC6hw1Bp10ODB
+5TOAZhMDxLHgNLtPxi6UKSfJI6PqqkTrSWwCuivC90NYINWdWO+MmdGo7TgAYUREa6V4j0yFXtK
iHDwFfKzNhSSFCuOkhVUvgG73MCfZyh7cF4cjpx5gGz14/Wd+X3irxLVduv6OcxKPkwrZMALccUR
M3AN2oW9BeEzDdo2RBmZ3MNt2NEXFIxP6oUjXi1q4XYdy9zZd8BKizAAEPALOked5D5QCYa8t+FI
iOR1R5hwmRaIHFkQo69pGqV8A1ecw61WZr2u49Javt9PdvPvtruTTU2R2v/5SiabWufyQGfx+ysl
64bfx63ZKpaHqk8kmoWSJl89NRMue+uJgx4aKVUhcnTLigi6wYOkLvW5nZNvwywJk2FZI3YRw+Of
WjXJDiceVWjDe1TPfjSgxS4sHxP6LnJbzkHpELBa+HHdDTnxsfROllwuuvRLTpIFj2dd2/YJOoaL
h7KNwqEMIdqmdQ8T57Wq2ARM3QVyIV9LN6DSOWrgfLSEBbEAIUDpaci3TA56QvaRhtxNretGrbdt
IRQk1Rq78ONND+k+lcnKeVg4YUVrdUFrE87l1s1/oANfcIa6DVls9fRvdUZjkcAPU+T/+u20vrLh
yxqGxdkeO0GG0+TYguTIkEY2Wz5G6TKT1oo2rs+UJsHiB/n3EHZpO+bRrfBi5nZVlxDuiNctfK7b
pGd9D0oIGPYwiOuacZltbpdPOIMH/0tzCSA53nDClHD1ED8G69uWIR51RZMSSqAAgzyluOcrJkqp
Lyj7+nHT2ID+E19qVrvVmjvgPxduFoEOizb7J1SHVWW0WfChkJceBVgxiF/v0BeW7Xq1aSwHrVqr
vyJH+XJ1UBCQKxCOVIQzHX9hprz8yClJcXUCdaoj64mQlzfxUhM5rt5eKIJYWU/SPEi9JrS3N9Gk
dZqFDtwxk+Ra1i6I+kK//mazZ6847QekM/dzg8psLAawtu+NcNh+cmR7jmm3ury6tBHeINVv0+aB
/jbheR9KVh9ObX7yO51ULMKBz0GspuDhsr2XGIWQm9XQnxiNZj7zJKvhdt7qmfRBzAjwlRzyHtNb
ZzIIwVxIy/JkCHR0k0/oTjELvIi63oBbwAOeURa4xkRdFTW/jAhRoya5PVr3eVcXEVhuksp2AdDc
+rfq+FXMkfyioZggpYJrexyjHnAx/VLGo1Y319vN5Zs2sm2wD+bljdVhm3xEF8YEto1nA3NuPYxq
6Oc7pnC/WvXwSw+8M10NCqJ65Do8MrDABZVLWZKIbDZkwspweyFaAwdCx+BzvsqbYTNZh9209jPs
tB5zRHUCKnUoepg/MbD7jB0dtzzSoZ65cV53EQRYAwHHQ5TNtup3CAw+EX4E8X6YDLNkNL9ZtIx0
BHsIyQ6q4LCOtdjhqO3inHaLa9ZPrxtfMAaqFGD7CxMpo3zzPBquUmTqH6qIEDKuP07tZrLgb0L2
o/LfMvtO/VUrhTh7z6fS2xkt38Fo3BOB2t+F
`protect end_protected
