`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2020.3"
`protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
ZI4R5vypoUtJbjSqxMcVONT7PWLV5BAxWx9cixOdjGYQW8e75F5HSfR60ZefwzGAhWjULoUZYJfz
DsdWZTLBrg==

`protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
mrptmhCSrUG9kEHdjV5rf93ZXxPKiQAU6Li2tXHwqkWJmdHr8tvAO2KkiLuc0KlAptfFm5HPxRAG
1X49jn620J0PGA7BwW0z9qsWnleQ+M7snUb3ZaRnqdJpnb2vPOUtCF2mFhSrxopGw5xvbdsthOEA
l+I3rGRfB6PP8ul1nPg=

`protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
XhMiUBuEpoKgxhLm9SYEgV53xJxs2k76AMARzBYcGx7rWvZrP4ONJU8r+jILaqA9FRFJGSnYwKGo
YC1fPVgIWKJdhFF6YE6N3KwzBYKFktK6Hx1tFK3z5lwyli4KSVb3mgb+EcRykEAmyHcfmv9mGpi2
J0Yx/s6oNOyREuHBDFjke/QSNT6msc6spygTMKqBNGVkVo9EySAAUMw4Efra4ml2eQuCl3lejgSH
t7lGlycKbO9HrInPas79cIfp/6GkyMR7H+kivZoF2GP0mEptnvmQj7KPQtrKQQXld1lHZkfWw2MI
HREtg69nl06SeiEsD9f9OPoTxZFSjh2rMUrVyQ==

`protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
KXDWcoHD21+RpVtcLpdaAEXu0giRygmxX+V2t60Vk5qDTZdeFjm0qvfu5fdvwy1lemKp63E/YsHl
a5F4SvrN91TlthJ/wz+cKTLz2YLJeE1P9WQKexMBYxpSIUI+c8D+zUUbUgWXd1BjGwzXn02RL/4D
jPhsLLFiqqGXhiYKemIHv6xyntDLINQLaViU2sS0Ul3ueSLmqFqy6qOuOzKym1fcb7bIjk4GZhxy
ojmJQpOS/Kz/7ej79FHhDmHsYI2mvNZC9IMCqJTKqAxH59GE66khpk++DTOzIZtDpPUJLSwtCtDT
BZ6YLZ0Ov1/nb6enDgF0nU6mt5cFDo+mXCDzvA==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VELOCE-RSA", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
Ju5k5PMsCEalrB3X4iBqx1ojyM54i/vmyPnlswL8OMg816CHrwze3Ed7bIqarPBzRXt+vQqJv2aA
Wq3P5oDdE9e5z6303HH4JehrYc8Fd1SQNwER36kwJnGcQfGk434Dg34UyVsVxXOTPTYiP0Z2N5Hf
c5cyOLKplYRWrB4G59Q=

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
nF6RaZkBhBrUn8EhEfwPENHgkqvE51fGWrecla8V9S9MkWkuLmw3B8o73LB1Jt+OKASVn4HTLLpo
5ODgbrS34mfquB6ssQPQ8rTTcg3XEbwZP+2JGi3IWiIK3txVjkmEZv83A9S2IRwwLqnzPHFR7TQ9
qH3f5dq8HEj0nNs/u73S01ekLIGVZfRr4ozbjomA5jVFRv8DGjY/SR8gfu7WmqRkY4s0OtDlOKpK
bRr1Y7jMI00nRJvr0eVL3ada85PVVkx/O0LlLMAoXvt8bm8nGuUX4wueZ8GvXiAG3yXYA+m6Qz2J
58iDhdHx4qOX7ptX3rR8Q2X4cCv4C8ZKtImOwg==

`protect key_keyowner = "Real Intent", key_keyname = "RI-RSA-KEY-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
4aoF6bRKJGX0QsRQF0/K4lV7NGihfHwSDRq52mgBbPf8vTAlT618VSH7OJIAN8J5GUAG+aDTiFjd
EIPOHlP3yw7hPAWlaObj+oiedCkaYAX7J19cCA9xJ9nhGm2Ax0Q3YGG92+7ktqKYf9Sy1otPL5iC
YAJ476bhQAfmIPdqzfSSb8P1MHisXGUzKqPi5dPfYupnirKaw2tJWzTpy6SYqCfpftBFxVORnyfC
7inmd3TPGLvC3UvJZ7p3L19+eulxITiKoazNQVwg+zfjyjivFiDpb2INO3SqTBs9w00ADswdBsN+
l2p8QnEEjE3LK04jfB6OV0BXlmq2qCelxtmR3g==

`protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2020_08", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
g3ml/fTIwWEoJWHqleFKvQ7JAaCkDcvxaSw2N9zNXeB5M7T4tJlOOWAeTM/i4I1nJgucR6052hsl
fCWLThWRsc2i9iHPawU4MJIgjmK+Wfl/CHLocg6YoGnCc+tW1qgHvdDnpd1ngCl1VBoknWfSubIn
cu3I965QGgfXfgSZNYuWe79H/9TsHhigKPrEwLIIFL3RfBueJmZ3UJm0oMKg6OPrrjBhthA8V6Ze
R+siVwEW8quITgeFF0Km6xpRV25r5gmZhjhbUxcFdW6fW33dlB/a2BJK7H03gpx4m5X5uuiTYIkM
6nfhwMXoawapgtg+vLUIXfpiL2x80JyOx3H/6Q==

`protect key_keyowner = "Metrics Technologies Inc.", key_keyname = "DSim", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
nADnYgPUjMeH/6ggHU4H3JBJFAL+hoBt98bGdOwc4BEoTU2UeWsi17W7I0wnyrJooOqnFFDMKMgx
py2IZX2tysK6JuTfBW2lWGfSFNapC8ZdzsR4dqCWfh39MOFNNz4aOYQ8MV+jctIe+D66auVdOaf1
wfTHPyVvRYNZwNlOvKc0B2Wn8Zgts6Te3OzEpP88HmVk9de9kTKouayrDK+C9SNGSlUsc1xn9pxE
HISZmA3Wl7inMKJU2e+VMZEZ6tUzknL5vQF33HK1gAKkPCDMltQNzgNwxgRA/+tRgWpyQePAHJ66
SnvT7yVpLM6ZUVVfLP+sBFkmzy+cgRhmwWo9xQ==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 60576)
`protect data_block
6D9vAsM58h9FEOM7j8uI+AlEyS0pIqSAH2b6HvgybHSYPLm2EWh0JaTKJXgVI6FW1mcSs9SoYitL
4V8c9fjavMfNlKCKDCg0I21gRRalddl7ZVrs3aEQ2BRbC3Wdzvubyiezt8WH8fh9Edh3W3scFN1g
QDe7oqds7OLO2H0nbmKQSJIveoi6h6mNXZiMViZIWcF6oPZNqLtppxnyw/Dd1bhqJ5qHJ0sL51SJ
r0NZzNaGrlwbh9faSMcCkiQFIw20livgF8CnW2+zHWKRFA/lZmVLcD8X2kaDo+6+nDtUtf5u7HfA
wpfppp5TXIFrlqWCxO5pQF8qNHQdSdvTqU6rgphls9zwc7hlSsvxfSJOFdlQXwf/2i5mmDTdb/pu
itG09FtlrGqIiUU8+CbNn4si12zsI9EefxBtk9r3haf2bfuRzgOgJX4+laQ5SQ5ovASavxMWzMaE
5pv5MNI71kpzuzf1PgXhV1B1mVq1f8vId5yQRU1Xg+wdVXWow1618Tf0ErnaXWHO4a/4DQUatfMg
vpqllq+k9aDy1zqKQDd/arQr09HP9R5T+vJehruu8yPSd/Fcpq7pKjspEaEZh6EIZgwy/+F9XaLT
PSGkUxqqokm9djoTjLeLQQrleyhQdrknPY8+iH+40kW0jdAcFh/W/zh8vP4S5ZF9KwyL21Kg3EVZ
kjjverBrdLl1iIMFWAnKewyd6KXwh72z4ZAfMBKpggTZi3ftF+WeyEvGtBm8rCwgthL0Eis4+r2H
HKH0HcoPF3twkgrm/I4r9IIrPx4fArDs0/5lO+TT6A1yM1UnBoYVz/41JdRZN4pz1uPtgoc9gNJA
bHEATZnc/g6SPBb+I0DnN/5QVCO2ayQoCFjUmViPyjLK3zX62ORWAA2qQ6SW3Ee2EbWP37n/SGAP
dhk4JtRpG7lWNg3uZWBP1IuNmkys+nifnnVpG6KCDFVIqqLdf5bvF/ewW2G0qFx4GNjiRtKtA6Ey
BxanrHI+9F5+iWFw87eSECaV9DjlF2dW4zys3zj8lU3evwwScJ9GNYg0gO1P6gKhgkRH1FOGDWE0
vuuPuxfhFivWUayGIK7cQijItleTTMIUP46PkIpqA7vhBrTP81h/j2jbZiKS3+DCqnoZS/mjLpDA
MAbiq8IWvH1xMegc/vPzoBBYowA7z+5nrhfH80bAo3vYVdegHA2LQIK/5rC3bVz1y2pJKOSjVuZW
XXtdrCxrMOuK693moLaDG1che/UGqiQPw2QbCnGxNHAQx82Y6RLUEC3GqDE6pzuBEKCdetChBu5O
/R2YNyrVth5naDAGzcyStWWBMl5O5+JFYsJbA2Wdgi57hA9CgZGNU8oYI8EO85gcjuVgKHmuxFPC
hQE2sx2WVNp6oBgOT7r/O7NduYFCYpNm9jlNAdLBQzqGL5rO2eBRSyV5fgVnE097xOW0wPzLk0/v
kqu3dNoxgM2xqEGy9sxUfXxcm3LqV42WJSdlfsUFNMaaj+Df324O7YgNZwyNvIoiIofeHpFl2Uj7
XPHTxErkzLO/06JiFdVncCa4i3FcwSodXJ0c3xNL9Th6WQNNRR1phY7lvIcE3FPHQyTmzk//c2es
2rvgIPZcrOc3DIyRNmBT6U9ng/e07WGRjVWJqYn7ydssa6bNNI3sdtvnzH5H3asD6seMH7mIRBe2
v7NZS9aoebP7xYYQuzW4eJyuVaZgFUuh4m0b0raG6Snnh1MHAP7Fuui7snY9DLRjSe2k8gDVHgDL
sdMbDAwhiHok1Jo0P2Oim/Rq02WMSolaIcAXN5sAYyRaLKU5SQAsMQUDS1e8C1W2zkHx1aRAHvVw
pjrKZh1ZWhgZpRJV4fP6nIr/7eXnya2zpyuZLIzAnLjeoRCz3mXUpDULa69jJ/vTUhouPLXBvXkM
y/lsj87wN8HfXQ5VgorECJN+2muGYJS1yT/2HXLCUnO+FUFBR3JrhBe3RA9KNoFQCjuX4N6PpD33
ia+f6cvp0tJounPi9w/ZvRnlUPk1/Xo1XFgdVkcyQPcrq9bs0V/duaEU8+VUJ7Qf1lRuaGGwUTK3
6gwLsUFLBGmTVkQEF5bMZyBcn9oVHM6OigWkhyBD0Unx2J/Q9A1KlqDFkLqaeR7w2SWWCqZeuCGW
DnLe3ygeGr6crPFsboPgXB2hceNLhEyXTz79hTSI72fvmUIPcWy385fYdmGa1VNNDjcrdI2r9UQy
MMlgov+Ruzuzjv1HzSwMe7L6FNkauXp0TRAEJpk+Wl9nRj//XfqCMFu+CcCYIuqvV0amLeeQAe6s
Kn//J3XU73ofiwqYKJSjUOHR5FF8U+J/sU7/lead9czKJK+tQdKg8ItcS96lGvXvBxVMKM9Gob0z
xL4mrdACkhEzn608dXsqDF9aXTkCXY8rW1YeRLAZVogt9wfl1YYvqn0kp4q+3xaMm9IsS6H9LjfP
8hMmkpvtueVpYGzDpwGRhwkobGJPP4FCUuIsVGlMRv61JmvvxgeqVNZu449w+Ex/55X+OEsdYvg3
f7mLu/+yqQBNZmGFmBiaYDX6uwF8cgVOjgEiaVvWnc7u/Y+yZOqybSxO4jlHjfxs/DTfCqq0Mjo2
Sc2ylvPNJ1jUvtJcqyL9ycCZbZwJTjdmzqX6D2VnIYyZXIwdVbPGMIkgFBxeRO39t1/86YeIsT/3
m9cQEP/PUuKyyvoyYxGoqgPm/BIQpzRSVQOyNsLptjHfAQqUmYB8hF9Ify7/3i2PfQueKG1+Ckvt
iOjydkXBsI3hmfrG8mdi39jlpIT4mh3BfSY2BV4kuztprRBokEI3ZxaYc0KwPVUWzPF232ATsKnP
+pjaNE1rnvA9BmO5vZwaRmvGY7vU0BBjGjzoydifcOVuXeBhzW3ezvEEFX1UJSkg0jvRL/ApC6EN
ppZEm95ENPp1EGJQi/xz5YS6JvIunzYzMpbo1JsY4hDKMOej7B1PtUEcBVqGIQxZiqjfFQtwHlfd
FrfXT0o07olr1R/NZC4kETLFob4KdQtMlFR7NvHB2uzbcoTST6TkUOqaC+w/HWZa2inu8l9TL7Zh
zzqGj6ONC8eXY2vrC+Tcy7uqoIcAoIQIrJzE4JD0RnKC5/+7E14e0s2tEzUw2xAyk4Cj/AkznIcc
kcpdXH4Ow40WaEpOFbC88NnkiQAomQ+LQl7pD1QpfWA4pRbxhhnVlRAjxHvXwra4klu0uMHyukFl
Bbow/fkMBODx5ulHHPpDmf8/MtNl+O7BFk3hoDOMW6b4mLRB2maETIzcqTzfD1yUCwYcrcGOmU+D
fLE+z6gEkf949TTqQSLORfvZrN4UxAfE6ZE2lnwkr0GmfCGscQkCeZhPPU/75i90dlS7tiLswyjJ
iDqI5zwzjfwKGHVnONJI0asj2nuPaqwgUK//F1Pt73vGCd1esagbguuFUF8479kgYdJthMSkQdUP
P06xH7+kpVeRC7dUxRvbAEdZZSoGFVUby0ArblM942zbrKy4Tc7TytqsmF/lpfbZQ/S60DMrlYmw
Zkw7YNWL8AixTgWL2QtH85vRSmYqYVvxxLZ+EaIZSChsXfGl6KX+I7ib+U4ZJrXojnTITrrCSjm8
peU4gK5IpP9uXafgT6zmFKOHoC1Gp7hZgLjaqnWmzxnS6xzm1CEsWoQETkhaQ8oLSZXgE+nM7WSI
2uMnScR4OYquffY8gaFZccTMxwYOEKrTVcR/WaDdG5z6fwCxie7uP4NLJ/PlyIYMruoB6fCd4tWP
ukDijlrb5QjF8aarVAqD/wXpRR7m2FM6nnSvIQrQ35vibyuzubwBKwkFFtsXjIZ8fPACsq8UM291
bwD+fvVXEFaomR2yZixvf2XpuCCnuqWRQRfsOP1Ui4YUqm0u5tI8+OX+AmQInot0BwKnyRglMcVR
5ooIBfmjl2AS9GvwG91nZbTMRQ/nYoblDyFmD+k/uoySr7r6GS7DiUeJam30lT9L2Ft0mNK51Vqb
6zYOUQNhMIX9K5e+3nbi5bgX8eFCSjigrazO5qUQkEEMqHTzI2ryM8I0PLmv4zF98lF219kkn7j+
AL/ygU8O4PB9amLQKdJ1qD0BzpAe/UIoLNMRUMr+Hrn4tZiep0YhrpjdN3JHdGt9pw+UDYlAdywm
mgEyarnype9KdYlGnCmPjz1/Lfb9ph5AJLxP+SZ+JwIESp5BZrUpUfyhyFF5GLUP4Aho9C3mporC
KxKy6SD4vU6jR/PsjUeqXtaRmmYPO2BOkJJQOkr1sU1unWn+hiQOomh9Q7fjLMvJq9kgy6f9G3vr
wT5hHxNNMfJrrPPI8t7S97iPZnMtsWmOxJVaSAVrhyf6VzrqPeYObHI9Krbjy3lIXOjy37NiSlzJ
5Wcv4r3O/gTEfE/3hjemdZ8Va3PHlARl9vD3YCHB54hWcKRxEE8/c/dWz4gcAQBQJQQ+XZKNTwwO
q1Z9f+qknyLrOHB+GkdxxvixmX5wz8nMGhLZ9k3T6iEUsUSIhXeFUTAETt7Hu/GAExQyQykrxId3
bB4kyF4bfNxt3fzGX5kIXdwfCMomifz/tjSyTZbFzaaegAbHnqWQmNElcZcJA6bgCNdC4y/eClnr
wF+J1swpCqp5GRJOOxt+ESDJGkOZ9+BDkphFVvn5+mB86i5gc5SXxGdPhugxTxQbjq3OnDEd6cIj
jGhAdFRiYoGsv/rNhCThsaEBpZWuL8/c7niJR54eUN2ws1YX39vZ6ftB31mqR3838NR8z4CXHo5V
h8DSolaIngTbxU6JOXnoMVa//0IQJm+v8cX37BkUugo0pEOzectn7kX4KAWg0Mz9z0uFmGW7F1v7
CQHS0Y6MtRAyzf4E2HmBRWnc5zxPXPsJGTdypkKI2uLnvcx8t0gfG5/S3kuCxgSJKXxXJmoz1khN
u8OqQlrkNaoWQ2S6UK/iUcVgd85NCZGZDXaW8gQG63vtEfNXETIMI/jcN6n1d+T2kP7RVaf5eejg
YQW1UkkkO8g2xariPRkhjZjMTAbjKUNfZVV7ppmnXaZBkq2PqarJwNOgsB5OS8TKKeXKtJBR3KR4
DZdp1ANbz0MLH3rQDXcCPtSITSvF0Ucjb7m3Al5g6ZMMT6ngY6QkF833PmXzYqIIUvfoLLpx1DLE
HLRyLz7vhSs4JxpCJhQGM5aG+y7zVghoVMSis6hw8gn9skQq7Y7x/BTkPuyuQyxN4ohpfNzbeEYc
d7HutFdhctPeiayf1knbnOSr0+Mg/MgXzfZc9lRjQqOl6j3IZwWHtfLjI0aXVUKJtFrDE7mOOkQk
IJhIQV0+h9fGK9rO+p6dq+aQyqa8LkymY2mLLGr5p/8izrYcKQHVn8gVuLANfY3NTUtWpY2pLCl1
gcbXPW7KKAJlEFaox6yARrvB0ZWfL+jDUZeimpDiwG3yZWONmM/rhbGDrnFsQxc2bxSgqLBrG/1t
ZiItTbmIDcJsAEg13QofiBk9UdDeKrqiArJX8C+WZutCMvQ+P6Yh4LQ69KyxmIWFgU2zBwEWqr7/
oz3ZbJ09MNd9IEMX8CQgFDRNxMqZE8l65uK75TFA+qTrGP3pZp7S5Lu+IXI3we8rnUKOBBZSTTgy
CvoWDfa0+cTInjDIXmnd64vwqUySScl4/l8/SXSf+1knvXKVHrE3RuTN06KG37n/jracsD8ODFJw
skNABDfQTjapbzZJcgCxWE72f2siP0Tg2O6Xm/nzScPAg6CWRubShSiRhbQ/f+jo3SVEUcWgb4Gt
+XN2pymd8Hg5nOv4vgwGImFzR8VWcQ2hmyZvrjXzUKdROSo1LBlExIlm31yi7A0srZnymZdwzfy4
/fCHbkMEcESZ0T8IqahNoEJNWsJQmm6VQ8+S6te9RRgq0YMd4NCCRs26iU2ecsBH4W0WTfX7+MNe
3GMjEaw+XXsx6r5+FSwCrE8dLDiV5S+yH/xn6uIC376ckO7c1+mgQfeV9CXLApdHDKZf/6AmZEfQ
VLT6tZ3Glcrgzhw9C0gkw/qQqddJxTYIY+2VxkXxRQLrzu9b/Q6ynFSLFznuGHPnONPxEjFuY5s/
GsqyJBR6rW4Je6+11bS5c2+C5fJEpPhym/91f43pfQRFUYZbmfuQzEwvzY+u8IT6+yj/wEbW/qWB
Uqpfm/M4Ln534H0aGKvkgzVdKPnPu4i+lX/M+IC0RJCE9j0JBk2OFsU3Uc9gOFFwl4GVjv4SJYzL
RnYHpVgrceT+GOz2i4Rpg9N+EmywF/2DueZ6pW5btil1qZmzY4Ne1sl/z0spvICoU8ujvgu3jl1v
/R0pC+3s44pJ4uEkAZbhkEAjjbnznu+Y07FyT3MiNzbdntViG5YiuMP2i00UdTCduFBJsKAiBZol
Q5b+stSn7Jlud3XY5MMJdlnVpZV2HLlF2GzDRsjQ8JcoiZkY4iLAT90cPHxXW3SZOJYZGDx1lX34
294AbvMrfqlCkpXqS5K0hPKZjC2c55G4jxqWebg8eoeff7EgYo98Tmu0aX0CaE9Y+ViB0g+NVbu+
WawH5hJ/Q/zda82xIFRfni2+TFdqHixzftEaKkDM8y6Nw545v40+V434bUdHCZPKFiH7mphBwAP9
jMn6X7qWaBwdh0VLFFAc54m4rPe8dmmmsqSH4KhoQ0PLNImLASL8ufq86d0FPVglK9O+Ly0PAua2
wE/XJ8PD5rZvB4Dil4PKRL8Gb9CPOoFyQ++xr7dCmdrHnYBm+2c9aSNwwyp3MTezd1j4Ap9cnO6i
k1cqEIqJUerSwjyv81eeQ1aUYsyy5pd9z6W/BgEFh+rfjp+AEuIXKra9s3Y8qmFXBMlJwmDuQa0D
jP338RFFrNLIqDRRKxOfiDJE7J1FnjnIWgdCKPTGcXyHVVJTA1QVnTcKcmzmsBR9sLTebQR6/PwL
pLyhURlfsToNtGgvFggO8I3Z9Vso9xuCRajG6G+0AhRZpIIfjT03aEtseJM0B06N5VDFRGoNPnp6
PKT8W92MdhZ0xLZBOXakQktx40MQNkD8a8NBc+5dcitIWxz2jukVGTMQrwg7FTDlKmfAUlNID9V7
rTX77Qv2EDfxIZHoojEybfPLPp0552QOmucPJ7ndM4qMs22zOOiCv1xIbz7SPg/cuSnF/FItRGXW
M0GzAtk9d5QXgTjvzRlvfctdydHsUnipECyklfu1D1jAGh/OvivfE7pK9xuuFKJKdgGnpvAUrC9J
ZkWH1woxBJfG3jWHviGoewWOlZb0Ug8IDXkt9TdjJXbHmmWDvrZ6ousfXHABRA5frxYXYLEUJwsW
f8Wnkw98bFrbyeDKOLbfpKUOxXonuyTowjlDBpj2r6EHICTm58uf0h+1H24JE1DiKrHB+dljZ5uT
ZTwTn5ZlW1RcOrlWLUcF9itDKqrsretdwSLEbZA9oS80OgpeWnkRbo5l4WTUFtqb+lofOB/tc+cq
j3HyA3zvdpOtC1ntBUzy7XDj5DDg9fhd9734WZiTYGiAZwhgvhvHEHmojdAn1YQlyzomqjSvEdtt
eZUqGj7NSW7TkUztEBaHZmBsaTNHdbl4ion1cHAOqZxliLPqVRYP8NSkN2i13be3eAejHWGCDS70
/RQ01gp4FOoTMApRxsutMZcePk5Nhs+FJO5p09pbEJRcvXPRRj+KYIWOR29G6EfW+GWiXPbdG8sa
Y+4COank4X4fUUwC+vzu2Xr3r+n6PZSJvf6mKSKcGl+q1yi3/cnFhoYINPWm9I5Q3zOY5sZPx2IF
6rHVpU8zvNnCxkI803g7w9f/eOZyP9DGhH1E4QjWSMCGH5TJgI1Ra2c5FTndcdwq5bWqzjaEDism
g5xd37Wr90XTzZumnvm6L8ToCTcgRjmSP1T26iQUwMlx9EBV8DYCn28v3uPPaF8Qk+a97fZcZrD2
Z0dUTyd5WHkRyyyR9q/rNi+HkXK2cRVF9Mhl7W+UDarfOCfT4JCWcGDWMRWxVe603SEGv/LX8ZHI
iXblPcaWuX/fR2KaBo/b4JQi1R31mk8O4M/5pOB7OqDXDZrzCX7cnBi2cved6AzJRwXtoxBw5cjw
4o4vNyzJMs6ToNQ17dm6uXj2z9LF8G5TqVDxuryoTeT6B6IpVLgbIQ4ZnXAF8eUSLCnGAbEqSVIB
zcSyc9tox/XE9+KfFhJuZb4akmDLOwLqBVHZHIUV6B3/SsHuFhuUoOhCr90QfrXsF9PLoZ5dOLkD
SBBircO7gnAJbmfmpUBgljqJ34pXlXU2C7jOHxMCDmQIvDbHZ5q9lymTEpsnlXmwp8JIFiX1iWxD
C3kVK4oWWMjnvpFxUtyVbysTNOjw9A0RpGVKQkK1xzw8T2EbOVhsz0dbanrxiWedFZDoik4epYpb
7PmM94PF3g9m+AI5DGHafm4y1mckkCf2NwMKvUaL7OMKkJmITNrUMDkMVp++FyhZIiMc9PP1VKsI
zDgCNlUG4joKIMoMlsElYmJEMCIv3QmtflUicW3FnPB1ZgctPQppI+LsbM1ufvj/h3tU1l7RnX/X
YKoEwDCOFTU6ZmhwJlUxSy5kkTVIkXvGDO59e0iamPC7st7EGffYnfQtUmQ8G+pV/MJQW/0zd5iW
LotInhs1TrQmSNDzBehmiK+dAXglyp1CmTKqQboBTCkcvlXTiCuXymD15tThSnWjtKaRGj7Wnakr
x/+hHa8+zDGjPeRnCnQPVh4x4ESCl/klw5evoREVncioDVrrcfqYLWnyD3BaN7qlKXxke6xZ4qKO
66K84S13Umcod+VLjKWf6nEJ6cwplbf1MNuHv1GwLG3bjL3JOKUR9aDnR4Wdp/qbnLyNwATnSy0d
Rr3EnxljI267n7wc2VY9AyoHKZOuSCOJj4i9dSmLfw8kA1TXcgY9by4pIvAdEQmvGt4uUnDrasIX
iH10WVi40ktZZRsd7InVv67n0jH4SVQwIxE4/1lcxbh3FZj31eGbUoVolcoV5iGB2rgJz+j5U8PT
W38dT0wtNrjCtG7fG9iafnF6PcUDi1SBpC/1BXjLEXdGm9dXcp7WpIedjc4wPR5nyDS9Qo65bjj5
qjmtmW4q+n40Bjax8EzUZaLeOWFtmZXquxot0Wl1JmnaXz2DWNGIMaKNjX2dacyLb9gtixplVUSf
DF9yArldhcOFQ12cq9ALb0ChiF6GtzOyvNPZScrtt9YKQf6tpj478+fZcT+1f4Kw23yo3Sf07kr/
MjoaMvq8tZ0bMILJUaiPNsPRxCqdL2ru756+lzh7GzpeFNws+j7DLSDDXbi2pOj7UWreqULajsPY
PRbdPAky2ZNkR3xChFKP2aLRKGxpi/YsOv6znba/1loqc4w+Ri/2YIwUBfPeeD+YVTYGsuiUODj+
j7pIiscvVfKTEGujoTsw9SOmu24swOAPU8W+YWgW3ki4V0SkSR+UEKPjjMPDrS3DWjWPIm9R/Ucw
KZdRksaZCZpvh83xYQeEdttSAmT2B48FzjfCDY1qt7O4WGRfOrO6T6NEwB56cod3ECGebXNhMZZX
1//4Y/TI2Id+8cipF4061saR7yxtDb9mFX03LUMLc89QJoRvkNW/ZDPa/ELxLKendqRT/g22kVpm
nQKtVDljL6NLo+XyMHPeBjZQv6REIFi58MllVn4dmqigsL8u9ovgYausz3ydWg/2EB5SnvOUyS5q
khhg8l/mTvlo+pI7kQ40qDHQTOT/WXlkYG6JG6PHRkgjc5bZzbRZpP9ZkPiKxiePm+zmil0FeDnQ
6KALGhxqZZgPzcqSWD/2t8+ZiGc0lkf9kbVnB1UPpKUNc4Y7/IH/EkEn9CQxAIRlx0bkxul5Z9f9
Zkg2TljRM7yFHpF6VUJyX/pMjaUrSYs636+AmmKHeF85P32/bCmnzqbe54zNT4LZ2+rokvkQ2/hc
iLbe83fmP7rgKPIxiKBzdYNrFPX9U1CkA1JT5Ws2B8+S1dBWTmHs3GgU91goygbxJnXv+8flJ9lr
NT26v5Qte4v8g9XcndpAyj6lllStrqyPrDsvMPAZ+2+l453Ximh+BU2E7EAt4RgyDPz6/H18ZrZx
TWMOY8lW1UeI5TJp0nL76R01sCF/g2VJ5MyQE7rt+0smRyZXLpEr78/HA2NSx2fliNUb2x95mN+s
RZh2cDuECPnWqHmvWoPE3/11z89NujpAUG8cABIs9PDZoOs3+i96vbTjFMSQaJZvsaOxFBBUPG5u
xBTzgkXRE5s7747CCIkTI408XquNDy5nvMSxPMs4hsDdyfpszTV343sE3hcXGSKCVE0xNY3DMd6t
tc0iMXQGH1d9cUxbWresrVVncZnyTZjurM8LYJRu3DDnBY8fYnnpSThxtlHA4jIEMwisAglvUFs1
7FwdvsEUeCwSNg60bZ4R80krlVl0ZksURvjNjmacu9s71KGSYF8BVReVWp5BoZUe/7sQAvRyRy7b
OulGMGfC1i74gHvKU9L6Mr7vdgwUvMEgpOoIsFiLXwBFWQGWp9zTfVyNBDSsjYD1B8xqTky3kfvf
8oQWadIzoqS7jyG6jqfgUxJB//azbj/qRd4xFoOKEAwFNdWF2naKBluE2cqw0oR09yw/md1s4mEp
IzZQwsUk1WF4hnoWDJPRtYIyLGzRoKjxXAycxa8ILZJEXDH6JVDm4h0Wm6+XpGzGap1Euh8HbY2L
iRDwEy+d84xmONCL0Gv525OS0eZMG+XrOp4m+2hRnlxj03Si8WF6FOYhYG8LfadKYx3f359SUhfw
Sucy4mxUXDuESHk17Ur/oE5yIep8QZii3PnC4k6RtiSqxPvOMwsianK7UZ7ohnXh3VQlqbW5RyeW
Us39dE8bJL4P11VSwDONqEs8N1Bx+U+2K8lc0WjgVubBwdGQcSoc0VbxMAllR1652lNuQPk7CakY
t3cSqZCTGKYqV6OhSxjgA7AlxwQ5V0wBjj0JeKkRa1fa78ZC4DKRK5G7HnfVJ4XTeNY+xbUVETr4
b/nXC77SFFvfNXHcf7Gpexhr6EGWME0v41ke/PQuJu1VJO216SURJlwhTTjJxFdN0N85SMMwhJBI
9PSokgQUNajcikj0wyiklU7jJcumfaGYquUJyjSYgSSe0OUITRbcLDavI4VdbjlQvW6Hv10h6dM3
LrOLqmz80kAKMnWXR1ZwZDrUvDA5s4RINx5LL43yY6VzVEGFhBXt6wi6uRVjNjQhigRpFjjCik1F
tQZhYhu/ykJLjTXWOdrNyPX34Qd7Xaw8Ho5HkfRL2BbAwWD6ljuem4VKQWbL+Pm5wSakhoAvppzG
cs4xPhKBOcBGhoV/hSX8g9U7lcmfyONknkctc/IDevoz3bkuGxVNd0G3d1WjMEAz4S4/lEwEbSfe
mVxyoTeT9zE18uIrQqvjx4umDaEv6TooP+qykIFidlCZPojqMpeo2gqtT+8owWQSWAKfdt4bP9x6
IvODRQRFePbR4MYcZmWhB5+VIqS5oyBiAuIZXb/aci5g81S/cbRHmYgwT8sZYEgPzE2LQaqVsikD
I+TpSlEbFYYC0TpB3oB3q+V3jzNDFHLerAujLE7yN1EWyoebMMDw4qHvI1gQxU0Go5tgFimh5EU6
C13PSVKucvQN5OJGzHW0kdbEXdHzziVQS5+y87ySif5hiy97higmhA6qXV4UNmYqQS64i5H34a+J
j8trWXVHzr9CeyJi+GJi5SZCz/L6avbcoyq0y6aiTUrOz1VrTkqV9DgedvxJuKQVQGlxmhm3OZGA
07fZOPXYPZGiquYWnF8KxrtDOLJtoTN7CzTJjQGbMASkD61IDiPXeVzfjjnnt2duYU5ek4uFJ0LM
261kvXzKD9KC8qjTHyD7hcxQzg7syEqlZuFoi1TggXCKZlaotUVa3y57TkN7pc9AQWTobHTV97cr
iSPQ0LO/vO4XBpjzTdQtQBG39kuGQkykOUMltVemjlbbSLG94fEVwa8eGLmjjQgqCY/W8QIR7fTa
c7Je6X0SjwNeqIpLJI7YQxr0/PWE6cR1ATSXycBsQ++H3H+a0xB8B0OBVj6lCiay+QuIIcZ5iR0w
vEUCbknIuouaHldJy9XCHL/TZ0YItpPIuAFCBqePjZLEu7N5l29n8uvzHwgMT00Rl6rfBj4T2qRy
1vyBRY2TdL5vjHnXEF7OSwQAsnJNSaMVhjRkqVTaGec0paJr2MNXbieRtmjEIwps0mAFfCxc4jfF
KgXltIRC3FpQjKPvcUExM/t41Q+WqPKlXMpHhYMn/fENgtNe0RRTqJDD3/2ynJ8k3Y+Ps0N+g5EI
gcnWDCWlNRJ2DVKN1cLRAstEWVTTe+S7CsaT95/7gZL4vVUjBd9Yg6pazdtZmVcd/9jysGDq4xN1
MutPt6mU2GOBUVv4jvlQqb1PbzyWD3SJEyAf7005KvBbfsL/43g5C2UHuesoTn1Dww94Kk16KVBV
FfegThYcE6b73KHlmETpGrOBJLWGY8HZBllbBB0OwHiNh+eR3R4ehuOWFQRYJN5Ai/mTKz46U59N
4OEB8782EONeValm0mvCAzShKOiy9E/qE4Qo6nr51P2WoMRHmU88rru6Ykh5BMKK9qRnluixT7v/
rRTq4WSM9qG+H49Orsyf7akH1UdCSI57kMFJLS3wi2PdCjuHkW3df7cice/R+olsBgld6GZa9M06
42uN+38IBrogKt5x88yeHwK3m/cklWffu4iMQw+Mt+RpEsfiqzGrVLwdz9YWddxqJvBb+nwOiIu9
9paxjHznx9RyE39V6O+8jIg6teN9BkhsQWtHjg37O72glx+oL84RTUQADi4ilqq/odCr5sfAWI2L
3ebTNLSjkjQWjteQx/otGtaeprQNnJxB39qiRsKet4rEIRBLDCx2ageL5/MtMz4IfrTcgtAio6wl
pVcigudFcfgNB/AnJ8lWRW5MfYMb0etidhFnyhEQkLgj1MN0gz2O2jQ34junaFTP9t1J+H4ussgX
mYfvKQmJ11+/KneLzQe6Hh2Of7R0RP+gYWmAd+rM+XBoDHy0zzyDXuqGVJWaRWvPYk+CmQ2gfKOE
5VBmx9r4xcQkG4hlROs/21jCJK4S+h/0cKdy20fU5Iao2vK1z8LshcWn+w4QEX8iyKnyxwRyuR0k
H0aYKquhEgghh38xoaaztH1Z3UpX7r3es1cTh3b6/Hzm26cXz0PRaOpSCTQ239QFBs5A/8cmyNrr
hfNPhEcpOGFTZOqdh2aUOpOwYrwEpvvOCa2orY76PW4Rmg//d+DCMS2gKTVxAyqIoEX3bUM0ZztN
3DhrzvouxPE3b3yz9byqVYFIXIdXxpz/CRGikKoiXEpHJGcM/W76mkDy8TX8XGBmQDhAiOmR4ckO
WuLhKyj7BglPjA65mH6vVdrbHhj4mL8BKpuKMwTXEjr3gFx/5pyMTOd9PBwsMx/xEtdi3+1Hrwsg
HHwPnRfVUeHhT0LOy8cPEpjyyAB0T6483vWYiVHh3xjIl4lOdL6sM1NIVoZWxnY3reFsG1ak3OaM
tZbXUhdgZ3P98JSJ/SPpH6eC1n5ZlVsa/+ICiVmWpd053DsYMcqW1AadWArDwXo1jX88LddOwFeM
8Te3AQstavnGv6SlbgLVuK5YHLVYnZoje0a7mShpq9EZUQissZ1vD3I8pAP1NMp4bABc9Bwhva1Z
wM36GFY9dXamHIsK/uhmo1+MTLtvRXNn1YYuUTOGtu/z1cG/uLSWYTrZkxZDv/aT1nxe1hHbFMKp
FV0HuieSDSrGsJoULnQ7bFlFFQVCNnfnOf3CKToAbtpzgmYc/7+6srVuOEVyGiMKljmp5YySFn5S
KpJ/FxHL8iZlE/Pn8vmt8mp1o5vyuOb5CQyQAEcNkuQYsxeZYwkmvUBqniE+z64c3ZiTWhEufs5J
XIS9aTErJVmdEMHlfR/FZINLR3XQADysTUDT3aZuqDHOBKAHI+EeerKWxaGyhFQuFuu3WvyHDdXN
Tqn9CzvgHpKrivUM5i2I7ARqL+/D8htJ9Ezl60pv5Nl2IC72feLfaqcaOAJsPi+h+rshV0ZksGz/
tiDiL2/9DEiCfvXuTMAx2FFG5lKNwc33LBXm4ZJGQepl/vANnUmI859KyRTMC5GcDCuzwxESLoG3
8jizH54dAnF7rKBHO0Uj9ImTuY4ORI45vLboSCYUBUMI+TO9X9Ne0LKy8qMBsbvzYr0ngwjnyEpM
qWv+HX5UhA92QFOva6ap1fO651TjbNf6Cppb0YNWr/jAVdAw31JzJDOf0jV79uBBtQKOrhMT/IGM
2LP6gE3pH91xaIeTUAn6TvkyGlND/sFOiHfcq32qBNReaR/yibN/wO5CTu1ONQTbI2kHoyKholyG
aq0hkYVuc+fuCaOfIvZjuOgPa3hGTMpsk9cK9Mrm6dHTwx8pHgG/ldlIZEyU4Rv8Jn3tbaG+7h8D
NGvceYCoZH4RqQOgur+Zn4HmEcp1Rea00dgmc0PRXUwpAj+Yjv4N948/QG08pQVolkiCYUQwyBu+
d4KIXZCb+wzk6QNTWsQkNGwKQOjO/IRTg3mwCo5RNQ4P1BLRnqAOUyIumLDNoHiRL4IDhy1Jc4PH
o4wY6JqDAqbF1ssBVHxh+AS2ZmelnbcLN4LTUFRCFid19/pxh79VNaNlQEzIdHsEq/sk7K+l+f8A
80L1HNCYddnNzMOuOponHN0HJ3DCgGyG3Edl/lH1gFsClz3l/63h17/Az/aGfTQxVYAjI9j4Laln
vBCm3Pbw+xXesVs2OwOOXw2SIwxh8pvFXNPQjJeeTw4HD8XKuHsa8/5a5EaVZg2zW6mMp03pm91q
tWgTuBVltBpezilJFm4SXKsawMP+rCShocI4goXS2IAB7ovcxRpepnfSSTB3VEdZrIyFckb3YIdQ
v8AjZU1kb0dfKmxMQ3f5SJkLUl+ADYeUpSFlnGv1DG3h0/pCWPHxwWdT3cQkCSNXYsoa1wKfraC9
iZ00hy7fT7M1baV1ojREB9kWDoTQQx5Z3j7rfW8qftrR7uzdOceIWpn+YNTSdvrIUjY6+mrok+mb
JswdxN4dFDsddTIVOoqfn/zKfgGc51NNgv/KxR1idGB+KsFy/H9sSUP5CrB0co0nBIXzGO26OnGs
6R0bjrpn4XMRT23qQaY0QvkXhgRvP82LNFhxcL58SjAbMKCvhG69VmVn29vaOc6bOlJZJVLQG5Xo
sf2bnlDI/e9R4oq9lxZMBoCI6LDCzzcuWCl1Njv1Xxg3mPq6zI0XY+Rj+0w1dtlD8c4VZGOxm1aI
5B4heWVxBH+k2lklZcsuuj9Or2ixwmtxscey8Biw/920O3lOdFY7WEDEG55jD3lgSLQm6T/J200E
QjePPV2M3tBKrG1sqG7onA85K/YwUI15bRcYR7uBi0U/sVKk+a/9HnP/pkxYKLGmraMEYmFg7vOt
EGwBmi+tL35oyKEZ4M/CoSAD6sASIlD1/curidlw/P1OhUwt3Vcyz2DEi7KD3JNcFegGgRCa3uZl
tspk9Bn7OlaTeVYy3a+F4uAPt0fmzxjGAZKJCZRmQiPiSAa59p44AsBiUtMOn0vOEI2IqlyhbqB1
Jfg7NwYAPaKWyXjoXLJdcxIpqvrfF59Q0NCmG4Hvj1LIVX/8rDHd44cpH9zlU2wwU96jsb0+GZft
7YFEWebxX4bc0ZoXU3c0ES8stI92Nu5jy8bLWSVreCZSMnIm/9q1+YaYlT60H9QoS/E4L6XTH/Fz
MhTd45GXZYIHJh8NMRV0axsIoFLIdGXNSFe1gUDsugQTV+L2jspEV+ZecEGHJ+54Xe46U8+ufP6Z
e9wQlu5EAXa34zivtnNq1mqEMEHvNrFH66jVh2vSD6K8Yilg81L9i823dGGtnXlSOU06zsMlivez
ec7r9H52RbuaBL6YO7iJ4Ea6BhUQQ95F8mnLEF7ALZq/ch2NdHjTnchdhUxrNWGCpoOTeJIR3Dxe
wIL4SD5XHD/igWVHCAS/g1QkO5JzPtIb4bVCQ+If3Td3d1EG3rWDao0GXB3K2x1wAnqHrsx3mBTH
w3mGON5rlTSky7EISuB99Tan4FGKR2ET74Fap1rBHa3CUyq1R+TL00MIdeOwOZnElRfzU+0wYHST
yEeSYjczed7rjiZ8Se6q1Sz6clBAeP2Y9eUgduqXsbBAqjmH2yuShe7DVnqTnLIFjqneEcpn9h/U
O1/JnksThDbLpF2AuFJWpa6MAcfc8XK3+yzg8ynIubKgCK5w/NCvjHlJUke6ey6/NJH0DRIxNwpN
6U4MIHZvR59lijbnSJGak47kYWmXJKufqVREf7Fk7bRc1ELqJ56AmVmQd6j8HgHV+U3VlBOIfvM+
hdy5at+hmR3mkuiczl1ZBS2Ar9SitAvNqfdN0XAUJ/uzOzypIQAAp652mhrviGeKs92mqw1yQ3Pk
YvreDO+QfAC4uv0KwNU6VAInamuixEDGJBXiulEy4ko0uz4fF951lJTTdzT2BCFfq9HVgEfnqxwY
0izb0vJzj0rbJWUSaayEXN/qms3k7x0AvliQRDbMjyZxKPp1zCAq4DIE6T4cGb2Dy2a3fhXvwHiW
WPyiDAko4bDPjfGEL5kpxTEssfEZZxALKPuXs2PDW+dhXer6epOnqPQSD1L2jl0eCp6JtaWD88Xx
nf59eKzbu0J16T3elznEkict00ZKvUgAxL6YcakIbnPER6iDHz+zTq4HURd5DlcZUfsiR1QQhlmq
KKB/p91Z8rT5Q5/bhopDPAtu4TC5faxT9ZqaEp7w0UaRRSpHwejsyBRb3+G0dWPVuycBQ5/H7Is8
8PuhCPN+RahAvkis5oS9slKZDlWFK6xztqtNw3gkEHlGaLUO7DoT8lxnon0gAjbkdqlyZms5TPie
t8kmxlEJUxhJMqw8N1I+jbBJgok3hJ0lBdYs8aBdRZqjue4ZRilx0lahV+0Hhne5KgrR8yJxQ0ec
74Nn4B9ZoGYbbLr1lKH4+4ahY3JRdqm4RxZnIxaguw8N8T7KmRq2KsPvgK1ICoXVtCRZAozXrLcA
29+zMC9iEc9bBmmKiTQEDDDaN8PraeviT4HmwkPrNxcFwngrhOKRqSVPyZS0U3yt+rUKyptlte+1
xdIViGcM2Kxaaow9lR1Zz8T7Mc7UFz4LeRmYvVKKEgalJRzoQOsxzwGV6K7EH/PBhYkN1gLf+pjy
1FIbdWc2Icr5fznrfW3NpQYiOjmfuY/0ncycZR/f1UmgEavgn8IFPaBtYQqxXRXnThHhQPvN6Tzy
1AvSh3M+KAP4AK2BpFIdPQCZGDqYaC3+pxwgvdYNFikQn3/o6KOtC79LL/ncn4Kkrh3E04p+VG9M
7LzlsDIt0iRloI2c6lyhF5vvI68/fqCQHM/jN6M2PCif6rwgKqF44Ih+yqgrIkaCMk8WagPeYCwq
u4+bdXd9jrMJMvoNkQ+OK9TDqi20uAvIhDy/yfelMe0NkXtg9/Oh2UaGogsB/w9AHY9xGMGziMcU
1znVHmKgb5xZT7itO1uRndh8ttNTjcFeCUvtWxBFMDCO9ipBIfO+oFQtwIW3pMytQmF9Te4ngp0C
W4kh2tGYJfu2LtO4phfF5QyLYNfrLVYdm7ij99Eo/+0tFikx/FgYpXMClT+73FcanBZgBZnUlkaH
Uf++ElZMXXp2r4R46J2vwnKyUpSUAjlD0T31zs23n4rDBnhp2TPi8y89DvKh9BHZ7Xxsn12aULBI
jo0JdgAy5rSuB1/Ht1c3AUEEJehsw4E3TE2zuT6dmQup9ed9M+FcX8prE+n03CUJMMDf4O9nJC/E
MVDKSF1LBAqh0BBedAkeGkBA3Vfjv9FFvuGeCw37t8usGAOljeVqMGiMJ9BWLFmBpVRi44Ev34GL
I2nfP8YQSUdiZSofyE1AYubqoI5WuQtaJK7c0cj8L7nPGdCxx1MR8ck8n7S5Rv2B+KrTbrJ3voCR
iwkn/B7sZ5dA+z3Q93LQYAsZ8QHuoxBRjLBnwjo7v8nxwF6a3hE0mwVT68sMcxnn8xz5rsfNjQ0F
m5z4ORDMW+21jUKBnndCMkSk20vn/QJi4GBgIyqf8GGtqoqbQi+JmDTE3uPMEj19wmsd4fEYxIao
UZilXdEKAi3aGbfAKUK8U0S0Rdu/K0VKxAsBA+SlUMOTwQfeKnAvLPWzo2Pjc6k0+y2OobyykWbd
jYcXVibTzLBDLZpz+fbs8rUeXglyGovFSO2Botr2A6u4ND7ofShi3mMWuvPYSPrbfItwDZbO9/3v
OKfDStqdFrZHfXbslfeeeZijWivIBVk0JG2m/5P1hubcfqxi4Je3fq0Qlou5ibUTaTMUDp8z987h
/uVrPnGA1XhIFwVVRQDjvZoZCNuXDdSB/eEzr/s0xFjq4X+ofFBBoX82x2RBxROZYXwANA1HeS6D
OXBGRtoxIM4PsHkXehCxUMC9kwIglOVkSQnh4bQl34uyOvwwLuaPQyWvd955zKdbsk6hzxqKBki+
rDqMR/LGXbP8PyIStvLYmGhj921luO05GhCV8Qz2ywOtktEb13y7y+iEVfwNudPaLm4yT6MBw06/
F4gw5tj6d3otss3NvVADtDyyVb6NS8O6qW6+LMgNLSGQp0YIEsWZYvNGEVx6Ke6KhUPgrnI+Svfo
QwejhGBC9qJDZn1RCTcIcqEZzu40fAvCExQwLcUrSsCqjIk2d/ndnjjW1HtfW0KOFnqTYYVP0ICl
aG6Flch2FygqMR4Cjy5LyUs7G8z1BfuT8d2YeAXRKoeTh24rcFB8tbAPzghGb463oXf+iRDQzCCu
sPrq2YRO+DfskA0MYHMaDD4HLzBqn2NAjOpEgZJowLJrmhotONGJZa4HLONILqX9yBZeHBCODHK5
NNFu3KoLqkm9ahvkh4y7Vy+JVFKGqY3ll1dZkTQHSUui/S7Wcbvnw1XcLQBHztKRDRnuznMS6IpI
x75Ba1o4uhhLYXx7G9JNDtz/71rX9l13nOkm1Cr+49T0BOW8S8EhvCC0eh1eAby1aCpUo0iEpYCF
HAjuQ8Jg9qUI9jLh1blBSCJjw82ptaujq160Jk7JS8UheIobzwAyogkOtd9awTSAF+Y9wmCfYOVs
q//0m1ovgbpK8XYo0CFtDSZF+sCk0cwTYUxmdUQ18oHBu0O4aXEhA0MXN3vBF2ljSH7O6WxtbRD3
vPMAOkn2U2xH30tx79+UJm0uBiXLxurd7farMaUlL+z9aDTWNjj+e2zPJYKW52BzASuHTwUrnyJ+
y1CH+EkVcrZ1TzS/lK2sQ24xn1c4mstnPeaedliy/qFhEs5gHzWWrwXAev4nrGyqvrZ2S7fyjzJU
KX3RxQhq28X7s6lapRbjgoZJvLGi9pYeoBfx8HoTdEbY+ABA88JnoZmxQFXpC6XLG53HpsbTdy4u
F3G6jQJejtBq9xYjiWuyz5mhZ03BCuGz+CN2/B1xYwLXr4eove2RMxZsPlwga/8o3gmsNBi/lY1m
iccD5Me5LjrYrYqQiI7tJh+cFuQzUmEyvrLUtHBCHRsxFOOCDq2wRV+KBaX/N5K0LNQX4EaQvJ7U
V/ktL4jV2kKOMXO1v5rfEdtd/gK80Lx/9m38jG4PolzVRjedLi3wfXG7n480OuC6t9TCVWHe2nwX
p6Nca9ZV+iF8eAw6kaygTXw3GwIi3RvMClNJPADlLOlqvxoIYD4QjNpmJuYR25CCd5U7OsLqCuvf
ZH3sFhiaKOLvbLimv8xn7F/FTiPNJGEtSCCinHU+vHjba0XDj4N2HVPWCo1T5yhVxUGBVX4YRO3Y
yFdlbN1Jb+0FBy5jy1mjoVEOomadi+hEOxKbelEJxOeS8/v5Fqy0GS/jpxCwtcDJa528p/LrKZlZ
uQgx0T5fWW4D/kjSeQZF/lk6ZjR27w8ZaPU18pnufRc5pylmrkpIcvWm89grPBdDLq+C6TfTGlZ2
H5OmeuW8w7unSySkQ9yndsX9CYcNEl7ZJGlsduxKjZKcAGuqT7knY5/HmhKJErXr2G2hNIkvgYdS
K7vw2wRWnqt+iJU1eJhoTo4RQxYZ94lwxxWsaSw1f1HcQzOrRShY8YOyxTPiBgz3yJsJALLS52qY
Bf09Z51OlTrsTKw6SkUiNqbUcD+8TSGKkqGuafHeV2jlIAcfqN3WCgS74d+Bai8odDZ5YhbnQZxx
nAWwWZuE8J59f4y9HGVJ5U/6wufJsz0guLsseNjE/79d2Yyi1Gifh3TC4g1js89iANxlLYQ5KUn2
PM/+Zs5uFwl7m+JdwKFJkc2sOEZdZp660jOfJ0McFipVnUpGLHo6fNvdbr5ABF/Ej9zEcld7h4r1
+6qt3/HctbV+s/U1zUVXyCriDO6T1D+oVpDU9sA3zqB8tj9C1TeuwQRPRTQ3J6FTsnP5w5mxSYCR
X9oWHkGInhs4bgtUlpaBQYEJKxZ18e6GhFbhU/RZR5ZVf6H8boiCHUE2UudQ7e1ENwMXFOPu5bGQ
sabUQBRhXf/wpinX1KsyqGU55x5YNRHQcoydnKP6MUzrfA3pc0/lqshos/2/feI+3KZZODpme7Oc
93pDsLhjgJbpmXTDYVNyj0/ApDNqFP90JxOBgBp2weV0uZIXkZVfgBgVbx1u2BoURx1ARg08u93u
Hzc5E98zICMma2T9ErQaZ6kya4NWOGIGhTmSUiH8pmjSGyrNP57/jn5mcFxbmFof+a1UmDo/VNyy
s2KANe/Vwy4u5nVO85OW069LjVQ0QSRtTBxZfEoqodXZSSOBKA5tCfGJzrAWE4xvtupfsnq6I5lC
3wdvqrzj61IBRMbp/JSJ7bvpWl3WA9g7QcLieexeTxmKbbDEdBMjjtEKbMxPaaG/8EkvBoQFbY63
f6JoLbX8tt5Ywf3ouqBCc5Qkarefnzzi2wPZdKWJQwJg8/zC/SToJPbCcVBHtdVFEse0fx25nguW
nwL9UImW3pq7Chnq0urzlKDUpXdS6vDKSXBhrfDiWzT5vWLCWyNXrJawSIDLCC/Uiw2+HppmGjy0
Ow3arkhVxITt/JxY9WLfLJEa6UMsgz3LqQvjnnLZJLUDGrmhrKhIVYnbZvrEAl+PuIoRPQNneRc/
ATCxWQ5fKhvsG/MtG3kFHw3iQ3Jm3SFwQX9ad4ygBKuZpg77CCAWZ4X7qaUnYIpHUXBXtokrqnqP
pp0y+sWkGxq0URHQJNpKwW+K80TYhv5Vqw51GOsflUdtS+ak714S9BXlJeNZWMz4OeT5t5FKrMdD
5R/YpyHsCv5UOWMKy+GeV8s17fDqXClEEtIn4Ae5xeYkmsAkDAhTqeHRMfbA33Npc+VcaeIzqKeO
AafSJi85HJYjdkS9a7hBkiqH8zf3gRDtIzhkO3EkvOkWsvLdao9idneNgWwDxI22JdcG5yU+o4yF
rSn/OEQfjKNn75HrNruSxbcJKMlGN6RqTB46BUOwxVqxsaxLuzpcIEiR0wiCFVX8VvxPxMe9yK/x
vO8MHyGZh573L0nXyHY12BRtd054ZP3BDMSqYUSvvER2ek8I2hvFeg4BgrLljyYyzbwEKLqoQ159
1b3W9dcF5Zms5lssHx1DkywwNAgw2FDx7dd0iWaY7FFCICehuY+4nxvGXvaW6H00NtchFkGOmWKm
kjeZipsVBwn+YMq3egaOfRsAWmcXFyy98RIpTSLRNnLBS3RIIWw7y5vI6qJUI7s/cNj45rmMC/3s
nslT/nNmNGMX5CHNr2vStKnDMMnTD5J6EKV3i4fUDo/QvSMh6Bjl4WKG1thdCQfoOgejPn0Zua9c
90SlS045pNHiUqja8PPoQyQmM7Z1pRwhl7zU96T+73HJMseYJkrGepe94KrPL8l7hsBAwaNE3THO
t/YhHm9iaEQaWKFHzw7lvgX9DEg4OdVbhHrEedo9c80bGjWFwDA2QpF0fu1cAgUILSpSkHMnBpD+
zQZSg96GBNbRs7QI0B2TLJKGRDYZqIWMKIzE9m68F9qqvTgNzs6KR1L0tua6cpu1XidDTgBtr/Ab
AS9DPS4vtCo6/VexfquUU4XlOhTtKTifFI0OG1dSPUBfWA0zY9QKvpbTFDdOUY2JlQeaJpysV1E9
WoRyq94IZtjRDe7jnkK8YGRsDuj1XtdxHEnHQVXUvAEGoXmt5BnX01S0G1OsLXF8ZDUiyrmpJx9S
WXSnq+stSOOnQA4OvdiScOOHQnOxlga46QL5su7gI551MvKTvRHxHe+GTrl2Cg+68V2Dr0BRZbc/
Kh2thEhMXnrWk6VTgK2hGWEBR2SepSf0O/xWp0iX++j8K852GKkRuHVnGZaitXXW+oLF2FOX6LLS
Rbv8ioFAFqEzPMCsZrmMNEE/iRCD5W6QPpiBuWdkWIvGFyKer6G0/hZXKj6JjYDrxQsla2GWX5qf
ntl6+tOJJYB1f+quxRyyfXowED96RgQLofjkr1YQwlCyuwDGw9Ng6MYnZOOCu1qwU0FZLeZ+GDf1
7wnRHjobYPJTYKIK1MoxQhkmm7YxegmFAcOANHSmY6nwj/gLSElzJmR/Bi19NVFjdQ+efMhl9isL
YjkXsceArhTWHeEd3A3RUiml04QmTt92eVeeQGOXxnc9IHvUX5bVbQvkVws1K8p2q/5yYulNXpPI
89VsJ7jFLfjM3qL9i0j/qGjgbVjFniDhh5NWUrr7GwUZyMsr0Kel37pkm9I9tblyJchtfdoyJAAU
OTjpwKtRQOnzA/af/ECYwY80hil1O2ScnnP4mtvomtvqUzaxSJlA5OT5QXmPcxY7yVQrnbjz0Q2r
1IzM+5wweIzUaFlKQd8d+MXmxAYcfWHY0EO6TtjLibCbkZBeVR/rZRJtg3XPdcAntGtBQrUM/c9S
3PEGw8DXMuiHnJ+kSNuhRzshLw9QQBisX3kOQ4dpmYsabssu1tnWPXYaFvJFCl9/mJljhyHzH5Vo
nPqSbSCSM8efMRR8pDhamAN2jnhh/fXLF8nmVjMK/FfwwPPPIU9C8S5EDDGNnZredyr1nK1H5vo+
HcFn2Ey0+KjpZwrUmS6Ps2eZ9Pdw24BFL6FXu9jWeWTFavZbyyS6D4eI43CCRH+3nz9LOgkQEYxV
9GDTxd3L+AqjHsn43NjRQfK0XwOATAeQT6JrN9nMA+6Cj9p6BSEwj6fmRzD6o53VojRTgWCdhWum
608CL/gBY9x3H9HedVFythWPT3bli/ASBfsr1890AxCXMVSKczt30Ymqw7u3F8hwiUhtUTZkedhw
D2tcsfjhbGvUd/bhbdPiEhvpTrMKws+BJsXhpwSyAao0lbXVHU/M4fzxgq0kP+BeSKH0p3dmbVJn
E3PvlF7lE6aKjk6fS2XKN2+QOvbXiDyhb55Twg6OhewDxZmbqhKuR3dNrNqORZ/SDa7xxfJxFx8l
KJvy6xq0ZohzKcKq13bXegwaOjT70iOQFwxiOZk6zu/jGsiqKdRz6WbUpRRkTYqrmm4M1+OMMLjE
Q6r82GHkDZx11vlirrwCzB45j4FALwg3tXikmCk1NGsMlvFG2ujrGhbXvruMwbXS4f+dS96Cdq9q
/4ndU28YLyVJ05+mi+B+4FJCw2RkAp/Mhs/v2cmnZQ1eOuQVbkJqVeqyTRPOGSHyI5x+8Zetttt4
QM9oR9T4fy/hrv0G9d5ZG27jc+rEC9CCp9VpVKWJ8YdJwrBqaor3MWJPSrTqwNGzokdudf6nxkQS
8D7vo6cyAFKB+LA2zaZ40MtREWCUF4eIQgdX3PLRRqUG1rHJOWmnBYmEFdtPN2uFRfIa42isFG3X
9/M5C2LOsQOBS01d5xiYyeSWcKdFbRoF8fbIhx3kwzAhdnYfMrDIMUPd+RQtpjNvFn3PIUpv0jxK
Q5NCobujQapQzIxjaAto6fHBcn+Rec/P5Yp7vOVVeyArdoeBeHvBnDZ/6j2HHrOPXL9hNElOZoZi
/bW3O3SjVXBmwlt4Bzc9NpF0mMVlmHNKRgh7TkYqdm7+6nAABPsPDy+4M0ChDyV4jjIq2JLBepNS
wcNc0uo4qx6sNO4WrRP1g2eveJFE9KO4iN5EuyGTN72VLU++YnQC7zK+Z9RrVmOe8gvxQtiH6XiB
LHRxbjV1XakfwA+z53MhpZnOBHQHUlxApa4j0/ofFExoTZmlRCcchii+RNVG84/LCXNrUtpqGBGn
tP5BCijWYB6K7AvqHLwhEzp0nzB9l6UqVm2V30dKv+pm4bbRBfzEfN3dbr7NbwNHcvKPGEDFQB8F
NfhjTv+DvxBfol1guYdy7XM7IRUg/7BK9r7s+WD+ARY1bfHdqOocbEcbFMTTgMeGYznxewTogcCn
f/rcgPrEyqL0Hu9iW5jBGK/LvQrsk2ySUIWTHHUxi1+0NU0jYdPcJeh2HMOdX3snSo50yCTZ9IS/
thwLsQZF/wsT6hpB/JsMPF5+fl7TE3U773feZwduSLp9y3aDKRdP7fzxMoPb17sUybF2334dPA1p
fktEjkucpC4DyXaOJhsCRO/aCpBJaPMJe4/zFp4smkYlIAZopoa9rpaW9DwUyrFtjD0dDCIwLg3/
DZYWAsIE8KWYLnWwR17OI3Qd5mgr8pqigZ6Y4XyBl+bsEqEwgRG11o+DbcYLPZVlYl9rgX5L1vgA
xbAe9e+Iu7N0sb6sgb80JUJiwTPa47QYMUtM63XovRg4NrliXqWrMXk27kzUNTF/qhzo6H7Zu5vy
IKvU2plvgYUwgXZ9x8hwqy9x2/BHR7fQbPuEfHj47Z1Og6kYdiVakvuGjtyTtxY6Z/t0/1/t0Hec
yCuYBz/zF+XQ5x8TYT1nlxt+HMUt8sFeQkFRY++xA2H2Tk+IOH20Mgce9t66u8tGZ1G5m9CkFEaQ
7oy+tx7TM1cqWspV6GPegzbbWErOHtDgcxl8xGBSyQGA3CB9K9yWcHeNzuOrYIKTRi8wTMEfSf9f
/spwZPCkWG6rAvZFmOlDq2kjCE5nuEQux6bx0o4ZawJQ4D4RPzze7ZmXr45VNBrdmK9L80zueifE
gz/FYh4iNv1//0ekzgvv6LHwebLBylS1M7Ub8tG+aCgFgmEhZ8FdXTvYzu9482mmYH9FpG6+efbF
+PSQaXZN8VYuDJoZesH7S8HJ7te+rBM73edietUOS+w+HOMUsddLpsuos+du1yOArTtaRNiJlNEI
8XHLoY5Ffuhnm9UmG0Yzn1Ggl27rjX7rBNUUw/XSbaFJF737Sam0tNbi7H9XUb9pSizMccP0M9Ev
HNlPVMraOw7YnaNNARFjvPAt+bl9PN663Bfk4xO7J3h0yLea8x84vWj2cE8eB9iO1B/sdCWJRhGa
hk4iWSm0tGBX2APkez2/pqAhm4+7fEn63ZZlUtpYeUf4usXHnPuWxe/sgSvftzuwqzvqfssI/rb+
q5bPHWnv3YB5qD8L3iR7pMN6QG6mZURo0Tghps6ugKQwsxbtyzLNI6QfYXr71a2zKD0ykiKbGMMZ
C366DfK1JSRmW3NrlNbBQozJwMesYNt4tXJ/DVKdtx5TP36D+ev4BopEVG6Y+2OqFlJ4z3Y3ve7j
+kI2ZlPwce/f4NF5/tN6u+mU9qlXQl/W+13Cr5RRhSGDHqU4EEcnj4kWy/V2VarqU1ndrK3aNDkf
FnC7KClLfX8Y3SrOHjp1wFUhG1GDWd3RqAQVEhYGLU8HWPuNSLHqttshfSpHNnDNXvybPRR1iu/Z
6daDqw9n+E82Eh1KDLpmhwpX8pg/A4nl1vK2T3dXmy9e6w+kxqi3baCTRG/mxw03GYH1uR/hEt8Y
TV62x1Uv583htE7VsCJ3tvCo+yrcTAWi06HFAusVKeJGTSx7z4ZqaMFxcMrB+dP4yW3p250avD6D
Zit2ZN6x+L+RD7/ntCMllmkdkeB8c3Z9VkrDx2Ouklq7s3NTOouF9SwKy2E/76K5PJbsDHdo33jZ
c5LZZUjMqhc+queFab4X4iUkb3otX7qMg2nzfeyLbcjXrb9e2+oCv9NIFRLdo6lIbF22fdP9+dUC
LcRRWdQMH9Hl04k2t1lFT10V7Zx27gHhiZul78cjTBoUCIq6ff/grDB3tkGgpOq1FVy+rpi7WFmZ
0swgBH0GXoP6oZaaMaBkwxT7GOfAjphxyadWVgIQHVSD3Iokvpk7b86CDYt2A1sZU5skMrrkvZoA
yQt3wOSDOd+yJVe4S7Vo5GLz8AzctoHb55D3VzrdUezPV5oBhxN+UKNuc0WNlunfHs7ZD8gBitW0
WsF8sP13OoDOKqsaWgL7bWf5VWk2AQGhB0C7KiYm1QQ2LADUMHdIdU1kskNgJUcRYxLx2Rv1BoL3
uyQpiJyz6w//Css5v1RzJVyELG23FOHuaIdRdkn9EtMJqgxM3gqe64LU46S0nG33WbPKKjgfad2D
QXzFW7B+NF6nXY6d84NsBgRi7s77xsnWbjRMuOFq/EjVowvq/5SjEqdRqULcPMEQIUPyGpQ+Y1SK
fNQo7QrEO1aaQ1D72yemE3avEfT04VnljgxEk5vOg4bx3NB+9TfYYi+vb9r1Oxc7nuRAhKuEEUs8
u/s85/SSzhKbyVfjMB5KlT2vYBl0ynSieyiFOL5xWJCXyLQUcQRQEAUzvHCUFfeeb+YAStE+e54S
EwStesQ3pyYwHkGanFX6HScPl5nkQg2ltartP+p87UPMMNiv0j3JAiUrJGFu+7DwkcowKdk9ItmU
oK8eFUvxw4roXku6Z77nTw3PfAioavmve5PP1SoRaYLtvQGqOcP1lYo+2gEya3fYGbyYSa5nKSV7
PJN1RpwgKvnjMUTjtRyR72EwfmsU/BzJnZF+8vEMFjWRsZJ39m1MxSiiL9odGuUfeI+u4o/vFMBa
YUnjVX1dCczZkV19KAuodCG4LkOKifGAD5fEad6lF+QSmRl/cH7BdK7YkrwK2X/SbvPAZhZbpcNV
+2j1IDnqTi7sAoBmRKcoz7JJVhJ0NTXYEYkvsw+cV5FxBl6fbbYC2+OxI4MWTd/S6A4pjYJ5GpE1
SrXLNK1HDsrvlV4eg55A2BM477dJEH3rZ7ipmmLQIRlW8SE6u7rmPIt7ww+hND3I9FEJSJQ7xssH
fpkQEbBMKL9pnOBhwsk1F+hvuWiXjvQpvxzaV5o5viVewgmxiAGyRTagBLaRtIJ+vaIXa2MOZhoE
aOTyoWs459b3XJD8TbBVpdRcDGWsO1aQCv8lxsfBoJTpL5udWUnMhvd7BZPXSJOCfOMHzVb9nYxe
g9wzP6hmEiKOWo9aMEqGS6/NUgJTal6Kww3oRtRbveY5EPPCsx5q1M5T7P1paaGVlGrhrEAbriPj
lnVTSk89yfyhki9pNKgVXuuXoGjJzPQ2c49d86gMBhkjvPqY8wfXhrFgJ4j7ggZ82IbQtt78pnU+
OKSKPKVIJIKIdSLuICPWTrmXtaYHuB++CXSCcfhiyuk6UgXL234J//pDmgIMx2MzFC35nnwxgQk6
uu4t8CxqHRTnUOmB1z5AyUPMiz8s2pi7sm/Br0i8ZdpZiVTn5auQ2BmSIxUqQDv+0dkvnA6H46ZH
Z7Dw2p2X+d7yCq0fthFU7GtDl8J/u9skz09cAX+I9zdi4yoBBmbHXU+T6mOrq9p6KMcOCi8somoG
w9eK+0BnOyG4stu1WcgwCzCyvHT/rumz7FpkmfG08R3BsCvYmURoSRlbBtq1roiOWQLrOUYgKpcK
LS6tuyrOUmQDLg7RI7idre2M7OBk1cl+Kq9IP4Go6GrfCEmRcTyDD5p1w4HrQPo0Z5KDlP8T8+kl
LNHXRlIx3mvU1xZmddvAR9L8IncSKkyqOVNfBZtD2kCdbJOxGhWp2jKuqxmc9yT/aVRh4eVxLDHw
6/NULAfxLk8/i/Zi3SgR73zEgJQDSGs7EBl+OTVsq98QhfyGtiPY7CMCUbb3l83TaXdH06TXHmBF
liiHv42sU/WswclhTHL52hbfS/Kd7YdAfzZ/A0DfOr8Q+gI+A92/+vyuG+r9i9ytytWk9VEna7De
J8GoA3numniYs0BcZGMlmFRfEF3evWVfY69TXqve2D7VxvHh6lNSodh4u9vT+o93dhX9srHHzh28
O/ciYwlvCVNcq3un5lH5QzCa/MI+g2xBcKA/sdL9G57mKD55P0sumbt8nbijfHkdg9ZyuZ3KHved
pbyNTVio+xc8COnyaWjxPxoIEzmlnQnVAL4dQeo0lflkIvkeNnssBghAgQ3/OIKLVLE48inyk4H2
KS0ewoUkhm8Sg2KPBuj7h8Ch+EeK5LVy5K1J1wy0X5EuPmSFNrxeZPrDhqPPUqaP2gNWFr4ZnPiG
SmaztKI6T74i7dD4+oXe7iyV40JwJmUSS3A8WT99G/HHEaTGFAQl1jCVFoGhHO11rLF+lUvf0z3P
hbM1BIONUAAycD7+eTb/2lyGnVoZbsGM7OgEthPa/ORsTVkTd7CIMOC+wkQSI4csBDx3XXKkE1Ec
f0O2x3y/p0iew5+B/t3EVy9Khs3CPcZXrYEEeOUUqUzINXbobFiEeT6AWlEVOpXggbPrzuMjI0UW
oF6loglcPWxD+l5pjXCdiIIed9okCeDUMDObQPAMqm2lt/eulJ2fy2hUuVu3bpH6dxM12a3aLPZR
WmsZvB8tbDmmttujJBYP/86f4ENPWO7W2rI9gBsptT11NJTyGWgkL3Jk+gV7rJ2s0ytQqYkhhiFb
iysoblw4/Sh4pNex+n5EX8ccgwKHViri9ISrj4pixKqAwAc/1t9TMB994cUK/WKfR7XUGJS51/yz
OsGCYOfRXEjqob2uzGM8HrkcIqZpRTrkhIPLQAesVzDBDWoRejGR0ZOHejAOduQSXN1sIT/k1Xod
XEtFVBQfZSX24+npCoq8s9dhEv3Jf0qI+SzWdHXlUFVzTHu32r4TLpjFnxsYX5Q7e/iR+BCy1e0A
8XeTfmtb30KC3xSRZs1SdxS38EJH9A6BfOyOpGHy7i33JQ+Al9qFFd4ekrIlCrstYASmCCAljir4
f02Fh82BX1AM/+bSCe182ysJ2F1ip/zkeCIXPs7go4NiewCclO5unXCv7+PoEv1K8x4QRWPiyuFW
YlYn6RRtXWNV8dChHr8qmrPsaQsjnZZDfH9ULLSwkKIPwPz4QkTFQvuIowJ3QOZDJqUL+V2FgYjn
z3PTTxgl+MsaFbwbnvzCLO2f2b0bvgGfZ9ILMBWpCTZFTcezg0i/gXM5Gq6Y47/yzN/odF0JWb8t
plgfeWJ9tTIXCzXMNCvvj3gWGGgaRW0qeEIb/dywocAXz672UqzdeewV1JEr2kTSBtSoSjf+wex5
dXtb5FHrYtoEHXwfSP2W6skAjX2CjoIZId9vNpOHeyHu4jRqIaTAZ6ajWy5a4dEzy5K8d7HHFWVz
i5G+DBn4ExfDEXLVVLbDOExwciTKyw84ws9pEZ3EJ5VFNeJgoA070sbP4FmacZbdIdqkAWc2Fnau
QEflfUHwIzUXMEjjvIRoKq2jJPIIBCaLPS4W886aoBOvBIAYVOjIXcQcvJNs4HK+sjypYDyDCojN
QUDO7vocdLBHoeWwqvRJq3baNoFMvD7a78nqGpGx3J6n0OuMCbUJ2omfytoSf8ca36u2WmNJtOhJ
/1ZSNQfq+J2Run08+2B0N8LSVeMF+9eSYjKl1I7pYrRSGUc64mtjD7gi7j3jlmokhRT/kwrMWM1e
KMs5P0H2ywUNL7WR7dVbNumBJC0tWCj+rcBlD8T67iro58VWlkXtqv5rvs8Cm3zmX6CxXPvOmIZ7
3HoaF3+5qyeji3ayxcFECXEJ3Vnvl4cniuYKsJ7zhbiS++xM1zSdTEc0Q3ctiOAoZVIBqSQh+vey
qoIYOjsYkgQSMMzV6ii1nwiRvJTYNfKBcjxnovily/Cg71ZdVIZoPdfSZp5d7ur8qvfLzx8ZlFka
RqhSFm7fpv5KGEkE5MvM1OmDx1ryQwvrJU8Qlem6GePJjLnE6ohujIatpXaW6WeAJxJ1X8c17uwx
tIN4+I/mYbiWO+HBK2DaMtnrE8DpbZLCfJkVpQIJQBGVmvJg4ZaHykyVOwsZiBF7+6Aj7dQDR8io
4U7dklG2qA1FR3Ize5v5QDxJkXnIsTsPxRpPfSIW5JvwK9Yx5vvsOMNEOfO6AUYChYPI6WeOQmsW
J9/7IhWgDmD0PUQ49uhZ8A0PMrGnScqwDkWMV3fEXPGPQMKeiNRCcZD4NLPpVEECVbw6rbkRVNRf
9FXVuF6LEciggvsHlzPxfztWLHsk1LuytNajZAfa/IcsaX6qtBvMahk4h+HhsVHvND6d/LCdXUew
+2yDgVO3HwKXQ+9ItdOCUuxhJv2MSQs+OdMLBP+R1vGGI9BmNTRfCpjoGsHVC5p2ssfLo4KumJbf
8ifOtzg73auDrD7R8y2DivDsXTX2BfWyZ4NKpRxcnvElIK43x4fFbm5I6MsC6tf8u/IHK6fWBwyX
ckwu7Dh1EwbL8F+DaiHcl1DUh7J9LMw+Q1suRwhn17GuIbmYP8GpjI9TeMIPSDiMIezMVLYeoDjH
WaTgc7YZSM8wOJN4XDduwpaqa5996PoYIWt/tsc37GjjQknGzaBtdQPzuos8sYWTY+0EPOuJImAk
s4+8ASvC4EqIJoTZIuJqAV84OXw64hzwgOgS3tjJlK2+INSwJqQ/4K7j25Q28diqXzP1a02vrtLo
QzhFjCthmJzrH6++VueTRmLy24NLnot4Q6Xg037ov7akG08YTVoi+x+EzhKyvlz66v00FgBrYrgK
Mqbfr6gl+2i4HRWY0RR+KXTeW7b1UDkV8xuBxfABOrFwfdSEnQrrPMUa3JTTK0BR0/EVnUBaKoQu
kT6MRWWhnwiYZHL3ShBwRl1wP7zUjmGUROLG8qf57ZgEWIXvGqA6jb2LaH0Idx1CRToClzTa5EwM
6cJ16Ak6wRGhanKUqF1h1fsr3PK5i3ngujPzwiVxkh8V33MgLtDD7NWm+VeeftuaHROZHTyDlArp
9Atf411OP/3AjA7Pwu9pubn1lmohCPGaZvEqkQMpl1xnI3G2rhkV9bloB3VgVpwDQtgW+2LsFTI+
DHKT2NrH8K7Cy/KcvWHjHXPL8T33HYNgR9nTiQmCOjP5ZVYc0qnLK6xlyskUatAgIlUgmNA3dbSC
X7sojTFzSbqFK92xyF7OEWtkXoCcKhQM3W00veRxLIM8HscyEtJm8thcRpk8wwpDLbSwdG6VTRVV
b2urLnubldpTV+sC//9T/Xov0NfpwjC9q2avUxRpdSKFgREgmVQBpjFjUKXMVhWyuub5J/BZD14F
OLEH4z22MYvzrrKsN99L0ftnKCKCMy2tJcjA0NZwGskR0LWlJTQw4ZjPpRKRZklK8+jS1U+i5HJB
PI8C5dkiXQxmQHenOFbdq8q0NXMkziTvB646762DYhSKkJ0kICer0u3pIMPhlqUNzKKiobY1XbEM
nAfKCbV4IxLADlGXG/197cTVzzLIhidrBG9gDJaayugNMOYS8EnlocMdbVj186wJwGIu9fl0v5Pe
GEWXyLeBVVghcIHzqjB7yXUnRMFDyG4r3r9E3qdVsVF8sfmAjs/CGsut8EnMDTQ6/K0arJv4qAos
vYESFJ/Ox6rDAMPIO2n8knRm9LGefRrInYljUvzPHbZAizCnxkW4sEkNKLPoslGXbHSzj97KI64D
SBOPFeUzo0zNENZ8hPuUPc/hlOuJTEgDK0MxE8EmZnFwHkvjtCCpSPaYDYLA1IwSbExx9guRtqmC
Auyq/88Dn8sRqxZwlEA2J1VF/zu2pWFzosZtCBQ+Bg/dNHPPGpeu4uDfrb741TdPzE28Fuk0pFMb
R1FPGTz35ZD0GDridVfis5hNNKIurdIZsint5rY3ADUf1aUsmC53K40ugX1YRwsQtZwP7L7BFsd8
YvDA/ctd/BRolu8IyCzu1/vpSSZfRAH14Ce+6oJ6Eg2hj2aZJ3V5VuFCtovC4L46u5QOekccB39t
JsMK3zeLQNZdUxAXFSrYPHnOd1VwXZE3JFu7kcuWaBZx715VNzRYxxmUNxVlZtozhqQeXKeuMNrf
+Mhqz2AQGFIhwbmnLgIZpyEunNdz5kqkTIyCbuLbX64rEvTbVekvMulNwwBVLg1HXlKTbInSNhBb
efKKCM8cURHOeGItKSzXZ0jpAU94bDWSyNb8snnCOIwsYTPeiGS2rX88HfNStP3M9E16ZmLD1vYI
JUsCk+c7+4DzsKluhRA60bz3GATftOv+nIQscYOwvvsZ6rrH7rbGV0pjbRNlle5EdnqeZtJxjbkQ
Srj9HUCTZDi+pz6HIqWJbIKhSbWA1HmLMSqSRes7WADhXloqe534ypVVS3WuTArze9I25e8xU69D
6XgXVAYimH3WRMe7SsQQduqzzPzg/Esw0sGoAnHqIUUhJlA6SJI931HP2TCcyHAi903qsLSTYG7S
35J0ecE+FrvaXkVW0pNDPbZ8x4L0wwseeypN6ZgXNuT1NoPrV4l1dIBtDben0n3jmaD2DbzRuNjj
XgKxcoAX5jySCcbb0FKXBTOl6FJmoh56++wbXeLJncXsy9XG9UR503+znKjj5m5ujSnQIkmNwXbn
BfSYf+/YDeNLVpCXqhTN4pOZVBcklqK58+FQoy8Z40IhqmsO1SpiwObSHnBWuFulvBySNZekadWw
QVe0qSzlLw1TpSlsSn4MHqjufdPe8Xd9hjDDvSjoD6dp/iOTpfsUYc4W/rugZr7wtsoxYaWklAau
KkLTgnYhL3X8qDC/rPcZ3HCp2FnHEFEdaeRWh/8qF8yh53Jw0dmV9Bq/7O82ZbvXpvD8E3P6OOdQ
nBZScxwvLvfwoRTeOIQbeCrJtrXJfN1JkA89zwpJwNbpHxmVFhagAwdJjsh2nE3vINc8I74taBzv
p07fezR1FzU9FlCYE73v3rrhaNMiiGm1kBBRmTtNa8Y3rpL5j1nFOmrMthO2GbiNN2gSIJj6aO57
4JpScBQM8DJi437Wcd4WRRhmxFVE9WLpQQUm0UInAT0Oit+rs3mquUMjjOBBrnzfameKMkXZ89uS
WupTwZQeZmA6vQSN5zaC83MKljyCsmTTVPcivRoajxtifhZJ3KNmyMI6kKpv6egrCn5nm+dqpKPx
LnqRn8tJSQbkFsuQYT96NI6Zrot4esJjwJ/f1PbnSQajB+0Tw9GfIJWCWlg/5usHZDhDrCazWT3y
FO0deV6wdeI70f3M5qgVMRvIW6P2JpBTjNgh26paT01YvxTEFccbf5xWay1eiBx0/ZxMJCx6nkZq
rNGmOYLMmAbW2jQcG6Zl8xBNWxHd6TbmgZmIrN4v1cXMUngSqzI5j4sp7ojuzDEfU+Wg/Phpq3KQ
yPBtyjKPqsuF/nytkF9pbhcLS330NYmCsCupFkA+YM3jRnis8PSCcY1UfAhnBRdtYrz1BAdc+NIm
csCy92TnftQXh6FSPmjlMuqg651DCUmzH/C4tavLg0HT5TXVH3cYq/N5e0KgTP6Ze7Jrfu9ZWecK
Co3z0zZFZ5I+ba7nwYPsepgdUzYm80d7SfMSHb9c8VX5huzTMWtdIFJyGSGc1j9wco1EkyeGVRqa
G4jfzqv2/zV8FjE+yNb6JQrdkFpCFWyUp/TucSL5jjtXZm0wySbCgRuXQGfezA6rnX5FCfWPJkad
vFcrOvtUvKULiQR/Ve4NLaj1eJc/HOtfSRHavKqUl13lUs6RxN36MILmvnoiq/sVYrGtaqL5xTkA
7pkORrvVeOWkLgGmlMQID7f4ikL1VX6qE467j+0NBgnayjpBUoszH4975V7HbrPy9p0Vt3S71Bzv
VkKNFXYL4y20yuhX0zO3MmKMeWoRuOAWsQA/IlLb30Rt6euot2/PMZeyiIq3/hxUtXQb9/DaYAXV
Etotlx48fWamU+ZJI6D9LuEp/awdaa4tL7Y255SzYs7eE68RPxoL6J25J1PoLrDxKoUHKgqoA2H1
85Ybr0XyNBQSx5PcF/VBhnveiBXEJCM6f65112sHKTYjv45DiZAnUeaPiV53QJWQE4z6WXdilnc5
6DMO1bTZ3V5bObuollKX8WXCtPBHw6Vdv9yIvxTD2KfRXdWL049XfCJ6qWVSs40RfRP9I5491r1s
4AQVoPHaW2H0Lg6wZrN6GlWQ/Jj9tgvqPy3D//7vHb8WYmU13gVfe1Q/QFb1yxuv6iTWgKMhQraQ
s8byoTVv9vDzHUidITFD7ej8rpNebkg1BAc4qvUGB7T/zFP9G4II0khW+ZrDdot5XAt363A04fmc
C7ary6HDVm5UsASPQ8fEkVoi8YT+R/WywfwdzzscS+O3SYGl5ftCYq4BJDbmVDCNWRQSIXLHJl8q
ulccbaFFohT6j/PUz8FNOX1KcBGVDEc7z3SiJw1BvGhs5aaM3viPrXQ8/N7powF8w66xoL9i7d9U
vwJBb8HAmIP16z7N2/qi3Rrl1rkgBd0ugcBOGxQivzlUePflh0z5ttTlPUYFkVIZaJKT8kbF9ACm
FRrb1Avas8VtzGk+olOOYs7674G7McaYM/MpNj9SsNvLKUX+kD1I3jrcMroguKdsaJmUgRFrJkSL
HbzSXts/WQblqygGhomb8+l4NrDXCWlyH0KqLI7dHADnTYzj0KbShHETMz/+ggZVcwYMx+A4Ahpm
/mzczX3QDhwKNJ8fC1keAwzsGHY9yyCl4+v03Z78Pl8OkxSjc0dEA4Ag7WTztmWDrKiK3C+kczfo
afMU9qo7qJmuYnkwFlYL4K0u3oFI7VOovjld9hmbFDPREE/pUFauAtLhwzGQJXJct37VycLCnr+L
BCfyJ1Y15qgPdic6ooF8BetcB2L9Bfuc82kLLQ4v30Dr/90s1xf0+OeCIcrzwVIGAbK2D7yquwz9
rjbkF+XyC0WhLndJsTdn9/04T+RqLWdB7QJCqtgGapEhEsL/la0y6oxkybtcrHCnrHeH8Osvg1Jx
x4imwr2ziUDxe5/0C1D4mQwiRes9LE2925RsofEuBO2C1weCDo59oU8MF2EdB77XnJYyKV3I7eP8
ej9z7o+845Epqkn2HsSLmTSYWNvhE7q5ArepbQAKFeNnR8n6gojQz8JS3dwTeZSFP6IPpplc3uEn
iwESBrq1Z1vc95GegBPDm6Nm9xtS/w3BONRojhCErDYZyYRQEAISIzYosIfYwABhHimqAx2maYay
D4r1Nvl2KIIKsbUBpRoQy7N0+rfsrIkZBbcl9qGiaP1OSE17XvN2QazgeJ8hVCL3p7J9Dbvf3iEG
JDfrKefpaL70FA+8gGMROtOfvbxyZlRc+sMDaLTqmNYCahovUuqHlfYAlsicSweXKP2tOz5T6Alo
oJLIKoHj9LKfCm0Y9e1BvJWSooubMR28+3brGOsnPepkj0ceDZGtm4Q6UUfO+fLQmRCUU5NEWMOJ
dXYVq2h9wHJth2im7JGZsPPm8omfcflCOh8HauDM5OQngK/geGw0vVauXzVaJLz/sEuzAgyagz8Y
3+Ui1dF7yfu6oPAR84VqqSOy8q0arcTz/6JnNGJ7MBrXxcjp0KdYOXmLGT2SHXJ5zJjIeN8gdSoW
BDMZxTy8XDEY59USvzHhYAk/VJxM8wy+nSM/vdGEDm7j2/QE/cjUjCEjuymEjGydAVyFUEPxs8iG
KI6zxwCI8iVAOodAh7lCv8dSfhVyrrr/TqOG7a+AsRKBxt+GHSDsLTwoWMOWN++e/8y2y5sXhu/O
9ah18ri7hdnOYomkWPudY2Wubfv8TxtS9pCUoujNEZqFoieLW7BdKCfx36ttdElkPIcBfzs9pCTp
5wRvbA4t04T3uOiRRNGNjA0tiTfgShoP8SFTAGETAgxsxCAVPYrIRrhaf/KG1n/oDnYhdC/dSL8W
d9bOlRiciHw3U8u+4rQscc0Y3Invb100AlJuzwOBsprsafEyjYY9SfVwBVpngX6xf8KpFa7l07dn
pYKmKF6BTAYywcnndmGOStftQwVbT88WzZRT6xD0ypM1d9YJGPvUk/VlFsLvk9mnJGkz+8PphxcK
swp9DwhSNdXAIiGP5exjOMd6QVaw9mkQuoEIeU21wEPispd64rdm6mJimpj2KxUNl+/UPc96sK0X
Jz6qxiyimjCCanQvogWCVBIm9fXS04uctZJfdoMOmg7MrlHSb6Qj9hNbgdNmpFK8WCc4rNuBimJr
qccFu1o4QWcOuVUf6JzuqtjJQlZoDoUSXGsnLIBg14Pt/BRsYJTMz2MVsxROp6euH/rU4tW/aTvZ
jFHLYEYSmV5lVZ5yISprty/V1dkB8PF0Y6tUkWLDwOY2VVdzVniAJEc49Vrl6ybfJTonu6OqDjKZ
5rF9qwpPeGMU6qo73/QAzYkJ5bSD9Ida9arU1tQrnxXCrJuUGaS7uxq4rqn5M+D9K2OXFl5JJaiL
rEXZ2NzaaIZEt6BVIfgfnKIY8gTjNnK4APpewYKDhlTu0rXINf81yi9wkdMexzLPDF3oz3ZCLwWx
w0UnxIYOHQCcjYbp+vRQAoqKTx0NbuYrFdRVnCLZFZ3Gf0NwBBbcj4VRJUwd1bktWJRTILST+Rs0
VgfTSlUojRtgqCN/UB6JuKV0zMgV+DgA4vm7JS8sx048bQnC0O/2xSQa/Fig5MpRwqFOWSjVHYYB
mIpV480LeYkdC4EhI7bF85FrfDOzqDmbO2eGpDks6iPJlyEh21wCYLnAm/RIAObt8NZdkqgz2CIV
U4gp2ZYo6hA5hd2Tgk9zvjdRhzSBENaMcMbTkGWDix8hsOjZt4K2xOHm5CQwFHnSislWJrB3Nz4X
4u1RC9VuQ4paLjw8tOhi8Uis2bqz+FY6KiPgibK2ZQ+3H7ceoiY1OeeGCxhZCawbSMtCsfaui9Uy
nPVa0AR/puEWwNEvsE0tdkMJ+KWXO5TKiD1tRaLTTcYrZhs6zLuW5q8982nR5UPkCCYwUHODzuyT
5T7nnz+e0s6x1aXX20PAkfxUuv0R4wrdONERBDBgnJ76GG4gz+DIzMmpjyLopXOOtLSyYhnp/91y
mN2bzuIjALK4XfbbGXgi7K00ep0eLazxzWuldsVnIWSqmJZYEgGgFb9xN+ORoB6YE7LbFAuBooAJ
qsiCALPPzkWWfpd8Q/397m3GJdmKMs81/Yx9+AztLnd2A4B/4kXtuxymwad6/vwwaLcZHLJGnRdT
E55aq1QLSehSxO88AzRmhQJhrgA2CTA0iPcqJ5s3kniNUWaaIu3Qmvn8olVUusZkm5APf/woKCCr
QkPsh3oVccK2x5kZznxOFkYIXcLmciS/Ga+PfEJLghklnl5nxJjNht0C0bno3jayyBy/n2UQrJ8M
uARpn+0eJjDwsgQI7ahzNFU4iiDhzqiMidHAKGPoXay7f2PatInZjpGM0mk2UAM4bIZVUx0gRAGQ
JVxt1W92yBEFV7BgMhKX9u1crMxFVzGbidH1eVvvks4a+spJFtfDpLmuc7L5iiYeo2k+q1/CnuRh
qrn22gfVFy0pH3V5MuKES1yRiWf/2XIWE49ENbh0Y8G51hT4Kkis8eO1v8wnwmIs7crYhe7sl8T2
aGU29R3dn/USaXTm/Y/6r0iWXOzZgYrQKk0G3Rn4sbAj4Ivfd9CHtGAvvjv7spkya8QC163d/Dl/
YiRaUnP3H9f3qAc67LDzgH7KrahBXjpUo0bJy2nhHGJZ6OHpBPRKzHHHkeN1ABTINZUj36DLnXdA
NZ5qUhaLkqzMgYKb+FI6xfBDnxIrnGrx5t3VdVZ9UdqdqXBxzLIpG+R/2OFlyvP0lw3Y2hh0+ipU
C5LNdi3/s7rAWgjDUigvOjORsfcBXBupNh2fj5HqPqw2AVPogxwL3DX4MGx5NKylVNwb4aPEs4eZ
J8tKZBaTuJzeV4eBmBlpmLHYkg/1Ax1M11Fn1NgnXB5wGu7G4zr35/7/dj0UAP1XzDB3QSwdj2eq
1ElT2k+rckLnl4dgK77fdytwf+bEkpgn5KMDdIJ8QpdDVuJ796V38C3xOb6t+ex525WeEVe4/iSL
I8ngsY5KFcx9MAiQ2lhBYKAUfq1ro4oaEXDvaNmQnCySi1cl22T8ZVJBanaqlSbQxK0AmQ41PnAL
WwtkCE8WF3WfIoI18FTA4OH+C8/xIhApaZ5J3eeDsHVAm615EheG4zg1Pgd2sdczD/wM5hBUV+vB
/Gn7tgfd8STPi1SBH4qOY0Pte9OKOVcBqdSeBJzHljGp2VrESymwZ9oheZaX/qJC81SGyidD+6qe
9lfD7Y5vEFcOYCjCZ2okXJqbIHJ0fy8O/6hXIUpA5DxzmtsAxFBKQHokZS68lj98YzVSlQornInk
tIHjdsyEerwnMk8K8OOMX1OTbE5uD7vgnhzutRHmytJkQ/RuZkU6r5fuE2djMJpKqOnt9acB3bYK
rdc39pgMp5gdCeDkTwXnkTy4lk3xDCULo7GeHhmtdR49bdROJMdvPq7/d1Hb2M8MSNTx7SsqKtbD
1vkAuxTeU4ARx8lQ6E5sM1XqizENwf2h2e3wgsiFaSS8edvpu6ziifZ3Hz0kANiluIFtxk6ZbylF
QOPh6P+dG+w0RVKh2oRYn8in6+AFbJVkm5uVzZxg85xhoJak2ZpLpWrsMeQZbY586Xecc+KlfVQh
BeSCZIYTTrqypFrUbpZVr9eBGwvuN7TLOYBTeikgmVyLpXe2LhT9rTSIB5h+8JaNamibO0+DXtsZ
fgj9iVUttnfjKd+gkE/akkeXEpdCCJp60jXMqZl7gCzSwv7I+QHVmZP6h8Xvx4Fos1gVcVvlLndQ
8fepgWJH1wdEj9b3Olz2qwzUUXaFNGnB3+k38wLVZn67Dit3Nvp6JhzOjDAnW0DZC4ftgISqLWSw
0dVkUdBvY6eUeLEjiAfbDT8NxMzlQnbMgcHNYuh2itPZP7UDfdDyAruqBo2IFKTF4rfeAFp5QuT9
1RRP1rH8jQMUP9ZSlVIk4A3+bFmstzBOL7XBC+ENgB81fc82+7dkkX1LpxK7PJo1iTYMTcxm5bo1
ZU9sI9xXMHBFmq85o8JGzMznvXLJLhLAb7rr1j5YEL4mIy2q/5YPXdUu3ixqI3i2ZVMa6u3E/EHs
r4ViACxz90STqmh0+GaWLjSIbmGTKsHfvQFoN562WJJ9hhcXlISQ55Z0fSR2+Ucj+KLcdy1pcWft
+Ej6eXjAHOU9lxIRutmVE6aou6CcD+gKnaAsqNV1QtZYHn18CGwGNugiOXBXlwgIlL3rFuDNmkLu
cG0LyxOcfoU2dYnkH6cwI22Ii8EzVlBJEYI4/770Sk3HN+DuuX0GflqXgVcprzooDknHo/DTSSVp
8iS1OvlJopyxFEZQstJ+YfhAxZzEbnnAflMc05Z/VK6riTxf2UIe4hVkrpo4JWQsUf9IRFBsEvy5
epnEGcDuEbp26AVZrRcoLBUXmS87bgiMypwUBbiPdPHu9TheecSED79mcPDvg4iCdtdtCxnlBg7p
TSc+nO2MOq/KD9g6BrgbUM5/XGZWcNgN6SOXC4irr0E3gNTJMqFvFP4n3qnnRgu9w2WacZ495eDG
bcDqXIlYGtqMNyj49+asHJ3Ne0QQ8oMGeheP1K/kp7DFveOQJJUJVaJkMDoT0WnRAMD3x/HI22Q2
9JYz8LvFM5BEzeIm9trlzhLWinMSWOS/vVk8PKd1iXYCxmTbWfc3+Ifd/gpj4C0T1+DjZcnmSm7M
QcO/pezTln+repXrUa+QCJLsXKTYizXEZ68nQeG0qZ/UK6+tZQjMHB6pDBsBXbFNLc3WT7yxkNpB
Rcdt9WZcFlv0UgHiNuxg/XExId55FiwC+pkqIBf0Uwn2lC20ZTZkp7X1tobT6IotsOhqVNGhmfWc
QbGcZDeMK281doMrdH2p4zqUnJE/rGuhjv8mqbNFUgATFdTlYoplqUiC3NUomFi7Z7lvQFKPhuLN
pcrrL7LLG8vVqq3J2Wfl65myJ2u95NSZzwgbifAk1r64xaIDDEuy9TgkIEThOBYX0nQnRZ1FTQ9D
sUxyXHza1/eHKnW9ng28wtaSCV9yCc0p0aPdwOGDDxb2w8/szI84Hc73rGphLO1RmBBt5/qKkqwl
tgl/suI3U2K0bpSd2wo5CEvgxwHlxUl65uCxAR1+62iktAsz2nWq4RMNvY93n6h5vfiI3bRMyDRr
4pDpvK+AoJ+PM0eSGTNkU0RxZKkgKjNigIefN+7iCp5jVacjbJKpwXbrlF+WccrA3G5hdn3JKxOS
v4dXr8YB7V4vxYcmkndDuMKwdk88rkjdN2DtM4ueOxD41DhbrpAPWjCDMj1pJLM63hYY8fvZwrjy
lV8+1PnmkNXcMdYcScK1RcFU+vOkjzypp0ECnBifPLb75biQHewXKgXkmNJfBkM4TKMFx4wBDMCK
SUtlh9J+9rYKPhI+9T5/Xk5nYqjgQkKsQosB8B5SLagWpyjPjud4Il7ia8aildWTSUXGGmb1EOyV
Vc0bPmJU7EHn82D7vtrlQ+yEfB2I4dhW8A/B4aQUqZpFr6ZpdHHRolEzmcqT1pT+C97Ie39pQmkN
sJ+tsE48BnXX4oFf7RaG4agoEgNJ8LBcwYm6kF3Q8j6+EZzpSorEXpUGtYpmpyTVg3PbLro1uh3T
v6zZ0JD8SZMgZItNpun0wRc9zD9YjFTonAVnBpZsUVUdhQSwNdDYwETKEnw4NLNqejbjDLeFXwJW
T2+V+PS+rIamzALXNCScr5M/1lLP0yWzXxmcZeZszrIwYiz0o6JXjhw2+oo4pLf2ucKNK/JDxK9g
n3+09xHruZfMCv2ROw63u6JSZ0bNVmnl/BK51tC+AjjTUz++9YNZ0ynhkfQkAUdVh6rvOEQ1kqlN
axwA8VNYD1dg9haxBa1GU/23ditBcg54RjCwU28iMt4QbNxwDGe9aj65uDhOOmo8Abwv8wse7kBF
EfcLGrZU2NwRbZQqGPu9WUV2f0z/PNXOzfBcksNYiPtLJb4JJ6LGPe/h+fKvf45HzFhfojKGjP1n
CuxkHzvwjT8iRUtGpvyHf3hce+ycKLYoQprvc5VGJbprt1bxC2AOw9Sdatmp4UDQ7ZTDJkgSoxTJ
bh+g3AyWyHTE+bSujJDvOd0L1TxKa0DDEcQE/FWcYmZbkwaJBQRF/ib36SQ5RG4cM74FYv3Ut70N
pgsLzjOoz6EUwV47p9vtcuenIpRZyMDbTKUmSiJR52TDGk8MJhuRLhl9S2aqRcLcHEP/FH9s2y9r
+OUgV3hFMLCbUN/Vp3RR6730tMObxRSaCm/g4D+vBZq30H9jD8/D3yuXEKDA8j9046Xq/ReFWtn1
Sx0kIYQa34t9Mpk2KCXEzHlMNM0WnX5yCngbPa24h6erMVyj4Znprg2TtLqUXBGXK1/Vv/Ki24Mf
rnfInJDX7haz//S2u7kcAuQs2AjmzN7FNrp8qbN+38pVq1MZtKR1F48X5yrp0woFPge+uQWCAjpx
PujTWC13+4bDzVcrzmdGo/Bv84YXp3NzLVE8D//E5pDvgtEZOaVbw9l6Zq1gi+08/1nE5/ATiPiu
I/6BdExvU26BLyi/MlXS4FKIF1sIX2qLEk7iq8AuLs6XFg6EaieHxdd8zunKWidp4jHIzWY9JOAg
lTgC0VAsXflOwcNBOgS6rY8FnBYjvr1olVy6wT4nHNfSMF0tOltke2Qhi0+tLTlfr4TgqPje/hFV
0U08sZjH7Qg9/4FFbeZci/IT0UG8k7A8QlDKobm8VQO2wQu/8wWn4NbRi9Lqd1xrlbWpgTHywjrL
eLnfeHWGh2CizTZvih+xOC/9SyIyORU1xeP3WJDCU8IeERZvgkU90QawNIGcYNb0BBzecVwA23ar
c3fXt5PoqtzV7i9mkIcS8gv46h4KRd41+sUOAFTsasQJmkIbm+tGUazu4ZgOSDX1Ux9FVYlae1Pp
WjHA40yf13ZD6JMaKXkPockfgTUPd7aIYWXgKLbOJRTpbzrszMub+3ufGLx0+ztrl0xVi5uqjvFv
WHxCSyqlawZjtoPyw0GkxRpMRmjlkI++nVXUk23jzN0zz4hZIHRmxYACh2j9qywyraoHzRQBkiVS
vbUyuVw+pZ47hZ5UA2doSYi/8slG/n2PZSbbc7z17SkjrJuupjCyHfisJSzfzbQhj/DwA0ufJAqw
IristdrEoL9fS1tQLmFAMNknusygLDn9TJ80OJCzag+sZi4eGQy7bic32yjNeuEPAbMNxbVr0NZi
fCdYPYVNf5u6wIfb5sOW8Jl9kezaB4ZS4KDPRFRDkvCSiCqkt5UN4IRhvhN06qVNGs8mkWzYVdV+
lXx8bqEV83H8T+qPrQxhnu9Fx+DkjNYH+WtadjUQiaYef6u7+r2FJUF2kJHTwYnutVBSJG/NJLS+
4qZCVxXoFbl/C9v1tWUU8/livJ1gY6p3B3yaZHbct8H5bN1zwzp+83wn6subupwCU0pgvM6ZisdQ
KhHHKG69C4SZITv03/XuVNJU8h5VzNN0oDeS1UTi0aiV9G4Pj30EXjqJ9qcdMayiGqsS/YvVu/2y
hLf9b+lZ+sejfdwzT2AVt33Lrhc4K0sVgOfbE/mbu015DFG7kw+SqhIQsDdBo3acr+KziHl6KtOp
FgCib6Noa42+6VlNEgigERQX479WNwDN5BeB1mEsimOiew6rtwoc1KCwPheplxOBd7uJcbvAbXIS
S8knpbaVAXuZ4irL/orPTy5U1D/Nn2tjxHACFOMDFE/K27VtR7tszGcMxQ1RherMSovxzg75wLNX
PH6r04LLMJSfUTEkVjaS0sOjul3qpKXxfAdLGP+b0pb6uKJ4URzPL9jMXNQmOIt6/jjneYCqE89m
GVK0taKYILmrJVwzzL5cJYTN7Ym1QKImptvOpCN1LRPGkNgqGELlZYnmJt8n/VaAWHZd2X7ldp+9
q4nt9os9bCdpZLSVMKxtXVgyEubQKuJih32q6bVwzF10T0XoLYLK+9GScTU7gQshVC1HKWLsPIae
xH3Kn2TzXj3GruCCGq6tNRtxGpl+7gJBzQSuSb/UoteROL6xa+P0qw0es2G9kbKeIc3Hi6SJ4Cai
Uc5WKnoWQ1DOVjjhYd5S4Uh0I3D9Av1/HMA/DVtoHv0xwga3sIkhIOiZIQ2dPSUnOQmNzYI39r53
lgRIbJgIuKkd6P9Aa4f1jO99dEC3kWyOHvlXTq9/nkTqxxHBcc1uvTeZ+KLl+FbxVL8+tGLf4Jan
zec/gmW3G4IhoFua/TpCAQSDv8c8KKttLnpYmV/0qN92JKUUfY/ZAgUhFl1RnAV5Dnd4vfi/ru0i
Ef2Ph2Vppa5EpArL5D0GIAFd/ogtEn1D47Q5IbLJM3IEQ3cSP3Zp6fE/zwQ5a+XMNOPgGBCKspG1
hYb6Ax4K5l0NZLlrpuzMrXHoozEqNT6hxiOZ+2sJ0IF/DrTVTacRWqcfdt7sdPYk9u5cyALEM05b
XGLY4BoTann3EznCslMGBqawvfE2jrBLN9bqgyS7hvG189HJ5v/fXSwKjGmDftMcimIMUEFrKSl/
ypmYJnVf7s4ZzSBtlhgcT2zPBkzOL1mgF/Lt4NVNFfhHn8GbLEwQYBkCAxZFFhjB7y/YwfsczPWD
4NfyPbuemgMLP+yjSTv4fG8fBH2zQmrwjD3yT+9aAsFS8aPUzmGiJ2knz6Hpw88+8M6vgViFrjqf
qbPFBz0W9+VHJpRavSnra/qfEuJdEK3wK1dqApws28lbGgDS1qVgfjpbYCbEN9rSUKWnzHEncE2Q
40k1ClEl2DUF609tPF9kMH2A7BqX7Rn2lEQExHMeY0xZXqxXzdvGLq+AlYLjXJwoGZ5RPlnoG2CB
2DLx3YYTBSA7m2qjtt9DvTSPa36/RAS9+GBNS9/I/PCkJzZkujo62lWIdy4FWHl6dXGsA3X/Hbad
Ixpkuh9VXgnPNVWEzL/fxcdT1bIfUhr/JMSVHxWQqO++M+tlIvnSY4mgAx5Bqi/TBmI1M6Tmcfa+
CegWQ/cUaw+kR+Z+cShth9Qx00SZMZcB7TGmyqPxG60pl3c1NwrBQ+5eyImu8yZO7YxiE34G1dD2
I+LccQU5S4WPbVPf6BWlHqyIrmt1L7AkEfkZeBPQE/aket8I4agXpxZlwiDJGYiBHccEDOL/Ysyi
Pd8XmHD+owBWryNVv/psPRp4JRTn6nNI6zOZPUDRvoCZjvmVR26yhI118fm2B3uNL0TTYg3JzHjY
Ur5/a654C1xiTiqo1DAcHaLbsiYgAPBQZnsqgqZWufS6fCvxeFZ6I8XAE0Madpgf5Nz24gPLMHcN
mLZp8TuhZEebuPNdedhUfhiHH5y9sIaIMR+gdsBOCIJ7rYNfxY4kfBHkl35SM8pSFCL2QzMGbid4
UIa4snslP0HKU34zSPihWk15fn+ekWe0HBUweXCeBxAo2V4Q0zgMA7p43pZqjvAH+zYt6IMIWIbS
aXz4YA624ZO0PADNFhoNnhPfKBnCjCcx8GXQuXPU9plAkoZWOeALjHg4J7JVm1CsQP7SBXyL0jtx
3Qb8qNUBVTkkrhNJKHbEgkZ21K0KZCcXhxqs07a9DpcJpamF64htpY9PpYcOSEahSCrC2+x8l4DA
Iqjj5sLYx1DZU6M4UUrkRtIe9TeSqJMNEnl6HcoGTGx8rv/ByJoA2YwM6Yk178hh3w1s0mZhwYvb
XGmjfxNcGReCUE2tCUhmGMaQRHLzo7VeNmPQE88BGSK1pTPnuWJRsAcSoKt6Ny0Z6Bqih/F24oBM
U+yEM7noGa7Gi9XiBwdQ+a/N6X0Ck+ZNNlbUc/Cp4f7w8o0e+dpdvC5BLCJPqBFlyTBRwM0crt1D
6WI8rtN3JC6a/o8OJbpvJmZ5dPWOj2Wyr9ty2/8RTyB9CpfqlKYrD4uYgL4kQZGz2p54BsxR0vJS
Fm75uzuwKaO59bhbSkVK08bJ/Nnz97DnFP3dTPK4XNNoZJFqDHVpPDehAe5eHaXDUoDUwvVpj15G
yM0QDfH924PVn6o4qlOJpYLAH1aiTI1D3bbPjd0JAg8FGVc5j2ahGZ6LgO8G+zxnJaLRkn/TQjm0
7FgcWo4873Q/Li+Eld1oDjd1wfnkwSLxcXGbi+JlNXtP8WQSJJibAlMPFyZ783uIQo+NicEoR1VF
cgVFAgBmBFDgnTrjTrWTRySbTGkzQ+j/iF2CdkbyWNIlnMzNY7FazvuFvVMEBr/vDHPSsyjck21x
Naey4OOnRt5ZCWjiGJo0LFXsufn7d5un6OtLxE4GAsqY7KMNTIcFE8dDGbjTDuydEHStmypxSElB
Mdz2+xJP1DD8hxz3gN8zAttblfnE4QDEag6Cn6CJ48rhFWGZB9vtBb37fWddSQYAdGshg59TRyLr
edvT2mf4v7SUpIHBMRB0HI2URTDWomQM83paJK31bCAbx3HoX/lW0cFCog00vPZc41I5MdcrvHGu
bx6FslmdICgs07S47vdtoooYDmBxSxen76SN8eTjsPXkoYLAY+bz1ZC64eHWv/MW+DDYj7WUuOv3
f8zfx9lo5uv80KyJOMdQ7oB1iUTQfpjKVJD7dmuc3/yQPF8s5OZLVrA6EP3WnxdOHzpG4KaRSt/Y
w2FGTBBwYNc5MVt7f0B3SyT/JQBeFArCmu1pLR7NvrdHf+c2DkUbX40WPD2sTKNPaR6o6F9MveT5
3ikle4HeA2oj7UaRNBaeYjP8FWzscVEoy7io7mmvqv21MyozH/OWEFnUnZwWNyAoPihhpuWbPTAG
ACoapK9GCBz0CV2xRpN7ZX5bv61jI7PbN9qKH9mtp5Xoa4W6eMf15pLgMHE2Pg74C6H3sU/CWK0K
ALo3q9w63qa+oRDJXzHI5br+OsEd4/29b+vLjWfDx5peL9tu+d0J/ahZgNcVcaZJ5QvH2ndQbN2q
yZIEV0HXY9scPwaPDEYETAOKkeHCk7nUe4CAaw7QRvb8Xvd/EfF7OfFZV5ti7eSdCDQCPTNrAUKN
RLWzLO2uo0GeNobH9+6QJ4uEQajgeqlJapqlmSoP+8PkA4Az4RVn13oCIH3BCT5jXkByrXzg6Fkw
8SnIlcaj4OBuplihEzmaxWe4IYcQkzsK/YCxfCZEJ3XFdLSVjoXt4VEjy35NvoxiDHSmZbSxe9jS
EuIYMAZ9qpYJO7gQyR4Yr5cWI3tRdReBmKEn0SkSKgfCstwEfP+AaKOzQvhgveFT9XlcDSA2aZ/D
stzGceu2G5mNNv7h1cUMbyu2ClqgZN6qsVLQSt+I1Sq2YxRS2KDgvrSL3EFRjUPIsMJ4EL3M069O
a19zZ95TE484/A/zcGa1aro1Ieag2SMtNlbdw0CCuJHD4S1GH8TqP6qWO6fZ63fEUfWzUsSkt79n
U56DVeeu4uexZenfnvpZFaE/Obdln9V4fnPZJ15AzRNxchx284vxUfyINV9w3KHjKEoRw1yYfv6J
RMilVlAvW+m+7lXe1qu7JVJRYwW4bE/c6LyqmgFT/mpAy994CRmKPWZqMvRbUonrL5424ySsf73t
A1TrZB4wcMM2KcG1Na72t8fpO0TbuTgcOL07hBnPV/xPgWGRk59rrWfgEz3nm5H2rX/rPNPUKfKE
SUywXcmzn3dclphW80ceFqxVuZaEmS4b6ITgkgI7cS+4aNJA/Eiy0UQwpAo9PG3oZDlcVTz0cJx5
t8nmbPXdLWxW6ZPwufm7Ys9gvms8qQ7Ar+XuJXlxZkMEh0B0ceHRNCZg2zPg4zls648Ooi/zJrow
hkxQq6Cd8UruH71Uep0MtA6+iePIx6H0n5UYbvJYtcmiHRTP9VFq3JP+EQQS3jH/xqo7DNo+81Of
Z1wxknV9CmXQ8AY63ZE6x1FAF55nvRjfEEBd4SrSprnBDwU4+FWxb0g33FNMwQ0F7G1RCFNI4Sz9
+qVrJOC3r0LXjYCJvn9H0MhyYD7ry+W1zIh9s7A6jC0uWdKKcKXvN1LWFlIsodHyb3TYggmaX5ZS
m94MighjjgGa4yXE02bgw1P80DwEA0WIZGUXaFIIH877RVR55K1Kj/bWu36HiOiq4ajT5dZavljr
mf3/Mw64MoA4mFKWa4gOih0PgwMyZkGY589g1ce4IWXevVxFt0tXYvHFX8Qqc22zAyc6Du08HKRk
PpByN1FGiigT+CZ9/BAoGGAu9w+djt5BO7JVjjeDm6aDE65kk+ZYlALXiRn434Npj5BMHubKWWvu
ktYT9eoc+Aw9li3JJ22Q0sN/mrLufjay4pTj8/fHyzbq31elQ67M9YujS9sNq4juKJhZlTsG7wsI
5aJ06mHxeuwIVVQcNjozqwPp+U7Jz8uVE02AfZzqwG3Bks8JkBYfayH6dzeqYvpPkJnWNSTn6xok
5rFAzmju0+EbkrnR5lRslFQ4RJLOrVWY3dNrGDp8/Etnka74iCskZv19kYqvfeb7IX83kyudEsUi
PXBxdcgQ/AmmUOKBL91+a83KsBdn3m2Qv+x42Ib8sNMKHhCxq9nbqx7u02JXHr3dOdZOYe0rKmbd
RpqNRmZwvIQWnuN2nD8Rn7Fs0DleDSB0QlwDWaHd6rbVpSeV2tb+eeumXbBGLyeMCAaRGb1BGaVe
qA7o9mcSNCvBOPH2H27VaVgukcyntXvNwwYnaONsevr/m8zRfFY3LyYRAO2uWXybQx0Vbs7dgbgS
ihXfIbW+9pYuwh4WELPEkCsP29FOd36je9SCXxEYxuBAx15fiHtCcJW0/qcMbEE8dH46/nlkeeW+
/ScCHKA3L4MmY4wfHSCY1RSGe83/Gc3HyCHJ84uxHqCIwRVOg6xL80dlzOGS6Wl+7Vth8TFBIeWI
sjLPrMbqniNapJbCKXHZ8M3HleiGhBOSP5QEGmP6o5WEOifiOJd7rSN2qOvJmp9+4S0GgUrLH01L
zGStlCSKzMiga8juGCxiZEquk9e+OOszQse3CJASaRDI9ZiQHoDAwhK5vduPzB23GH48wUyIHEci
ouM3Sc5QPbX/r1EmZ3ZKjbYl9E2cs6tOYwX7X5dKZbfdBwjf6JJ9LpSuQPwqF289mLe9sCCOuM1E
UWZga89rffzzR/j63NaHeI7kl22pNBLEujteiopoONNf5iUZZd7XZiy/zbtzFSlE8fPiGry+MUhE
nKvR1GQoRb0NYH7yxe/D/au/ozsHi4fI1zX0JokJYYXyjrioHgh1HI3srYWkVs6S+BtsbtKF95BE
3Fl+fXIOAStcrvDXRD+JRwNAzJKGqPiyu4RgkXeKZBDdcqblN3FDZXF1DgDL27XWcEpInanpf66g
huS6ASj4+YkecjYA6ibQPoo1rRFIr+EU6xo8M2i6wXLaerMmjgZbqXNVO/z+ueuOQ9RvQFQ8wsIl
cDK/tm8XwkL6SG7a6OUUJ1480UpgsMXYI2o35K95ESJ+kXaRajoD8xZG0zojSD+zvxU4LitCGH+f
4htWUpWgsb2SMbO+78Cdm+o/jFNp71QEQW46BJZtdzjsXiih34TU7DxHdC95QKTwJqWu50ThXGf5
OYpxlJF7oQPRFPj0on2QyLvyWn/cihtiLM4rir6j9seYM8VWAnFsMTSAerzoFbm7v/79hRrDO6Gr
byyzELsVmyieu/90h3n7rJbi9sotP1wMu/FOBX1khHFkW1ZIQuUwA1jkXbyaVImYJ8kJdsYn7Q6p
rgIljkUGrKu+Nvw/MzKybV0CJuEeXkkkNZiFUrgM/xHMcXlWGrGFXN5WMXAeqCF7Ux/f/u7MlxAP
TTSzB5i1CZPDzQ+7Wk/90gwM/MQB1NS6Q4XFQYJ5dUBJfjDGi6jzGNT3ZlZZhZRkMUrJ8k/UF6bb
iI4c1WpZhapz8ds3krNUuWjymh0Kod4gJ57o2Ln2QzVBfqINI8NDsTxI1vKz0j8IjbPev+W4yHYD
NYexyKseS4+ERFLW7rTz471jk7fDYhDT4PWyVpV4NrMmfNjhCIylMVfwcttsN2Z+FkYux2BAXqmJ
LcRbVgHNzMV+KRNEE2dI2a+djq4wqMFqPCK099bzI7wTVq+D3DCk7p9N+1u4e0Fj+25/YfOUdF+b
G2MgPLHc3MQlvrcmbGrdsOE69I77Hu2Qyj9cCOJDCGTzKsDgzKQ9Kc3S/VsQVcwaIoMsyuMdy3Pl
yuNGK1umusgAjn+byM9/ure6M9sH40d5WWrRJGuDlbeq4IOYqzthA80M6Hr9xBjqJYwuU4w00sRT
niLcitK+g4ItwTGdupWcHfh50hKfH365lvd3HFob9XzQyBhRXprcBbXC6E4FFgB1XrMbeBPkeE5G
my+qx8l/Adchc14FJ4fYFVwF/jdpZRSuk8LKUIng4kYo2D+BVJtOg2wHXq5HE7c+iUUvZ0OS5xYT
o8J7ti845lU1Vjx8N0iTZS056X2H3cf/2Whr95ZGFeHLsCijAhGn0ew3OPEWhwWvhe0v7ZXnHnVB
BdVGl5Qqc2ywnG/tQkrHVlLlbyySLnS4XKta/RixSjJYoYO6SlVbbD8sTjvcKd6MFqnLvEk2mbKz
vl64+S2RbI4MEA8663wBFAeN1vWh1gE/dG/4iwBQvuQ56LCe4qfkgtvWro3zshoTo6CpaTZ4UGpE
qpAsvvQ9Kb0VCzbDmqw3W5qe1j+oVKrfQuL+5gKQYZc4dbUWtIpH/76mx+HYT35TSWAitLLVQkzG
Ns4wkqCb7Uuvw/7dfPFLNyK3shjQE2Qg5ERsPoezkvNgKCxZjsHXEDBItIqy5m73GS5KODgvg3ZL
owYvwMKpxeE06n9CeBAhNeEUKrStJa7ciP9mtsQy2R0Pdpe5ObGNd+MOVHSttvUf/OT95uh+VQS5
RYG7TNA622Ac3zCUHD7OGAaMsAF8bxYpSMLUPGnjhp5mEPZNI7Jq8qTJj37kqngYkeF3uC5cH2OY
k1DJZsOscdw4A+tWQZc145pDLgHFMq2ehWDz5YCc9SI4cV2ofiqyqQ5zwUfWyiSOFRR7WHYxJavW
U0fkqACZH4mVTJh5Zusq7YTeaKAdsin6l7+OTn4ANKThzIAtdErU9ehBOqAOAa+RA6S9rjYhyeBM
WMlq+I0K792PQ7JYRIcTN+WvxU+JuCg3b5eCPVpXJ70a+LX1gQSr/++9fkqt3pFuc/mzbqErSOqN
/HvR5k5qxWuB0FT3AByfZk0EiuYbSWDbCGG/RkjV9Ci/ROUvIgWwpoKjaGU56zRjv+4fB1JvYAWo
NMWET4ZRa5qbqPFmOemiSu9xoggZ/HoJDudXoKahXwmMDgE9iUN6FBpfpe9cvjQNuElqBHLjx/h6
x0wA169sizPrCztq36mpPJTNuh9/2ba1hcD9fqLJHhG7yYExDl7/ft64CGrTAKtPGdJDjANYU8T7
WusRo6Sva8sbY8nOdKJyOwSTIjacuF8cnl7wQbO4SJ2AJQbkwm1XXoS5bJYguk+hEEOmXcPo7Cwc
SofSuCiqSaLYAY5tXvfEfSuv2GlorkXvQ5mSJqbuEjZsEBOVebFa35DEzQZDyxh0hrA70d6oI2cf
4nG/AFmJOkS34xApHokzVp9junQfyUfTqvfFafu2f6V0RcGrHGeyxvFbV3PdT1AKFi0GJS8nkmsW
EcO6e9fMYhVRg5k6UoxDdgUYuszKZYHIkqKeN5+OELCtTMPHkXe8puzf0SnerM8tKdnturuCcIm8
nzHZ1F3jBKFOihXZZeMF09J7jld6KYvCfHdSGJPkR/BzhiZfT3lq+z/gTafrNzW89JaMUs6K9BEf
Li7QbPPjFHgVxJufJtYEjeQh5NlTQheL9Z6jDuiE0wtzM7POXqeXQiSX3c0UHgR9E/1JYPVQjGew
eT17iA1ux7cuLk6lClO0AtD2BSXXlcgakRZp6GcW2xI0Y2KvOTJ+kzwaPEWJeQMpWvG9jS7O6JFb
oDQznP2PxwFTzdWkTi/8I5oZ8Wsgy8oeJfp7F8RCRdhhEclqdHcN6QQV/bpYpGQ71Z4YvLYXcXr/
0TL/fhaJC/fATNpO84e9Muq+D7Qj7w8iE69F1U++hU5jaHOMrpGjD+i4R9q06VfW85BM9nxk92N+
bD66tIb/s9EWobqCfeHJ0/enGBT43T3xuOXOgzbsH4oqQcMAX81bYjfzUhrJ0Bn4Qg0E+UF8oR9W
+4sdc99K4ndjzTeNJo4VZTz1Fv/tUG1IUZOaVuBYC0wLCviYIuRkNGYbKsPe1nRl5yKGQ6PDcB03
9NL4qAd+x7HsXwcPIfb68BinPp0Ff4GXUaTz9j70xH/RZ3IGgaAAORmHKtKEIzj5bUQNuZiCs/Z8
1dWG5GVsBFLtVX+s0gbORBJoDDJjEUS5gUbaKLKZ5EwyJvmzqpv3tkvZYZlXZ3fjg5pO2EUEmK2d
uDR7wwhuD3Ntlzh8psIzCZF81muG2W/QBh5Ss/5LQv7sWHCMjeXjU68nBfvXTlL0gQnbh6jyC2HI
ylQFXoU4Lyw7fQ22fRJgx+vLwr8MNscMw4BFcdITRqzIVYiRVdCK9g0Z6bfDo1bKzMvsl5DSVpHG
oYL24AoL5qwfJ4ShRYnmdvX/LmSgg1D+XQ/UA37PWf3rqTyQcr7OeM2+lnfhbKGxqc5KzGJrxHl/
A0agfO+YqOjyVzp/qTGkO++5Vtj/Qokv98P21DZP+hqWoSx/yIuZg6JJhfQ6I2XE12ys6JSEHog6
w1sgeIysUCrMy5rFCW2yY86pdgOLHO1bBT0V66x/YJdal4ySg5KOcxpqpDCmQDVgRmHVcALAO+UI
ioWarEPz4jrEarlMRZU1IdK6IW86d+YxrTPWy+AEI1+mgHA3OWtQiaW0s1T/ovqTT4uIWPSP7M8k
OBvWxmCOWBKuE3JbQKPOZ/gK9kEiB1zHlQIGEZfHle0qSuohQiWExgj3FV2Wfc0p5nlKb27kx6jn
0w33BmA5X00qKFXy3d9Vz1KdccHsl+2WoU45EE5Gtk0A+Z4tcxUJ0hvMJxLs+H7xuFMGsvBppU+h
WIi07+3Zjx2V4qlWaOi+GAe8U1RqgrYRzGbAXsWpWC00QWYqY65TE1gjLdkubw9urHLtATpUF5zW
wwgdbwtDbrfo6+3USG22Gt4hUNnWOTJloU6h2s12bBioMJ1Uf3TYfyhMYUdR2hZPQKtKaNcJxUXj
4LQEOG3NvbBiTECcTdL3n6b3c+PEEpVehPvTE9gw1HLdRRvl6pO42qEWpUHhvu6fqE8/tknWX/k/
IJyieH5cznbrA6szWK7Pc+oGbAwMEkYQHj8RYrUFasy1ifgnBin1rCO8feYP6Rw0uHReisSQEAgW
wvRmiFYltYeGjnGFsVjxcwIF1yjur5YFd9Spxj/q6iIeaDQM+gm97CF7q+xmsDq+bsrCORi3gqSg
pu+dvD/Q7Gq8ROMeDoU6F123m7cYL9m71cjFctoBt+NBrIj0ddF2X0CeeypK5nU1ZQ24ljhJlJ+H
U1PXXXN68h2GdeAkOyu/1kHbqAHqXYcvhzA1AWEcIdQUwQk0QDW3goHQpkLtoRHrqgikSmlBUi1Z
dotGERx/ND/d0m/efe4UeEY95ch0hebOZzAMijR0U4+SFNGO8aOtyP94OxFuiWl+IaasnUoN2X5A
33b4taZJrjlpdQ13K1nXzMrAVfXoBaQIkLwM07QgJv6prtm2W+bZqWwmgqOItBS7M3olcyYFHnYj
ciuCivQNbjsiUqx7mTWmeRfYfWdOLNpGO3a8Ztu9xqMAJhhNbowFi5+5BWUJBbFeg+M9aYWgWB3W
dkToUJorSPmfzbHslNZngOeMoHhCn3+tpVbggtJYtvvxTdQWv9KV4BO5I5yqlumwWEIlxuY58mx0
U3MPMHe3yJUivJ+k1VtcxZn1MO/bSqlYiG7OUsbDTJ+Nllj2/nIhVBEGgHLv5ALnx2XakyLXu7JS
S2SJvN0VpdFAJOpFiuylDgsIuo4bpRsfw2biZEgDcr7/Hg6+xrPpleG+PN93h+KuP0j7boDBhpqa
82h+VZlYG+/I/HSwb5+LAvVvJ6Oz4Zx1LY6MsJB3k2HvjUBL14d9GnjAyhMN0FGryrIRdNmQisP2
VduPLnLgBNiMrmkz5HRgX6/WT6UOZ6XZIixq/UKFDQ+S9sTh6filz4btmx7fv8/+Q/on1QEmwAAq
FhwGtcA+ykliDLF3x7Se5esMsVgklJCJzXTZcnFSh1FMOwETTMTmmrk5mhl1XWKno/mQJF7dVrQx
PzVV93iuoR9MX1RL7tqvYLcUjPiR1sq0xF00vqMdrvJyXFHzHCc9z7QrTV2a+QynMj3P5Sz3R35I
1SE3S9PHT9kARJMfCYPdrtl9THKTIdyN0N3GjPV6CUifn3SG4ZhAvwLy2vJKIj4a9q6qOgcpZx9V
2VgzJ3/Q/o8HxhcNW8sou87gkQF9j09hmhvDLDg1ShY7az1r/el2NAv+nf4o+V6FeqyWPHxGSwz/
q5Y29UDedyQcpEYqy71hSoAd+6JOHrwEH7bTNtW44MKxah0G8PffHA1ick+rT6HKGLIZbc5pfdNP
hsP6lJguczWN+nFl0oEKLlnFZd6vprF+TPp00GlKl9SOrBiEIF8ApOlK+bZssPrgZZXw6Ne99XPc
CPm9s5eo+d82XAEBa2BZOyoxsxEYBLlVY4hXl/Hx4dZ1qrz7LwKcRiqEnWySjMvuQXlCF5A0ReiW
GV5zE2l2NivL/2qJiUUuQXjHg7GTuLhy5jpRti9VkiEydTITagTo1mCtB9Yph/qOE2dcIIE4z0Wb
osL4HTzPQgTTuQS3FPsF3xlEZuAsoC8H9IOdDmstOLICtJrsZiM5AZJ+o19fgZC8xxRXKrmamWxO
JMB4Hg4aAJ5/N80ygOcjr/bbxOrMuczOYOFhIljazK7WxcF4xyqUOzB2eqpLhbia/3hjVnqttZCH
hfFpXakQxh7doArKe6/hdj+vv99s/8c6qUZ6mQG+NrOzOU58dw5aUZebKiMNsto4gJVolEWjl6lO
Ua4j867mXyjcampKRG/b/5v1INoakTm12azzI99lXH7Pi1x5w8sZ9ifwzZBVG7yVyHWGkXR52RfA
Z7DtYH7Z4KLXNLl9hHI4aTjP4+2GJOmevyJn+FE6N+g6wUhsr0haZ4LEJ7CtfAjCJjcn/Xyd5OZQ
YqgpTL27WfAKLiaX1oJp3IwQiK4Vjt4uD63egduDhlGwyZ4wle0LvtMNpkxjdsywLepyFPif5NQi
uyx5Q2G/H3lQYszATx0YTZTCwJJPlOHdK3x5JrGehRr7CeyqsVXBktAHmBWa5A9Sfoho6NZ2Wx1G
TRrvwCfnk/Vh3vvA6rymAQS5/sk1jQhBR3bVihgdAEn5pbfHkzF044MgC/FyJ2hlOakWR+qo5JUE
VQLnFseQNsL3eFuWQEF6vkVeTTgngCzdSQKZE25WSHJQXxzxlv70t6ZHTotntIQJytp++9GeuWGf
1bATJGGzvQdybwESUGUdhSVRsvlXI+MdQSMfpzvN4MQ0A9ttad9fmk4GJxto9K/jlennB8kbPgoR
iBdRg8lpVYxoBMffwx6ZGJztJAwK/AYYzY6wX3nC5ImS9z4NjME+vxoNgxdtSugs4I8oApIUDRoE
vkfAFIskiZ6WI7Ucxr5qH77DhUMKSq8LNt0P9Wt+VcQEAZ84SHXtf+lnYG03vZdMDhyF8TZSWfQC
l/GSqDb42P2VNil44Sozms3RqvHbcgW/mDl+9+hfI5wIdLYQv0h7HC5OkJiD273TEPBPeqLXp/ts
7sH78U01XG8F8cfjmEJ9fL5eHNov7OIFTqgnQiDvB6NE4eMC/OmHtMrKQeKesBbyjWM1r5wLUfqO
lK1UoWZLNbn/1gXqMewEoe1BzK0twRk0XX1olBdTr9hSTtf0b8PDb6ryLbJNcc4Jxv9DEJ2EAq2H
OVRC9FAIcTckHCjoA8AYFoQ/jgGD2twtORLEW3ArBSFePTfAhdgG32R9inen9NzmPVOI9kQoujXx
9JZgapjkoetLhnwUC/9/zmMeEWXeiD5nsqNoOT8ogkkJ5Gfhr3gEpT/Ujcza2BhffpwJVEGckcJp
depunhnI8eW6h+VSZoNg0zb27QKtXYG9Jg2nEhmALSo2eSQ8HFDWIz4URadODmi2t+SdLIFS6+3q
XkEDr+74kuQBBqz1K2uZBOBPu/1JxVFHkE2Qx9vtOfiissEqMTj2Vm1WG2cd3OocQTlydKYXdQ+Z
DEUvpNEH+WCZGgcvUbhdXNpNih9jR/D0r7Y+oDYSj6zm2HeLiqD5qaoTtEwlLGrfkDcTiuv5sTT1
43/oAdpidICCchNWasJP/MXwggO0sbwXqAUaEo9A3Cyd9CS4PcD5Ew7Wtw3iQufGsxNEO7CQ93cS
F/mWDbS4y1uWKHkbUAtDctsk6fXou0rlQqWgNY2CiYfpROgTx0VnTSCTyOJLcqdekcnSwbNqJle3
Oqn5SuSAQ2L8qfCo/PbsJ4eAkwimIP1dM0ETwxO3JaYZPf6ZhxaxNhAJ+uaCUqNXZRr+2J55NQ1O
SJCHRQhrs9Hdc7z/mnkmlT1XQ4v3WRrE+z/yn5pW75LfYArC3ZmJAP1/1y2kd8pPjwda5ZoEoVaU
5Sza7iSdc0wymYPGswb+8Zi92UUJFvMFk9uJb2YtPyQPGYOWCPAKDO12mrAyVIp9rnyYyCBS4TFe
ac+Tz52W2+pCG2e7j+rtXEZ1NoFZuT3mrKgL/ffHDg1Lq+TeoHxvro/PqVo9yXY0gCli4LHCcOWr
v8wyxWoPx3ZuusAlKeSMn2/q5xiEo6h5bbh/DlMmLESG8uerEbx86ZBsNJ/Y0Qp2cAmW8SgeTo8P
PHpJywojlaODidx8xpO9JJ8XPcjc7VRooycjUSGqZdqrwOpwNTGE81nv4qvOpEv45cdtmSZaJVKD
XKV44YCY/IAmLLIc3ePxiQEDH4xpnDOluE6USe+ulvVPcluMNHOxjwQM0uYqQbsrmNvx36cijUNI
YPcQVAkhwuN1j1o9RVeNCIugq8GB5y7jTHimtsoQs6/lBpJs0DaCBEyImdwd8Y7KrbO6b8cLvOX9
myhUpd2RllCmANgpZU7/Qiq31dB5eGlBTr9LrAEcj7+wZPg5WT8lWsXxQX9+mpP7yi8UgJdLTyZ6
nTp21axGp8QCn8faPRrxNlZk23Lt4jhfnEPEBUqYoGdIRWw3LDirPcDgbQTOp25q9Y+KRJwe7zEG
pVcVi0vPZjtiQfmFRdnWfF/gu+w6xJtIddx12plE+qeDrFokEF1Swj5kPs85Y2xbuLKIVk0F/zpL
StO4K47tYE57oxug5VUIr9F6lh5Wk6+eTGW6EpHBRuixfUzn8jf0rZuRj4Z7v81+H6WkutT3gvic
smunUioXY+oxHcCawz/UR+RzhmMAhAH0s/QOVt4VBIfIFjdhjuWXoxu8jCABP5g8sPH6NxuwBMUz
Uz3RCrZV6xRkBsy09hwIZXIMqgS/fU+CmalSPzYbOlle08U01lag/w5FRCJfOku0ONCCfTrQ+Zi3
9livcHaZz0uZTB7+iVBLsTyFrwdTOi2v2WsgFt73LeiKEDtsE/v3LZTQuenC/HytefbkLuURpJvR
wZqnnlAIIaKfgR+12pqgo3hpmaqmp8zh0yh6rLpAGbjJNh3ZIPI3oFmOJmLkCewiOADYtat5Dthk
DnXK4sIAKwHGaLPW+MatqSLBJ/R8qr/LIEH7HY5dm50qi0cHXXlqmG51kRnLagFmPNhVNU1Xv04C
2slvrZHlnDt94XC69hnAld8rgF2PuU6xm+iWPizTZnR8tGg4ikovbpyf23eNhMZgqcQZXCHmS7JC
QXLMhVRAMEcQ/x9rnvom8wUfQoScGKol7+Dm6YiPqKoZUoUU0s5k2onFjRTesL41+F17q/wU9XET
/Ns+N/fH37HknnWUIRGCYGyHjbxGChXoc8LGwRppoxcPUeggeEV/WFBZxF4kSJbxqjt/NdygPw8u
7FYVqRW0Wb6MnSPA5GKuFxCkThox7qpXtMdWFOAQJIAIXfE3yfKUmykhfow2oqt6vglgi5FJC1ML
9TWrwz6pxQLCwA4eZIZFQH2enmCOSw1wxwmVDzv7EGVDIaGmXl/U1vRz6NH8mOl2J6TiO5P9P6hI
WFwpTXqVGMi2HlIm/csE5oAAFkvbFJirMym6azThI3jxfmN0KncKr0FUNBoePDwwBFlgvwP+uSA5
oSk4fMa0KstC5PFRDqsQuwd05q3binPKJfVshUTEk+8QvNRHysm10dCs4ICML+Zjq1PQ/uV32Zi5
sUfSvxCXGcEbWd4nIWl7fvaHqIfNBMMgypKuwN/6ytXfXPv/jEXSeLFs1KVL56M7tNL6hGaEiaAc
W6DR4ZAOosg5ulm797glMGBLF4aCxypxqaUDM4TFCVXHE0XAkTbXzBikgj8KljgAdaB/PQXw8kKl
G0tM+j4xPJL5zo+CZOjK0N/EslQ/elhpXZWAPA+kA8+P87WOasSX9Y2W9F0TxtR2EwQE2BTDw4MB
tSHrOBQLzPUDsqoHZQtzVwBjbx5trOrWKanmW7FcSj1XK/WLcB7ayCUnbofjkjH3glaQprodAAXL
v0Va7Dmt2OI9fyHcH2/xeiepfd+oPhqMh4apm/Ait/xsCcXJY2ktRq4EewluzS+pUeGIlRLBunFc
vhe6kBk7rqjk+raKdmgyQFR5bpqTbgz4GRFnWWRv8MadTQLmrthDWd+RZJwQ2fk4CKDmyMrStgRZ
UNpkHFCKYsOt3IvVFfcCRYvjWl9WJSZPaCZRsv4ccbZG58P5YcN2vXk1Zo/hTvrg3HnT+qXYvJQs
cqI55O01bxuYjkNsGL+rlWqqTBqioaLzy8bG6y846Q+TFpgNrbjtDVcXAsK9o1IscktdIpIpPDQv
C4efRZPhrYhrg/EPKAu7V5yuMFlT+Oir/rPHtk3Vm92op4YsWz2tFtUlwy5YQWvKSOwqFVenppWD
Ho9v6ENpopmbH5F8SwHo5v9rVXNTqnYEDVUHhaheqAf1Y79S4ghHrPwmQAaSl4YpqFYMd0i/83Cy
JUg9OaLzwrDNjFxiAmO9twtkovP1npszeIeLhZP8tuqbQBvXkvDIhq7u0Pynp+HMtr+EAVNq84Tw
P2sDXu9WGSIA3FlBEUMks+nHtKT73cthC/swuVz0MBbDJj+0w7QyGAnk4rdNtTe6Ade84Cz4f/TO
k+ozVn9/fJjPm1iFDfSaAZLanbkYyNzRzSUkhTXTHI+QkXZHeXdCVp1xUQ3YE5AODhXOTXOiLgko
YG+ioJzODpQRXexuDEnzNkSH5GLDBKfS3DMYRQTqsIaTVDGyNyiO2Aq0eMlmLImugUrzwYg1s2wJ
U8bm0EPZH/sakvKpW4cYM2H87XYYGsG3T+Otllq1b3QqLGRepvpfS08yCfsh+25RIqMJGT4jnPe2
dfEgknqC5UgZBc7siGGiPyQx0nMpZ8maNQekOnTK0kNpYFTl36daEtYLU6EfxnYrdtgRPAn2LPyg
R3/jn+2GbMFqNdmXGZFspcrmBAODlvML1f8kqvfkA4rJj9nO+GJn0UmuX0MhRjiDPm+jZGETXowy
5IQM8/lfgVyJDw7hYaeVI2OOgePQPxUk6S8DZWPpafjkTGsm+ojMb6mkL4M0/GUx+BAfpUKRhDja
jXqpAR3muxXpEA+Z2hJWgMmH3nIK+ACei8MWnSZVtH/A07dtRMsoscPNcEfr6Bt3ux7O6j109JaV
naGMc70nNo0o4uWY9Dz7JEXIHviCfMSiNJX8QyKNqJjhpIG+Ea9EibLXhLxpHNgiCnCFE92NY56s
Y2gfGEV/O7EkUFqJlMDptTUWwVR+aV2eaiEuIuB0pWzu1kPeGT7e+eugIl1FcZD0Qa0Yl/PLChBp
4GmpjbkeLsIaQ19D4Tr2a35vWoTTesfAn4kmfpoq5HCJAXuk+QOmUaT1/jRvzC1bRUgFicOSyuHb
XZkAmq7OZgCqEEzOE6wRg2tQKzrq/isHzEncZrBalxyB47xtvej9c4VE5HWAJa4fD0lOGpevjvP2
YgG9N31LpDgQHPk4iReXGWmliOqa6orxB/NTTuOfrjXavRY4EuVwvorq/U+iObzU1ljjuK7HMldb
YsR8H0hWAhyveMCTyfzJJo0PsfJgrWeAGjKc/jLCwOlL9FR7sQkLGJsToWvWDv6c995JDTShOz9N
Q3U0gimAQPCx2qhWNmJjp0X4s8+iHwMwkKfzR5It7LkcKBawXvNJ9aOdU2oX9KTTQPw/ff2IK343
rHC/xHjAxoEm1r9MHWGeuHkxtL4DQ7AyRBrexEzTjidtUuNpPTH/KkGs3rHKSpKA+CMdw7gQyhYG
+gkXBtOdZSEwwseCR8uMzo53LYu9uBlfnIvGJdhlM6XNVwWwnhEcLj4tMS2h1JN4xVeCzP/f+Qzl
yRS5cvJZd6eJtnfgRGyQCVASYQg3CU3z3WdtCK8mi5v9ivCHQF+dfQlQ1PPqGBxByRfDdInJpWZG
jpCNwwv+mjIRWQS4TBHXqYKjYuoasQcemQcyYN6SC6jvrf2ROEvfm4v7N982Fx3P/j77qEu6Jxv+
h2c1cSgwAcxkpHCw1P+dL3b9ZIPdBP2Uas+W0R4qKcJt6oLLyQmQON+63GvGHuNbZHSwKzXGjvTH
gTXMR+SjYH1ur/3GZK2UsLcPvu+BRQoL71H1h+7j09/3MQ0z/IeXBt77TG2i3hxtGZvlZHAxz0q3
OWGsz/DAnv+JRivSs0CzBcmUTuElIwOT4dAaV7wIoqoF8Yks/BD7U2+lDhxJwuNgLKAGNQMSjDxM
lsSVwCjltY0Lq7aALbW+1Au374b+7zB0R+HuL9VBp8bpUZDYYazmoZFdusAc5BSIpbdiZR75nNTm
61wNE5BWkWknoxq6KDIGbKDRFGM+pwHayi89w5iIwdaTj90tkYKxyUqUVuZEAg8/DWvzmUUW7rJL
JhTXyFGx4PdNjlQhOMaI8YAPJNoMUftEIDrbVfZhtl2Ho+uJcQKs19rPF6lx0pD1Cts5tL7ik0xq
bPF1IPyTHaey/GCzDI1Y4XhcXqhBvKc0Jb5GQ8OB5YHGFDbzUZVyM3uF6+i6sycSOzJRMXxSETK+
evRHNOKz92tWoyjUSsazglNLydP1OsMFLmJA49lClbnHa5LC18gurM+3hahHCsmcvCgJVfZAy/Tg
zYGT4pl9ULSZlFlOMUA/mRdrgGNGD4+BofIBFKImzT28txLEZOp2THsU4aJrlpxNsAeXoqDjjBEy
Lg8eg2t/VxpthoSLAwSmXDJNl1wXrSgUxtz6wY8eYsRyiiV0kZ+hQgVSraoLkHjcV1jf5Tzr+Got
4AqXSqmmD/YQL2S1a1l9EY839OMUwXvCE0M1btxJf6mceLogfhYmnv4cSEi9Vpw2P08IPzOefhsN
ARxSsDeSKpysQ808sdI4PVNSJdqTcBhV1HGvJgI4zvTcgdkdZjatUeyYTXMEXRw4xdBIUzBXqOBs
2Z2YFUIlHnnHzmxtV/8LfWfEhJdHAhmhogVWHvAQVl5BL2ef0m+hMjgpaxlzFci83ELecXZ1SFTv
LIY01sBN3q2kAUxkfGnpNJ60+alfUJkIsTOy3mlYrgxhZifjKPxkaovYTRoomYfI1xyaEfr+93tP
jpnxsull/zu7Ix0vBW9ZO+lm9rk2Fy20PaU71rOVugSL5u1M1HzZWx7iEMry/AzTBhEymywGq8kw
UXH3xjKP45+tOd8O/p7z3A3LfNn9g6DAJUtEXmOxeFYzdESnunwwoelvFII2TZkUyD7c+NLy5+px
UpO9HHnHuVhrvj+TioxJ9dkj3SLTPnoM/E8GbEqCKOPkPc1JyIobugUfAEOMvrb1Jpbkul1I2ivN
eOZR9+bTXMRLd8GD/ePgIbwiQ9xIHN+EKRbFhNXe/dhn1MH+DMZT64i6uRzDxBT/FPlmxMkkrQ4G
D/4DuEP1M4UjJLx7ac32senJIMecelE4az7spSrmoDqRn05KTzcbVJPj6V8kb4+5d8g3nmL+rSr8
+Fyr7xJqx0hxhc20YWJdqvyBqliQvHkwS8JRa7mjpSkKEVVG/2T9tc36CnzDq0+5hIOU/5dr+HzA
chkZ5yj5ONypDHp7Qw8MERl5T1X2Nf39biEeS61AbiwsKgUOu3holnPEbCBdfmBf4YPeltwNmVm0
mcGV1zMBKh/CgQ1tTuP4urLp3vWzl5Xj7Lp7+ECvc7hxssm81cnZmXL8w2ZmdEifKby+k13Xgvu7
yWKDV0dyidDiMsnlsXVhBDafAflw1+ZM2XMqZSPCxnKTc5z5uhjwhABebc/6wfaPP66O5BcFC5fH
DNPT+frTpnsykOjK5brlwwu0G5OCLO1zZwPn7dR/24emXgEIWbtTAABDkI4H6F1bjpfQC+pqWaB1
7QGkA8w95Ra13lg4/uRRT7BL2+QR12Xm2/+uVrbxktNgSf20XNauR4AlHYx7naW1nbabGtmSGTJw
gqeZ79iLrgIn8+BZcs4Afw3UQkd0BbSSaFMNLNJO2CSJ/Q/yZDBkS8mLEcnPyySi7N2XdJfLA7WQ
UEqhHhGQRt0QFIM3iqYec/e7PxVnQyU4JAMr9pHEaBOX3JhDrmaMxFSf7mmR+tuPA5bI0fljiOyZ
KfdSmZdG/EPj5tw+QC3dJa9aSN6DPArzCeFAFIMpuO4q3XTIDKlOi/QGDG9iBoz1Pl8wzK3p75sf
kxSDLoNMacisZqMTZIu3w6bxdf+au43GIPZHVKJug+Nj5O9/yQR5q8W19oTHAas4sU3tGJtywffP
04/Tr4yb1/V/yZIC20uhS8OJ0db4X1vpg9HiP6gSmdgVxp7qpgkwYIpjPaVPupEoUw4ZhJlthdjN
K1RLH6lLg63ewMs4MEHu/6qARYzZN3JG8Q6QqxIti5zu2sfRwYVM7l2l5kLt+keQ7AM07m0RWCl0
fGQBt1l/ht3Dp+EW7ptUxq6890Y6WUGMPi1S44iS2KyHLKtsuE003956GNAiQdDOaYPvoH1yUkcy
FFg0DhmZTe8mf1jpQdDVAdP7Tz5v7gPkp+p0E6gabrso4cvJ0G6y6z1kMCKxuI/xIYEVZJ3PfQB0
CP1OWRdGbMc045WWWsmm8bpLi/JH7hnoHs2qVRBh6EI6yAnvUUaehRewyXXkY2V24F6jIOgQHJAH
5KKD1n8M3A2vQCaklfJAh+EddP+yYMVhA41SEhKm6GLWEMlkK3SbWMZ/HiJ8otC/AdcRMpE+wBdV
DaMAFCquOrd4UJbjh9ILJaR0EgP9sy55Niy+EaLVg+SwRC4UwjaohAO6YCZnocnBxkGqNYinFmTz
okHeef7ycxee0mI1CTbIWXxvIIuIgneRmeh4h/qijU4AyjZFf0KCxj63rbjxFD7KdkcWamxyeLAz
oGI5yOieSyLBbSyGnzbNCmjKFlW7dff5eo6D8fTgECNsPJzphLYSU+ErdisqIRhJUZZb07Fd9IIj
pa0G2dG5Y3347gqRs9yKz2Ga8RIPsIPfcG7BNE+bjTI1+gj1/qJJIT1hQYjIRgY8DaMS9+oKSQ6Y
XAUnYxujSnejCesEun/UYnUDTqLPKQlep92ZAVzfqS97VY2uFQ1LgXQsySgZXwtrK8H5OwlTdYbh
A2peoQriGYVVV65+QwiGT2zJhCfjIvIvP+zD++ITNaaL27gJAf1DbMbjbP7qLiSE/qUD2GM2hJMm
dZb4z3H1l/2S1KIk3k+5DucD0mdvldaXgm9yz0WAbsmBfqLDVVEK9/Yccx7gazFs3GGBPyBk1rP2
OerBFRjpkW34AhHE9QONF8IOp2/YPa1z/ZRj0b3GrmziqEy29dr9M74RrgOc7uhKYCJJpC17PkDA
lEFN1teiykGEB/CK+9tZz/xOIyH586c4grhsHbppnaPK0wrwsnslDwwuTBIhNBi+2hOtb8RnApak
oBHckjbwZN7kDFczoEgxlXHclJRksAHNMJzYI4FJqBg395Un+FOSQ9y3mrAi+hGS2f/utxDJmSdn
JiNShRteXaMEAZs390q/9j+G3yhkWxHmOQwlRmNP8v70B9AwFaffH884wti/zLfhX35nYL/omWKN
urwgbWNx2m9kE0I8CXkR56ntpunSluQh62O5uu2qz07GHnS31NmJxAbNiSWNc5DtGuiwlutTYyRH
mUeml2JZz5yAcyW8Gvji69Emymvf47OmhMKASjmMEnCfv8AlI8NvtJzp8YmKKQjpvyBf2qTZdE3q
L9ibmlSWeEUt25Cjx/5AX2biC5+tLJpyTBnv8JkqItf+PsCg2Xl8mSJZYnlZzRHLkNAKFTD35d6N
NSaiBJwoB/FYEDnnOsoQnuWxoSmNjVAlRSX4+Bv957nEhki5OTliqg9UiRTIq5HEvpMZod3N+6wf
q+N+Ci9nf1xdS9S+p3EpkI72DiNheEXgB769DUifzDQI/+c7q/QbstVVftakiQI2T+s+U4Ij79IW
DIR7fXy4uGzS4aqMgHjm/3hE+N3u2fOJ3j6xbLZnL+yT42p2x05FCyY3T2DHqiWuVR1c4doe8Yqk
Zw4VBUAO3RCN4iOPCWz/irbCNJ1OoBC1Y4ZhPH3N5H88dxZdjXrfahRt//ko1/DEPVeSZqw5/oVC
QhR27nyoeXQeM++7KCBNF+AXqcs2xn0+q8T2KIoir6JYXmjoJq6ZcBucahk6yD3DVGTejZve7pqS
RpMqutXzbDnNnh1vl+hE/KCMfsqmPDktz+l4nSQgr9aYeyelqC8tDJFfXo5mWccRGly2tRT4BZLu
3H+YnbGQtxk765L7vxT4HSvfu8iq4iyY2oPFy9vsuh4DukegG5yw3EvhpN4Ldg3agcFcJAAoCp48
jRUfAsHkGhf+E2BrBICl9AHLLL0iMJZHChHTnkQELwDiLCSgaYepV7kHuPZELihMIWin/a1giUti
MDmOI82H7wOzB8qnVm0gC7FRGhSTZmTsRIOodMVWV+QatE42jf9rCM4Kl1cOAgeOYlwK20vjdg5J
zZWvrWIpiL9cpW4n4NnutXandnnsRmDTE3tvCZjWLX9l4ZcGCFbLXSEN/D5ZC6Kik1QHxjg1zPMN
ecYi8WzexBlYceplZuFhzgqzi8uXpmmjhvQAfM0ckNUl5qh/cK4o310Ir16yudR561aBIolrPNvt
U7paO3Jwk0Tr6Dco7QwutQExDnpSZNXJkzSl8AUXwuAjKdYLTD3CUgvaJB/OPVQ6GCeD+3qbAx/6
VrrCKmhQ1AFlj8yqLzD4tpEqekQnuChlefH1qxZEMJaOP5siBGdXbt+pIM4K/YqMwdGwtG6Za8GE
xsFHKgMw9IhZGQ/EN9rQ5RWWIPsC2BDpZi5jQ7sqAAkDKV1t6IQ2p6Nd+dbhL4tbmQtD1+uf+Ai3
8Yud07Xozx3uGFUXoT2AW6dhQPkEXzHC7RyoQvDuwhSzNTjrD7kRKo9lBkBdFB1Yvsx7Wy+zI45W
eXHfVrl5MAEPZOg3szcYxtAjnrSTvPt2qOsesNXDNb3Ia5EvfWnYOBeB1pZFrx0j4hNEeM47g1rv
yaUn/efkF5WV/xDRURGA7XxSbbE3piGeId3nxLyqMnqXiuGoCgccH4zrll+iW5InauU/RfKKDnqs
wOnPI/cjnmpO0hz2Kh1VDXHiPgqxjtMxgIuuxbt7xN7ji6fbx2wWOUd3MqKeulPtkHDmKRXGi61q
M912y1t0oSBGUCpA1qWIsua1z8F/nQhgWhSPBiqNrfudfaQ6FH4VTbzIRt0y67Zzlq5BK7WNnS1E
PGfSswMjchbg3hdpFJn5Eg6P9hqVc+pCNAnlsjwzVUmkBsaYz7QE8/gphfW5qL0Mz33WyCcedfEe
MBJZg1EE2HEjiV1uHl/x4ybxPvcZ1LwHE4Tsq0Vuyig4Pm3n5hP0oHV/be2EJnaqKFPpsNHycRay
V3nQOVkQTd0zk8Uq2QiGAMdbs9zFtp9QjZtPArCpekld18rujnmgKRFa+OzdcuNTgNGhQ8rMzsGC
QZJh8mn1DE4SPKIP5f5pddArU27k4gKLVxSG9Hp8Q9Yh0t3oAtCZULn7ArhJ/PCdnCKayfEBa+Mn
qAfeDCtbmnSWLbSRjoBf9wmhziMdYLk++w/vHurCJ+uKtyGtyIsATa59kWmsWy7VVcLCVxK5oLbJ
YSyuKiDMDom+IiqrhhlHGCN0dGmN3GEWIYEEPTRLNei0rtoqwAaupnGy9YCa2TE0IPh0YyhNLJVW
AHauRf9E24B/NzjCzlnLg8LxqcxiACjqfAUmHL75iAjU7qHlQOBEk0j6a97ZxHX/h+V1n5yZgs2m
QaKHkUwpGFeZcBOoye0bje10fW8vRTExH5c1hdV7PHPkjM6RzLRTiatXVsDUCPhjk30edVP/IFo2
LRlmzY/IFtXBELEhN/ucjGig3B10ZtQznH/M5Ig+rB+xr796NautDjD2JLckfLjS4PcUFf9bXCQv
ue2ZhvSnZzadpFcP/QYK0tkbiUYPwpGLh+INwgeu+9cI3Co1LGkd5eDXUEQ43ePfiLrlommPQwKV
Zayv81IttfBbx62EFGMv89361xXV2Dy8RpUJ9XJPaZLAzYuE2hMq054fqU8i2r2H35tiZr2yVG55
e/KHXoN/iLAXQ+VQSJYbOBoZ2xAwDUaTnRbkN86fqo/WYVFzBTXrYgAAL/NXEJKLdSsFQPMt6XPX
KuOzpBrNE6PAT68JLIo+fUE+JbicgHP93MsqFcTHSCeZcRWzW5/OzmkOFGPMWzUm3q89IbIot29L
2EQy42a2jB6exqtJx6hQX7jytoG3ZdY6sxV8mqtgw6eo+hc6/JrRuuRj3AwFON/CTbljqGfYsOSn
GPM6oiQn2hComJqguF6DFm4faraUDkzfyKE3aaSsZ7KKiNrGu5ONDeFl0shkR33gnewqvR4Ph2i7
9W8tBw+Rvy6wUH8FtRawBmOkgucAcUpQLZR3ay76q8YijvwOnYKXPgaM28e1IhvvvsMhTHOVYHF2
udzQ8o76FVWZOYb6Xtvk/A1KCLUZSu16/WOsDPd/NDlTUD0rDZa/Bkg5UZXo2LSH5C9okBahr9H2
8CgF59UBmL4XsPl2BNhDRkomyVTy6HHi7Z2oK/CmFEIsBUxwNzMsILwQ3+MN0faRU1699jqfniAa
aBKgPAqCJU1+Tdx/CRaTUXRmZ0QxEOUnbLJnQ+cbykp7EFC5AHDhYni8pPrVlBYa/XMUMatNLY4v
/pLICydi3n4I/zogoqcos3keACSfGtCrxeTS0Y3jqFPxYqUgCSq4qXavOZ/1Q3UlLac36TUAiV6t
pDzLfvcgCX28C1TFFdGbNihZlYhJAWE09ImRh4f/V3iOXpjCp6vqKk8L5PBuSsk6kjH6hzKe4LZh
8/DTj1bFtau6RQMo+lMHKztZj+Om44yzUgfhOau5HosRjHmShfftp+yodh5OXLHPTb0EmOgUqiKr
lhCearcx3RkVzjGEUEeBbeK/PmjCO4sti/hydq8GcLBDkFXWIEFOXCJH1fhFgsDFj6akOt9yjO3V
YD1oTTdrzAMyPh0K4hxnwzjrd8W7dx7v2itBypLU7c1Rb4Z4cZ5xfwmrbxXnQZhk6YPVQbEsoES5
3YTsuttCzPlHm4IAPT5bLha6A++a0MdzhQhZEjD7I2xjhMyyGOhEa5nAZMTX6mXoZScufNPvpMoR
deldoqWZI+bWid19l3PLw+YFN3sbluCt1Tk1M1Hg9BlCwvmu/qdxqrKZ4k+3qTwLKf8GBzOxv0YF
X9LX1GYXtdexn1wsC2PVB7motwJ7tP4Nvm4ieiYCaHHiIKEUNkWcx2D7pQqbiG0IS00B0QUU6wBf
hd/p4pnMo1ZQE8rjCakLfRqIgb5AVnh0iOQ+QSZPUq+Itc6+LTPfT8osfhwhX3IEAbrewBZ/po7K
5k5+kCRLU4wViiHQno7xku6o6vGo2m7I+lls4g7ajMdfZSFL1FaB4pK2XyzBR+bYty6JxMjUOR2B
Qo6iEcCUplvDFz9eDuJ1KAHEJwcLng+wWeqm4GWFZ5BfqPor5lA3Njbv0o3AYJQUak7y2uhoYBuy
spk1dO7vkLeDA46iAg+D8uT2oB50r5nkDfm+Es/H1w1w90V2sGbElhdvbCTwI8CyN0aw0af8wZfL
AwFpGQdcdq/MgG29er7vsXy74m1Vva42SboLg5O+w3Hf0/m9EzESr+SXMjipJ1ZgBe4o9FsvVVFq
jGdtq41isHUpEaqmn8ywPsGJBdQ6KTe/fPQ73/XwLHKIoHU9PpmI0AH3EZFCCEchaDTrsqo9M/8N
UdFa19BvStocg1Dpb1HcttIYvdFtILaoOQEwcPwM5/OZ8pVcnWCmkhiG0Ah7plMAfB2Y0b18RuTj
5vLlUKg/++PMcRNV8YS0q7rPHE9IfcgYQ33kvJR8Zxb/8CBPOdGeHp5SuKzRpRek3pXmxJjQucc1
ixmIeqHB/PASWqZL8zU20l5O3ITw/mR53V12iYL6N3pcFL7m9MB5+jwz0eqwZgoiZFVXBP5j35cw
zJyn8ZIma9afCRlwO4TD3yQGIZNhnC9TxFue0zcWe3uhkhTI3Fayz2/0d8fj7jBL1xH/kvKL4CFh
rs4LoV0AfDz8lcwRxXNaxt+D8Z3duHzx+mPTwz/9w4T05cNvMV06GErJCqG6ZnM1G8TVcsJNB/e3
aUSf9RaC8XrdywIYBFsSzoV9igI4dmDylUXl+2mnC8mWI4GGtY7+HQhKF9UCw4Fh565eCVBq/we+
MwpbuGWtstYVHtttHV2xgz7JKctFTZ/8a6qnOZYEjjIvoQ/YzPd1S2DN8YzUaRwqrRve5tRAySXr
THMRhFZs6h1T/j5Dyo9sMVjPfMuLOIWTQSIkWNsk/IHJisHtFD03eU7Ep9NPZcTkSNtmTQFFQFLl
88TcYuBsTDfgWAE18WrNnfROrVIm8R1KBfqKtcUy7Y2xA/EbW9I/F1lm6r6rp3YQxMBpCntf6ujg
tM9EQRfpBHwrVNJqNmtx+aR6xTAoIylY1w8r92JFQMDN29bmHoaGvGbpfyJzvbq4nbAy40wOMvu/
LmXV8eQQZRPrdzdwBXO/sfdU4L5JO1TZR8gYQ8ujLxRoZNaAhL5ITn3o/HVzM+QXsF+uBQL8YPPr
tEHoqDFojCRR0A9PJScugUAE0y+veN7z7uGjrIld7MumWlkTcux+gSgguwBa9RxNIKZ6wSWFwalI
ombEkPSuct15BIw9iHKVbtZkuuqQ5sdIbeNTeCgTTBhhkmmIlqkI9vCywtZJl0u6wX58pjle4O9x
bJQfsKoHBHWKiE9r09Qvmuji6VnbSXvndnWZ2+45fgoWNXuQbvMkX+FXockY2s+qG0Em64wRwWcD
21lPUMOoC/ZKwIGMYH2PtaqkqBP+GkcYucU1YKmHxn4OG6zUQEI5MB9sMtjSOXmK9u1SjDR1q6/w
WaMdXSTQnAnJmaD9C6zKk7aNQDBRzuiCdZmZgSTUDDY5SHTgxaeYApZ9AMifyw0gIliwsJOZ33Wq
NYRzTJQ8wyw+zFlaW+Ual6RubdS9QGdJaeS5DmlVqbEjxSNMNsG1hqWP8xeH0YGujr6hesX/sQza
59y+D4Nb4rBwTjnhpXUannklOBA2pl00oO0DNezTvhyIziAXCmGWcPEMuxnNMaGS6U747cPFCyBh
FRbTGOSUhThkAAY8xqcpiHPPDfAETKtpDWWdojIwxAKuio9ku3NNOKMxYrqOd4OM/MdyXm1xGrwz
79WDWpkE7GiNNkPH35EMxKZVXYWxaHNJLAApBWBKZLHbb4EEkCdESeN7Nh8k48Lqxbf2tUS18mST
aun00Lfb7QEPYCw2vNdH8h1y5YUVvUSeiF9hIOPEryUiXWhy2J1GAFQor6jYbpj7dPAoDd/aFkPG
M0wXURnmSQLIhipSpUnkIhmHC5Q0SJsX08ZZNyZa4wv2slCe1gEHNeykl6pRhCU9dhf4hhJ/0cew
HsEiFSv+P7UWD3IFuPyg891C5A+WPBhi0w2NYVbMChn64FF5GL6iuwq/AcFX7XQuTnkhyGOX7gMt
Cwk/931KNv4yJQF3A3XoNKdt+Vl5uMX8D5I2PQLph1GiS+t5je4BGzM2PRFP2ISe+MWPSS83ACga
jEx4Rie2XQWJlEbw/vGbd6dXpKUhkkhNd8l4XYxD81l7aB9+QR3PXEXijE79/Wj+enjcQBAwEfvv
vXswe82nZzjwTCyjgxRC6w2wRU07IAnFiA+iIGOIW2w21fCwfslgLJpSUgh9IwDi8mbQOJ8JMoVw
IeXbOiSXl31or/kwJfQGJ/DDHQTaHBkqqfa9jg47khtb/832O6T0wpTCgVA84nzck7+xUrwcOprD
BAJofYx5lwNmA0T9GiJc8kbbEk/Qwh/g3gN49l2ggUBwpoTTwIRCbkr8ga5CUuhS4dqYAYF3yOfj
01D9ski2QhCh7gnFYsUZYLxjmsmMpbJ0GOJEzar9/COBA7SYE53aMM/pvue9cWz1MADtjv6477w0
jy/qMr2ev0tjncslOzzY8axdYeF5SLitKurfrl0xNeRiLolQKBdjMuCWDclsXCEm/SNxUpkL1CHs
zxgGvpYc1lR/vPmmv4YuoEVYfcvlJSIHbEpmHbR4REojuPlKXtKJZOXbfCgN2BB5/ZIaEKLoOKl6
WhhHD6kSGHKvUnvprvWr5WcCQRnZ6clG35QHc/1OCkgwNsW6D6ZRGyAjuOdAjolfHJeop9xCX0F3
d5mOE5BUDUcc6S9x9Cyb6faA6rVQxRCWN8UmuoLpoCroEMS8u7IHT/R4QYHuRqyIBQAkCSdmhrq0
BbdcTLGceAChxv7sroWz/nTZQwz0A6dSb/5mDqMajN9So+OwvIt0UgA2auXVZIdjHxByEC9Y5ScM
tRvKinyekNAIfSRvDZBhH3ShRJNlzvOJ8Bu8KeNPzGK7TIQd1uA6Wj7yHwsSqKjPYHhyeFiuiY9d
4d1JQdDPpoWjRX6fwASeiZCoXTdzRNL6YMbDZzwvlwAmB7A1m+UdErKUXjpyjc/tFeV+aANJRV/8
El/1xOmIn1qpFLeTgCd83jnXoOpZPJ2l92bAj9nJe2bjULTYHayDMzGP2BbyKvscHMI06zAZC7zk
1EWwLOqs7D4I827e7QsG0dxanjt0vYQdWMCFZ8Bm0kSFOEEJ/CkXFypVvWd6/ZbQWzyKddzbtF0W
Gv2SCRoxS45nyytkZmnz9FvqNjlOH9skuNSMaDvNshHGYBps0ctb78oZLYL+UinjpPFoJljB+1it
B044+DgItpNcWhYveBnUmpFRmuyx9Gr2Y/Cl7fT/sg8y5/7vC72rRBQ0w4BHglRujpay/tYZ8Z46
asSEz7q99uTJEfb9hpUuApWIUmbf7RcHsW43PExMtgaDCWeFQtjeRzE1U1TEmZoG24SfklJnuX+E
nqFF7D/5Gm/aoQO5g8DtK1VeSPcxlqaXS3ZlOmA1up+mp0lAbMUj9V1vkB7gNBFo2Rgrewnl7lBG
4YK/4O27WxHT3pipcTyfsfVKTY+Rc0VcNYq7uMq/WZP7L+Df2oqjAA2oYEj7nh1Jd7NQPqAhJNBx
I/jNb4rL2AG/i2c35cNi7X2jweqq1u23cPXl1IVYgnVZsIhK3P2Z2BAj9HWh/gBw/6UgBPmfs7vS
4K7nFx8baXy6w5z8qcUOD8TI9pGLyZD7T6VPkj3MQekwTjTd86xtIW/pW4IhR2dgg03IgI0m0ZEF
RJNn1xuv2xt8aqSbsGOHjpA9s3vzJ0vDg5KTp0dCzraMwfUCT9a5CVmG2PRwMzfvCTMEPILMw7fL
mV5gWF97V8KYXHFlmk+7wUeMfmmhfLifSdiGXtCKPsETuw5sSL9rV+P8h79IytVFnuOj3QMwyitr
AA6QAAsQOFMbUGa2mvH7JV3HFTN5eKSqrUmjl3Fa0bxS026Mb3jz/DtJAbvn+YsKE5kHQalTZntl
eCOYXBzyUBXP2k5XI/D7i1Z+/ObQ0la4X5DQXXS1esw8m4V6QSMfhzMXQaSRrWhnepjAelDfUJjm
i504jNceG4t8xyNGQIJ3aT7pnQWEk9kXC5szNUeRUvohs8cvgbajT+FbGGU9pX9e0n3IEp1MrPPk
HU3FPaSdubPCrA+48Eb6E8H6AUR+2++ClZKhUI1a/m85eShxMIMSd5MkivSp8fq8JGVuahTY0KiO
5PcpGJTwmONPHePi0yKnsM4rHq+Hu9bdRY0LIjdBfwY+oGsK9xEooRz2szRcOVURbuaEqfeiXoBh
FFCFZUYoY5rWTFr6NCEtDKi5RTneyLGbByNyk5OTiyJ+b/wQLmZsmlP2mXwHSmuFKjMNxfAAnCkp
7PpuSVMR9oBI518yEtYSoR7YoLCld437yL9u4tC9dTnHmlJXKtHn3Z+YyqKUNYypawzoRm7EPcjO
AfJd8rAA96yGeZS3SqoGPgSN59aFBp59VGp2xN0RU9tPoidiVMbIZLVdNixsNsCbkyFuaWaLhy/F
Kc8cz009o2kTqDax/Id7lbgB1qp3MbgiUKm8tx0y2IV7q4a+Yn0EIaWgkCummS7/52DxY7Ktjz5Z
uqb+Mdc/HD1wO4GsyYRwEYqI99TtZuMDB6wyJurgePSsWpPjxpLJhPc4Z8JZiezgMXum70XZQNn6
wfg6/w1N9mN26/R+R9G2lQSXCAeP7+RqUihiW2wP/j3BDAXqMZTFcnLt6xGzuLh7ZWRSUgrycXIE
yT9hy/tRTUOZWMpibL+HUg7klFLQOO57aOsQ0wOq0yUA6XPxkP3j/FZFaRRNYNPGiziqxUrYBMd/
lexqZ8BCebyWz28baZSjln5rQUj4tocko/y6Xk9FT7OFc/cdMeJHJijz4iygWirjzYWzYA1ccKHa
NVO+MiEs3gDRRwVf91x5/zNtL367c2nl3wiTKP2wp3zAGhdyf/GX06gEH+lHJoEFq0zH931NA6cw
OYDePStKDQeSkXXD6C8gwRzI5+ilFRFQVBVIJ+wMpYEyjctQctmGCAUIbLE+fOGMqI72Wfc8K03B
X/z5nr/xqa0nNFWITZQ60ytKsW18TxqqcMpZKSr73w63UnVBm76xy0EW+Dwb59rJPVPthxAw5Si4
SsbtWH9KmTlALSmVZGAnPOhNDhjPNF3zgfy4faG9LGRBtNOrBWXnT4iSaJH7O9ycsKvhRY+BJgX9
BZq/R5HfVqZ4F751BP3pY9Ayxihx17R1zmwxxkGMYdqPoQ2jk1NxNy72Wq9aOu1tJpX56SBDmf1h
aXvewXNiD++nedX5rwjKzAh6Wh4a3wHkFDkKi28lCnIUDUv0AzYBobT/zSMMBiGKK5sjqsP5rFwB
NUjCxz39xJ7tNUo+ca2qSGYkSNWtDo4ag1a9Ern8asxq/5pZHR/yKUiRVIhb3/WGm/nqnbFkknU8
SHEeDuvypkvBqaK2Ta5sEZqU6nVhqo249vVF6j0W7CNeYWYKjOePDoQz4qD93BGXw0ngSYn7LG5I
3PID2jrU8qiPXM+R7b8iwOD6iU7rXXNt0/Lbaq2gscrdjfnxuCSJsPBKUZkXkIULCBFwQ3LaQPCw
pRfIATTyfJHxRkKFB6HUJaCl6cu1G0dXgKdeUOcRkfWR3lF/X9y3fINUcHFhEWXQOZa4HQC3Hw6O
gXiALm5/KeFDn0fPgzn4+6SS8c6ldVEL4YAA0sdyTiWLoI1flCRjz8LLjCXHZtAiSFAwcw+iQx63
KzzAMSGk5IBeWVfpgSx0iIcp4SsLyF55Hk2FcpomO0dsZ5njhZZF7/Uq2gDxFIapn8zgaczXsKqr
0liVr/7CGNcVzEwiXYOky6+mYiTALJvKmL4xkybKIz9e2X6f3NPGFOYkXtBHfA0twZllLV/plKX5
XzR87UvYmonPCIAnUX2e8RAuue+96c/qbBf0E57nAQVprZ2+65Vxg5Wu5ASoVHmlNOU/imHp0ROf
EZ+nb2hKGqF1ygu7wKx+PQkeQh+TNgllYXsA3U29vJV5b49hbY704o5Dl/O/zIKrCdT5LkasJeKZ
M4jOJ0AZsmIXDzdBTaJTvGKHU9UPafKYfBNLoCpqKNgLvOg/8RnshHDVtcJKbathbJdcFj5TolSI
jyHdwvywZuSJwJ820d3ENMS6O6nB6QJWwlCsL/KSHzszxulnD+Xl6oge9gXLA/ZRcLiSjVBSn/QA
KNmY5Zgit2Oc4WnuVjRKTJgF43h+SYjDP/KxucRbKFQW3WEaWqbhn3Om9nDJoipBoiTzGatAFAZz
zcIRBn2SPo2yMlrAgQO+wb8z/yvdTXfk3zGM+Ql2hz9phsWvKJsLMwauj678ZD0EVgJZM8ITrEWC
pqe2wWuLni83lXg8krY965B81cJVIPH+2tGwmiuQzVWOSgi0y7zmboa3kE0FmuDxxIHQmqhUCCif
pKf0ALuhgRtGswqM4dgBLi7zkuYpvlAUHZLMGPgZuaesQJkTVECGBsNyIOlQchswn4dbZWEiINp2
anJZ3yRRXkH5qGljdTXuaa0QSONJE60sHvO3u25IxJqhoRuAxzAKTc4o0doEiuyVKAIUiiVxQTp4
BQtXcrpb0GbBV87wdbj+O1D+c/EzyfieYDTr8j2gjGqUEnkVw9Msp2IjzFgvXuhVFC0WZVHKLXaO
lOA6cuwoGVKeHHFOcdEh6tdaP9hnkVqtoWZrBC7lK5xdWTSE/dW/05wz9tiBW/44L71d3pP2BR/i
LapaLrTh2KsDdfj9mGoEsZUGRxgL5RYaaLSMrzbXipE179oO2AYvnKtmi+y17Q14HkyovRoCTfiI
5HsJGjX+sZH+ZIky/6P37jm8te3+hW4sB/FtPfgOzFIts3FE57MNNJ5Cn2a9xYKWLaxPrngP5b9J
XIeG2W5k0cct2oQ6zP7PoSF23/G+hwI1SpCUtNwOW0Q97lMGGxjhuMEtlr/seYk2AkGftrUOjDqA
pNteiT/1ps0X0KO8s2G9U+mtSp0FiQsDd2GkpW5yEIGsdXtm7t48OczxLN7mPH/PIFUPLkPoY+W/
96WHaOwFJJI6fh65I06U8LrypykSQHwkeW44XKWJUvtE0B2oAvsynygd9R6Fa49BNGSQ7IWrPiYr
wod9J+Obet+92ixyyv6xdWqH9Uajm0NzHHgKczyJ4iDKd+NCWhPua6fZ3kZLuGvnKRBcPbxCNxIT
gnzFAppbeiDsUqCrx5Lu15ophXN2K2zR8jqfdluEU8/B7PY29RcHYzGfQseujZ4gwjXM5eWbQsdg
lAmzO+UXZSnVVOTt9vryAmYxmw7g3oMExnfQBpoepcbmj78KMzvXY/fRBTijvyNLzCI9JvIXu9/7
bCLBb67gjLiDW72/M6rkuuNpv8oJlnRx6UC8aQBg/CKKaElX2WbXYUXEBwwus+7eKSgsMaXGPqJ/
Kdm9WL5qvAfHp+G7E343gs7GbBjLpAvvfcpKYLX3lHKiJmav1AzIWPoB+1VnlvPV908ThfnZZ2t/
+BCxTAB5Jd0QIApV1hMbtutNBe+1rB4nImSl6kaRv4allptX/68dtKAlBX9OcKtSW+V24KDzPuQF
lAmH2OdAXsKwktqbTVhlBC+mc/NRk4hQoXqoiqzhdiQ4aeuOdqfO195IcVidTqX70ZuAxR2WPn2Q
HoY95nPtM1tttUIjnI56Zj7+8kB/v9t/z1Vqcevkv/Y0IW6W8qgJAlowb+nyiCHe+PIM3yvUeb9r
OCHjrdqa6FDfNEop75Yc1VzArEimazQAXmywJdriYAMoe4GzFciYOnEROn40IFR/NySiN7euc2oZ
QRfJV9lrG+q3KE0taInTBpxbfbF5GftuQRDODqfzgV7f0EExJjc5IU6VVkaoGupiqQ8fUrNavVQp
0qURMEzeGM/t4rqcTEI7QSRJaqpstzcMQPTeSAxiVuW1LiSmuXRel0a4iEXGO46pYdKdsl1sDvXy
ts5/ZT/Ie9oO9j5J646NNbCFS5HZscJgGS4xDWHN4GuR+FfmpPfGx+Upe3D2q8PtGLYno0xAWfP0
mpeTP+f6nV9fGJSMB12BLsSQjoWAOxsL7XhSKKM0VCndh/nCif0U0StyuX1HlfKysK9GleK48wpd
F6gA0pDhq4wt2NyTAiTuBd1Me3wLFqEVKNXHtJTjGFVBYBeQPoVCgaIEdtipZnk4lgKIR9EaGzzM
IBZIHhw07EWi3o1b/3wrQW11RW40rTzDVSGQ/vrht7XJ1IiP60EpF1JJehqbX+BsFOtY2AKHZ3S0
Yy0ism3pxIdwAGEMTMyvGh+HsBsgQjKqmNzwshLg7jghgB6Si8w7hc/+yRu7AhB2E7ZqLFuuN6zG
8bcjMs8d2AaFBu9XSWuZbTZZwmWwUcb93BB0j+oWeIDSNrh0/oa8EFzQOIMhxA/5FJJ/5BNTJMEJ
otzDpiJYN8FtWvbXYWUluZtZRZFTL0mV01P/UjBqhOlCkvN/PN7uXZg20zyaP3ghLb0wJGAxfSP1
10jMHEoOFmsOJw0jGNIfrY0WdwcCJTVziECyIJ2O+H78h5+ffKzVTTYE2Xs1LF1SeozJbHj2Ws9f
oLn/PIkeYrEeO1yMLe5gbfJ3346xLLfwCo6AM7AxLM1w8fc1ZzH5Zap0pCNy7iKmBOOrcpYdrEpF
4iqRcYsxRCrh2gyj6gqfnnZZw4GRzptbKqgNIVPEYmJJOFa1rd5aXbInqqw1/9po+f1k56DS5xyB
LhMfRKIYDDw8wY8k7ddz/nffQjuS7jHrOl+cA7qh2HG2xcSs9racSoWjscD3BPM2FbMHSQSqh/xl
ix64SQYp/Bh7dBeb1VzxUUJvoEUbZCRoB0cBEMjRfpMwzPSqMoRNzYZpQOmH1tT7+m4olAvqHta4
I/LRkaLulXIB/2YoqlFQv5JJ3bs484gnq107UFzhX8uWZ1sGew9Em9X/AvfQnAJL82OV16Wb9j9I
+OYEMzDaMW60TYLRKWdKf7lxpenNYLWrWM7W/gLkannDNnLQ9bFRkAMW7iJStQtItTLG9msXATVc
hYltLO5SVQK7qGC11XdHypxQIum3FFbtlYK5fjZWp9pHN2xYFzPsdMf/q72yUB+bezRONOrN4X0t
k2MGR4YYpxHPT73LlQOj9e4BzOV8Y6gUyJcDt02M29ssoOfslBxgwloyGXHEKxKxZ4Hw8lLnGKln
0L56x4HOID7qkg3mpUFQp5qcbisO1sRH4DH725eagS+TkjHUTXC4pJaxibb2kXJ8jO7nQS+Nyhck
YoYzXBH0hZp9HDUe38b9qPG+crHVRIzK2vCK3T2pf1lhMxrO59bk/6mq7HQkPl4a+WWWDOVyJpw0
EXCqLxwGiLf+paX4x4eAHNJKRZf5lpXCqTWpQ1BkGyLLDo4GLiV/VqQr4VLiM+h+LOC3u/iB5sTN
EbcenjAn1I0+vMIxYLtoQgoEwzuzaCcaRBOaOrURp+Y+nVMiCE4+1OYe/d2BLw50MCNE41AqaKC6
Hmc4iHl6eisUQ7qaZglNYo+daD95KRsup5jsAIQtOyhxulLdP+s7xu/gcWXqY8IGnSidm8jUQov3
XtihN5m9yKzgMTmxbEHWMoVZ+KU/727oRtonMShFaAuEtKJQSsvmkLILoWzp+7Wr4thTzHNfq0+H
Cl4P/cVBcro89JPMHxqaPxROwVgJ/Vhz/9Kp5PcHzM6o5w2vMRsK+9G76oQ1zKbvVbeN8DBefsY6
AQNr8Lo5quEG4sradVT9Tl6XKYErkCE0IFc7CHGY9qzqAxf1StM/+R+nopy8YGhx4MaBdYd/7bFs
oAOeaGFy7r63LMpvWZ3z/M4YYXkf9+sIspFSvR4Y8SiXd2GE5O78RYy19K3aXsiDs96wUJlGZsg5
uflqrHuPG3zjJbOQKdASY0wpSqsYNnH+KG45i50Ji9dDuZbSJ0Zr5qm/8ifqBVnif4elRVh014BD
AwJMuNLyNYmLG7rwxAFk+0lIlbrDqcm2tSdZTRiY3n1gT9r1pjafrBHElKh6G+5/TRE3zGbs+Gy2
zN6Zdm5gzbkGvjeThFc6NXYPHf5Ug2yvAOE4rUf3BijXh1xu23eDKSFe1vD2zgAiWsPiyRg86AwS
XW6RLG0r36krWxBpb2vahnnEV/z/Ek96/X9tqB8+2h/8zB+3kJnxYyVdVs0sa+boy6n5kQcMrar8
Y38Ir+UoKMzkn/5W2wPD0cbDOtNAnucssBzWN/NrxYJtQSfWU66d17YaSVpfNMC0gsA7S0Co8gnO
7BMoY+A4En4+V22wtuW+g+7hUTaH5bpohU4WJa0tqiSt/kWK/ZIow/JvWE3B5+brLzSCp33mLmNQ
r12KCs3CQg8d3dA8VrC078kG6dhC9o67jRImwn5GBUGRSoHT636yG/QCq9cAU7bk+WEwDZvenwrH
HKcmN5qPN5EXEhnS2ZzEv5dLAX+2MCT8SRRxNjj/PiBKLqvkY7/79osFs/QwCAab+oDJ0P6+w0md
rpkSUYxZRO1XAi6ymUDy88u0VaL5n+y5SZzb4UvOKk44o0RiUcMjpXdGIm4Xto9MWUvwZrHI8KK5
dtdlXcw6YFYKB7p8wC04Kh6hViEM8NK30SioypV/p9BE/UJ0afpr2tB7DtZq3eN94IWoYP4ENG3u
1TeAdHf6lgqJH3WCYN8CTKNqI8wHRUnNHJI1zaMdO5yFBdr+LcIp8FNmgdS7GHvXK+oAzSnYP5vC
0ztttU8aiUVGyGv0bHcDq2ighC9jLGOdqqUOyLeF34Pe5fG3WStuBXMPQbsXIeUE/bBvM8stUX5o
59uUJlcTJn/MxIo5JJG8wY+3R9ZEIRRNjC17OrvShBNI5JmQV9neA7lwQePgkiay7KMoeqQXECxV
T/CH9zSZfGTjrkxBDPcsVQuf/J59+7uFZBjNifwLkRKvIj5KOQWcF6pYh+jTwKrsGnmJeNssBQLX
rL5/yoyH+RyCdPMUfSRiccwhNIze5BdsYA7LbNJkH44b5jtMt94V8Ul5LOm8BZ5cuoXFk5dB4Ads
XDFrSzjQ0yKcs7PXKMCgDvB0rNwtvKy44AaXBwuUN2bS94RCP4UyLMW08iJwGHyeXEBDlRebW4LS
HsNiRJAJgu8eit2Y/7OMraATnMLotMos7lDPb3HcXHRNEr0QpSmBEixByMGl91nv+zw7Q9T6ZOIm
iN61vhc4bzrlI9Acn+A+RgRyBJ6cCfVTnvOdHuQVY2aL4KVvKAe2ydTcdhLcDC0kDr1SEWGpVZpN
4fHw4DfwPnUkHvOEwThaX6V4wxDQDedlDFlnwOGZdVYPlz9nIb27TY7uOiccKc+TT9WB7z9O7qcU
0bSuIm4rKyeuXuqvLrUu1geH+6LDpVWij2WODZ1SCWhwu1664d97hxGE/P2iPJ52sB2MUDnC5JV1
4GlyL3Zr2xty0wX/yTEuf1Fv1QNNdTjFt+jynDOeyqfgwKrmaLLpq+7HEFAYao2EqXuK3MbesH++
VqxgEVi5KrjY0wzTSfQ0hLbodtDduxLEtp0/7GXMxc9bPC2w0RbTqZrHNcVI5wtiZL9TFRKpat6m
7sSz2Oobq9q8nnnWR30X3FEE58WCH1LCrTKFXdtLPHzGOyZIAkZDdoWLGjRxxuj/wCdO2md2iOz5
eDtSVPDlo3B+yuxSKITIHpE/i5nc8y03IMyol4D6CJ2CJiDtsDy1ESNq1QGp9/BUwZ2X6JgzfqO0
DT8G2v4Z+9rSsRpppJvab6FchLUlKSBhA5mVmJA9Nl6aJapQOD/2vTnucusPRN2mONVddPEntn0l
X+vduIo0L6MDQjU4cUd7IvBH2tHW/AQCg+KnssQ4OKizHIiX0RpMGSQlIC5SG1t/PooYfNcNMA9a
v9ndTEUgVz29c0cpNzH9KEqT6eXUtpxa6Y5hgEm3H312MbcNHMZKqwEKiFdXc+nhWdoSFugK2KpG
Lmmet3LUeBQHBfI4McyT9KHgW9Pv5EqFdZCi6iideUZ0IsT0/U175U5AQ+e94rHeaOQfCol3mt/w
8z3UqJtStO+x9gyxJ2BQDLKSGWfO2gyrhcmy00yT4ll0x+ilGvNPrY5uaJUvkDzgxPOAIvt1CqFP
SOzaTJ6Z+mMFUvN4JJMKmpT/eQIozQ72XwYQnQAMh+CqMWUKkz063l5eLXjzPmfeZa1rvujSGMEX
0ypYHhn2y3iycIP/Nt7+q7NGfB7/5Fta5V49Gk2C8gQHLkqX4JPWwME4ar/rqxVnRbVk1Relb3Zk
Rq3PMfEslIr3b6zB+9YR174cWupwqvhiv7YQoxVwT8Omv5cN5nb+hP27/VdYMmhDe1RmFZ3JSGeb
ZroZvcX/q00UroJN6l/jcn9RoHT3wCcnvIhWuopqYmerCAkm21Tb69SiYPDLJm9hlsdQndpNnjFv
cL9cNEdpg2VXvfJIbZxgFjXBPF+rBPRUx19JTzt4erz84w/xqwvyzS042KxOB8QeHK5Uyioew1bo
yo2Ceolbt/bTq6N+HwllfZ1OLHedtRifZfpt9IKGpZEDXpfJvYStsYSwRn4mStxfO5vpZClic/T1
1EMyCZD/qkbnCVEp6nC1miWqcX9pXZZl5lPWh9ZNu3eGufnmDjlGZ1lA9Z+pB/Apj6S31F2/m4lh
DGPwkGkUJdDm8VVhr2159+gtQig14Gx52Gqqpp3RhWPewYtPHq1Dxhtbv6wTcKUIEIBBXYZDsOcM
tSutBP3m1UaTz91lKHMOa8fY40wlYp7iU5zXzA7URaQHwGy5xZlwW+1mWWzCtzPnPWdMhARWrZSQ
h8Qqa0PrSXbtcDDxS2XFxJp8oGg9aw2louChHgPGToNpQVVQUSoh3KUFdRMauDsaF5rJ769Jsoi5
4Vfa/Covy1Mxl/nI+wJdGqrqtDQeJ3bwhjXaJ3Xp4oJV9KNzsM4JgiP9wejVTe8Lv3AU6Xl22l+2
n06dWsv+EV2jcaGwFRMHe907YDdIvSQ9p/eEXkcQiXpayzDZpE5lzotmMkzvOUTpvDmfzESxkJQI
xFxLYKj4DpxiR9Ag1YpXUulCgcRApi70fZ7DIWJRRJ85Qs366qMt+9t4/yPy1utyvfoOMnJmOfS4
9mRmOvpyQ7DlO+sIqv6kQBeU89ilTyeUyst5dBjHRQtJYtKWYIS0KrF7JMRx4f3cmfZaR4Im6+Qh
nXDDoMOqUVZqZkY6VxwbMjcb1CDbhCa+LhWbPKgejalP3DWw2NG0j28aJ6lBUJVK8vxzGxsopceB
erbhnODuV9SESAwQKhinOLNH4v7daRdkvrnginF9lhFjuwwg975HnjAIv/+WcD61M1Y5IUyuryAc
vGyWJnlCjwNbLbQMami88QOvaPnwcvNuS3B7UR3fCzDsQGa/O4RMMoMtL1t/Xlcsz1AF+LdG3NI6
PJRCMFLs2Vmn6m7jlQh0H7MmJvCyMJa/yXd8ZeMgrTRm03Ntx5ThMPcJ9JaVSpaEDm2xJ2sTMgOs
I0sZ4eznCXIbGc+xVS2qwuVdgAfOxqHGXVJHz170nqg1VY5UbehRVZ4eYnwoW8XW33Pq7BxkjKvu
rIGufFi9/xwdfZhrv+YSoUrbDyuygHaxuWN93n0i0IQzi95VJgBCI9ImHXqV2IHTP1Ui1jDLy02t
DJGgre9NMuaz7x5JiNg0AJrBPNFUoay8AkwA9sxrgrwBTmPyPoAUJZTXs9UzjOxNQKXXKJeBiHUQ
3kJy54HvT9tW3y6vvmZQBmdRnnu8ARsv8sMC0Qxvx5r9GVXA5vjuS3ORI0kN8UmxG7cd/0u2zWvO
ODXOr7RiT2CsXz9B6x0FtYEMNHSLBVmLDhZU3keSesq1qWeA/b1HFtCIkg49RRTsoRTgBk4HECpg
ksdoEOg8j136RfGqTHh2T6RbUMqKtfxQZO0kl7jg/qZl2uM1ftpbT//hbfY3LjIZ//q/KZPW0Gti
PYeyPFmQo36xsRyNYn0RJew/RPsCwhbljzIRfMazVb9iFiId5GrpOISXZBAT0gqqqcCkvYYFb6zs
mLTuGhaOnzBf56NsZ4KDLh+2ZnG9LiQmSSZ/6JQaC5WRPMZHtRs16GQ7VlZHM55LpSAWkacjEQQo
46v4OkEUM3HEtVFCK8vX01OjhpIaDkocGtTiyC3VTTbGfn7ezGONXAkqx/SZaGky0npq4YWzn5wN
99HnbFtslA08AHBRlQlATDCA48UWU3BGIW7vIGdaEG1mIQDLalygq/E56OjylXRwx/ibg6RN4AaQ
EGC1yCHgIOHMDq7wbLOC+cCn7bdZNN7qiLjcCazJgAueWxO6M1QlJxtu4AhdUoDQT2ffQ7nopwQn
hqEDuYWLYj5xiFW17i/d3SKkake7o/5MivqGo1s9Ss5+w0TxnGNRGVUd6W7f+6idra/W2CN4uI7h
VRAQb5LIlZZaCaXCe0V7d3n4BD3Q8LJnNmJqzUpnusTVRcj3BmvyOxLr
`protect end_protected
