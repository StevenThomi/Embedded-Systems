`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2020.3"
`protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
IQHB+CIKFsAFH9iLcGZD4mWVRDfZidh9vdBxwVRdynqY3xiGlUijBcr1+11MXQu4VXIvL1/m9ch9
0x58YwSukw==

`protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
WdtR7fF1H8L9aDf+mKYTiP4GkQRUQ4pF8RFTnvoxNG5slJliPPwSrmqcsX3UXUIrLp3qjeQDH3he
PTjnkfEIMR+B9g0Brlhnc3OopXUpMLeVnVsaPSa0vyGPT7RSKAavfXbU9V5AymoDvLP/baxjK46V
bw5ge35eGloUnUCjxck=

`protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
vEhheir6ntY5gdOh/GMlA5zGTVpf2tH0qv9zdgSVT2CeE1TXCyJl8rJINMVXTTf6+xR3nLda933n
ZP6OE1OXU7j+CvyiVUOoEwT7nvVFjlyDnunr0P+X+9Id43I5jdtirA4eEzA3Tc/uR3HTZMyyonp4
h+FzxbmkLKwKQOq1X5GCTzmsAYTksCTuW6meeTQTsjZGAJjRmF4OK1RwkdTHDhUzo1PLIxG3JMJO
FPCBgMNVud17Qvqu0HZeSCEvffB6mCBRftt4lO0hRw4aJi2Pzp+jTbxoP5tPruQVMU4++wnSHZie
owE24VSSOW4clTP1+wnIhMoL4F1aufK4oupEeA==

`protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
IH5N46D3qVRoJlCpYMXOW7CBK5y8/FQ+IAT0ZH0S4BBL5qsRHkIBtl3Gn2NRIgMzLeQ8JzI+llVx
T+dYWeP4YIco6bljHyLqoarL2le2Xyhf5utwrlbtEguHT3aHrTe4Sbi3hBAxV72C3JVE1sISCMj6
i1yW1hQtwjgY0/smY15fV1JKc/+wi160DP8OczQvPhPkitM/H8dvGwGhxVbdnPD/2gnhpgYqLF9h
abVMjbiDK1uiKd32IPQou5R4Dj6Qlc/2a0qGWXnHzAoNX5lpAXylNAcwzPcOtsQ7LQZ6HCVrPyCw
wP8hoQh4ApUkJibmngp82sjrfnHY6D5lj7vzmg==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VELOCE-RSA", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
BIvkZXEYCWmEqKtLavgsdLxN+vJiT/Rq0io4ou1ORnRT4FXu8G/HTTK6Qosd0S4pcByn2K06ATHm
4T/amR9WdXdDN6BAnEa0PZCepKkwJI1X0IKflPwIW8oxoyfWcDh/swCavxxbkYPhidr0d6nOtk0o
nRKxA3uK9E08aWgO8bo=

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
b7MY7iJq4wtqS05GDYpUAmbkGoWOTaiVCbkiajLW2n8tb8eaGv/5BjXEC3Dc+Gv/mXE7IJmDoWyi
jPP6fi78t6SVv9Fpr+RZcFNrXiQPC85j7+WmqkPTA+e+z6a/TokOe3BWs55IrfM7EB61ARI17p3r
hN5igHWaMLVnJvkC/nGav1pzHDPBYfsIzBM3Jg6BoCZE+rGk2CglbUyHR+G7ipDyil0Wj1Sl1gOi
D6DbLcpAlRwq2eWnwBuIEZyKWrXH+mtvcZpLstDvcS8oKhrnAqOFQz0eI7o+SxejbbrVBk/7YlXJ
XLTr0uSdHHBuWZZq4kyojOOH9KVgX9haJ+l5sQ==

`protect key_keyowner = "Real Intent", key_keyname = "RI-RSA-KEY-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
m5WOmgONfioXxSFwXvZQNmst2GJZVBRRPLArHgAPT6YPMbxu7R4G29w/QXQxYf4e2MT4EIk289IJ
Y7GDx2LdonZuugl9WpEnmRp0wmBtsRZnN8AdWRJ0iZb3eEpNYk4BE6FigTspdfmiuJDZ4BWIYzfz
5gd08CUe6M7/siN5joqcna35YngpsC9ciZn9WOBSkjWZCrtyYXZD5EHQBTYm7joDXy29gcjtt4mP
bhkzOuRNCWCqBrPpN0nm/1u350BjThlVnQkR5lT0PORql5x3lRuTveqaDVtegYSuKLZiCL+8hldW
5tfsB9IdMa379kbGmXSJ4BZy5Nv7zimMt09Idw==

`protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2020_08", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
R4rNp9KCefSDxfXjAVj/jYeuNK/8HvU7IfkbEG3p/k/43SD6oLfuYEJxJzeVrqcccDTqpNW9PC4p
wzPNDFky648C7TVSDjF9KTW5bN5HU//Uo4AOlOHTEazrMwIhUZeiZ1DFjrR9rqnufwcpJvqoGwpn
YLoKC0TTqDNV2S8B0OziOB1TeLT6Y10171UL7uHu3Wjm8C2w7DfbYSj77xhI6hzn8VWSiCAVfoHS
FAYAN/D6vMDRS+I88MxwD/KU5z0AbNStFarQvkUhQKIMeP5VTM3Dzr82JWXc0Ee93MLGUSOXkYLI
c+tc10mrnyXQy+/7iwNpb1pI5WUwN4WVYvYxwg==

`protect key_keyowner = "Metrics Technologies Inc.", key_keyname = "DSim", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
OieoK030HC6U0FgCZPOXTQKk7ztE/kV5CVJP5ob4m8NNst64p+IzQ+dZebidkPPueNlAKAwCju8D
D0zFJsNn86UlnPb9u5ljEBJkwpp9qZ8SzHK+GhxhsdgUzxINa1svQe02vCsdyh/+WM9nWdC+hr5C
Qm8MCVOwKngdPz6DrsldxdWLBeKXiEKEgm49pHibTkmlKGJqbekih2zkjLXIxiw5LIp+QHnFRlf1
hUR/TioKl5OALM11WDownJpkdE3JDpbyPIDmvmVpKJr/AAKzX2PQpOXH1w7kOuWGwOvIYYWnKjit
3I/FrETJX3Bn/sMnNTJ3ZWIwmzXseKdMV5VKqA==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 1559120)
`protect data_block
b5ubrrk+BFpt0K13zpClk92PKoMzMb13IwQLmUZQuSbPbWO8O1Buv3xQ4eCzTho0cJSr8Wdkwd0G
evXZ22Kpk3NVaHuMbtEttkywOrwH0+LG7T8g3qgt0mEpeboH0u4LOX1k3TeKe17+OBuTRG2yeYho
EpHXrb5E0rNCM86Crr9k/Sn0M1Lpu+6euRqcfP6CrXDzo7f+gnTw8CALWiEKR/OY7xRDLSIYQxTi
ZlCcF1/uGHIv9+5uIQ/DOtT2hIsjtgwNjNq+Wfw8nBDIt2nGMwawLLzA5dwXElorM3EiSC/zOgFH
zmpdzwoioIVvmzga+18ho/2kttanNM8Yy2J53drNubmxQ3J7d4Ch/7+XQ8/sloxCtKAOVLsPS0yV
QfoZ1lWj7Q4NAHKmNlUc0WjFFK9bkD3Av0V4TchhQZfC4gWwxYDSeBXYY8BXAbkJ93svngQQoQfP
vE5j2CkW0Rf9Hi3INIgiA1VrKXRBPGvY3MdjOL1czCKl+LxsFtTyZaIZKCIuuO79AHn6l6umNofi
ZEVt3Cbq4UASl1dffO9OMK3JraRrjfzSMC3Wlnq9MyTraJoUN0RzR5+Z4d5Dn3u0yQf3CRN7kyok
VI6L/+PoR8fLBwU9XE4YN03YPP1zCywYN8aMaSLv+Fb0JqsnO+RLuLCl/I0eLyo8fombv7wMzKIj
MoJxh6Vu8Debw5SU3ooJMx75GPNBQtrGXJvrdudvJHaueEWCaSt2Ypp0HRQsWEk9WAGVa2ieIkE2
rDYvNuYzP+vDBp7uwGMJhqoVdWkqg4pSQUXNNDLB0jb/mDQECf2mhO6ZVKeoUPXYJh1+c3rRGmI6
O9uvgcFYJxaCVb5iSTFqSCVd8DQQh15nil/bvlo7Qa6zmjguyKR7q27KmdWI9gCg5QyzaeNNBnbf
QXuMpv+qRUPjXk2YBI/W9FWx2nU/n2Tn7HNt5XYB0ankHvNfP2isLYlt/jXQOWdFHBDwyDfjSysf
LiAZBE38Na43MKqirVTPgg300WoUFbteF73DgwgTg2qOcGwcaLt3p/lIGx+wDdctVg2rfTlUfVlq
B1Okx8PVEA3hDvSWIZZc46w44oNo7H+AuZ0k71zEk+Og63BoQ7b4Afy44k5GKkELVv1tTAcmLlT9
vhtBDGxAYvJtp1JagfQdNldap6TiM+VAdxJGS5RQKYWW0l3IKHLbV1Zg58jwdysLWEdn1bfgXqZP
Kr6eswx2y5VyzAg/3EzL1d727efLL0AYZdSjnCM2JCHcWpeKkbLgIqzLljFbrmaHIiw9LHCPTcAi
qfw7zoijYj9ViR6qjZJePl9t2gu5E4kLO5fESYuJvaUgzm0xEwp6Umd9m01twwr6xD0iFEBKBKc7
dE9Ydb8VVWjAe5ll9MaCRVuoSQZZQrl21LEYdiDFJ9D5N9nJkPS5JY2p26gwtLQp5QV1fXdZF51M
qItiSuiurke2B6/IdSwZGb4cVM+GlbvdX4FT76ST7/b/5PlNkPrLU9M1bWjDwQ+IZXnlPdqZAX7R
4E+H2+A2LdMWk57eU9Mt8znwc2NtOHcGmacXhCvhcYrfUgHvo3D06K9cKmjYD1hhaS33UCHkDScc
vaW9+E8773mgYCOFAuu0v8+5YhVWvRxeWXY/IeI3EytQoXEylOhSu5kL7OjuYOFKYpserR9WCswM
kwPI0/PZfF80BgMFhKuRdUPk2G+e39QpSKHE7TOQw5NvXA3DeZklZ6l8dLBuMgd7cJerDxDX7/rE
POiZDVIk9o0B2GVQZ9Jw8vQtLqG3qkpTaYrs0avQTlkQFxZ4rj4iredyf+gL6nVaDT3/VSwyRAZj
akvPgeGVIYk9ej7bVzVYUQYuRDomoq0ts0BdVeYA26mE9YGfBJ+nOr5KDGYo+ARzgBB71FRCtd9E
86c8G/6ggFpYTVMzCA44/4vyRIBlOMJ/Hhb3yU+yHZiPQvks+wGIUj1EnCy3MFUEoEeAwYGVYd0v
jGAbCVD5QU/9/ZNnateN8GkFAaNLKlkb6NcUz+cDySpLpRaZwhuR65czgnEvubQfwkhjPPwWXOZw
vNqA3dEU4ceaPqdm/XNgY5GuOxsaw8V4RXgMIIu5nN0ov74p4AL58DNZXtcF2x9rer3/VDJbVewC
PfdcV9HBezuJ0yT/ANWwZp6XHi5DI1t9KwIHA6iVwRP3SFoMXOoFwBx9cE8aaWmlVT83L0pRMOks
4DPdayoKVzJ71s61y4Grx3R55uJbWdlC3MWzEKF7XWOJFZugTJIsQM3UW7seK6P3ce+O/hcSmEV7
Pjm8Rf87mXfUa4ze3m4UZU6YjJ831U0gBzUEApoSoKCHUGju7xli9Pl4uT0TSZCtfPfg44R6SwJD
cgLA24SAhGKYFErDiav7SSlHYMA71HNubMvJsZLeO4maVb6HwcNUl16eikK+XvVQKKfFq3RmuwYU
d3rDYT573dAGpKWaI3h9Urd6IBFN2QJpePyEHEjMbK05lJSCo3nGKcsqIEoQdA1Gnzeei+6iu67V
Hqkpy5qDdpiIMI0nnIKHIDe9ERpNpjF5YNXF+qQML83cRsrHHUVO69X0+pNVQ+K1+LQvYwYWTjFl
+Queahh3GauUGWs6DIPg9wFw4Tl7sAM5PR7HV+xE3K8mYeefGU+JWIGDEl/qtYtmWJddZGksvM0W
Cm5U2fuF1NWYkihwyWa3A5PPV8QzL8OjdOD9Gz31I/vKrTSY4Ro3jswehmXuIFHtq4SQkTUKYKn1
dPz1nwktJhPDOzqZ3TzWLBlMLWbKu38VXjMFzzOocNxmrbobmoi5f9dt+r8od6GF6RcGAx/UTQev
nNey9T9IiSJF+OFpczrLcVyyfYZznJvdpduysL2CF0hs4vCsHlx61HNgen9kWTK1XC9yElgKv/gq
xnkLrgZPB7ysI1wVu4sTH/G1obSwynk5UszbW3bnqrjPZMSZxImOYR09uKVUjK2KiF3OTS6+fH+t
ss+HtfWaBL3LAr0VT/3y++x/9N67mtgrZrJDM4o5AAPCI25HeNPoT8Nbb+kEhVQXSmJb1pv6QNca
mkHc38+fUdmLXqnGZ18Djdl89ovReOyj6VXOQce/lCnUSKWdEnEJCrn0A/jv+uZtgyon/m5546x4
Sw0hxaX/zXQxIegqb9nc/kDKGRcVWocdJZjxcriW8W4HlwsQCHcELGHna3QD+GRBNT1h8Mxiph4u
+GnUuxSM9cekO0qPIeMKU3qZw9rCl0Btlwch5hqUh6y+eyXLGWLQ5GBHn4VvflhCRKgQBGvQTdw2
iUA55fjS1SGPiVEI8IoRDzLVGst2y8PICzv+pTOlodlttPf5H5JrA56tiUZxw7Dk7dalUCTgfQDS
D2ahjYzPaB78+K4KWckHS6HtHAPqBwgi1qWUy57U2i5zeBc+KrPoRRtsEJdGtYg3C090icH8K2nU
SUlxMxfcQxW+YAI45D6d9LROYob/e8FTQh8oynRk9FEdW5tMdtYAB85NYDwlCtlxPwY6s9kTGRcd
qOgU44/+5fk91Bx1ASqy8O9ypOXTIJLlCABm+guKN/92A5kcVdGNNIzi/yajXHdnQ9hwIKdlQP2u
PNSMmYuqS/vtrUpnqhlP179l+JVtsyHrwLMHbKu1gA2PgFQDBK0EjvfMDMuLv8B7mGAsO9lnhxrn
xJI8GgTr2BqVrWU3IHi75ruyVgQ9Y7spUOeZ1WA7CUPrMt0blrOvB8dnHo9ZpY790cvzo8pOY8ze
j0oar3L15avdzDUhvQB8vshKJuhF1AahAOTyT+7JRfLP35WIb5xNaqCGROQnKvfyWOhcOQyajC6+
g486ydZszz5cUSOHJDIB+g90Jv6bkOVCYIyBSurecFtyNrN1xddSgzNKoTJV4CYilL8lviO8FXPS
iKZFJlOG5dyhaK6nwDG+cjeVhBY0XrZ88MfMknExOzT5fuRwQQ76YervF001XWsOI02cnMHRqZ2w
ZwnutRN0H5pSGC4dZHWbcFqL4HQXLZKyYVGT2d05ajxJpVcf4diw6+yh/DRwdjA2lKzskHZibZ0j
hYCWHPnsrEFnl169Am3mAcdJ7srhreo8VGhqfNpBSuf++GZwV5j09LnCjhMmIys6D2HbIdz43wrc
yQ1xiiCRV2mLVZu9pBS0JEkfVoIVmJAZKtUzG5PQAukSB+OSeJdTtU3wONAn6C/ncI4WqUMYuEXk
F8Wo/zvuCkEVUwQgZAHwTSj3c4YdCnug2OLwBKoFsVpchAyk1yPBfLbCfY/1I4lKfU7bcAklnGt/
vbPrQE6dmRK6tOq42EIgGbdbO2W5nVhQcUFRQTW5iXqDiLVZ42w9/zsuR/0jOoNY3+C/FOos3wlw
x/Fp0S6xbMs2Jx2Kh6CTKKHMv3CfApdzEwGNZy95/Y4RXOeHC9TbiBo2Fnn4cD7zYsG+fe3lFp4v
fLAzOSTi55pZkwOh2hRxcBVBOLpd5GJC9/R8sR0mDVFl2HB8PZg2F8EDpFW015MwcAE9eU0IeUWo
U8LO4xpr0owbXkrzo497+tE6lQ3LxbnuhtrNXn6RC4c+S+jewdltO9th5ZJgkg6Prbubg9ocucTY
hQTI+MRkHl46mm8c+QZ+aC/OGNDpOqHiKYoBBIaxTe+GNlRvbWYIZQCbyR5ZD4KydBxUt99DXbdu
8GpioHfKM/4PAGH+RNK5SSUNUIDoMh88qZrL1Ma1z2jLS0UMgdAN/FYt4rK0srDa/TuuUple86zC
60ltFoYVxg6gm7fus1glBP4IktICyD62ZMA69ajHNCHi8X1Dg3bUXYUKiJHFa4hz1zmBSCY4GYIR
afClWeRBFamAjBC8hmr4E9QjHTYuU0p2I7TuvL+Oa8FREBOxvmLhg6BBv43Oq3KVDRlsQRnwyCby
kT9i25a0/SpiSdmdcNHj5Ul0gT/4AY81w/VPN8V7exr7kRYmLYfAFLLnwMOTKQWZsK0poyub67UI
oPvtXlVXyZcGKf8spEfBIsKiGTAYBsxtT+AIQa9TM0yRa5oULUAFw4NTS0lXNIvusNxsvKhZsuZX
h12/+BVdGddEKGvjWTTrUbjPFLhqq4nS/ftpb7JF3lhmtHPdPLWaZjf8DbdMx7zWjDmsy327Okel
mlb6zRoAvELcNhDBzO8TUKqKR4fq+lxtdx4mxIwlgP5mKm7nd9jqu25a8SBkhsof+fpCp5oKHRgV
PF+FZfC5qVXVkbzSHXkRAKMw8wkfXB+nrNCHfRWvRtcPYM8hGbfxE4+w7rZBfQ8C6Bl3sBq2qTtj
fUpH4AiXzjGcOxViRfS1LYKoRhyXvaZfXscGu4JajZQxF4OrUQHatiK2wppRmklt2MjGiiFekXSy
2RU1k7Z7I3ZwGobhG7qENCBgxVqH9hqhOWMUDm7W/vSZwrMp+OhJ0ywapBApPOf/4sibyck9sh+8
r71Gv34BasvKEpa4FjFXmQ1Ls9FALyUYy0bkub8xzYXR+sUDzfVhnUyViX7tZIio4Bduo9GxZ5kc
grRBfInsdjSgUv6CgQvI4i7AoaNlYmIfAn9B2rhvWDItnSSrxGYPAPX+aWM7oYmoOwDH2Nb8H3QV
ncARZ7VY42GaxC6DBPAfdDwmgDVdmn7XmJ9btjZZfXbM6M6NY3AovbBf0OJzmDlweSFA4wj4M6jO
YxBRi55jTGO8oBwzlVCp9cKRX7VGCjk33slpIir5qCQVjjPdv1Mp0OhR6Qcs73M8a6XCWLjzOV2s
ZRY00aMOtwnfWgXGsZvbKKKdxw7ZPa96BOjhc7LtzP4WVSGhDqXDrPjmF4TueI4V322xYt9TzYG5
epKyy0J8YydDTMiYhRaeH3nhYuIW3v4P5tftIknA1eY2cTEAAjrw81pIc4VCRhycW6QJFOOxu1xs
AK5RMfI+4gEDTmxrqlaISAFFaAPKRj0zRPpR+v2O8CsS9ZYpmkbmrlr86/4aAivZHONl9ixVX9L2
l0wMTwPk2RmxcbM1mJ1ozIHNrG8MHwQ7fxtukjqLOR7jdvhTZULDP7QioG/m2RC43JcrumpEnNQQ
uRPrYa8ZUW9+RCYBC7CCIVoqk5DQXPP1fwIlBKv89MHJmRcttth29Tg3u/IoS72cLT4YYTxbpHFc
bk6QpuvlpqqPKKVSjJf8Jebq2QqNLaHIFvreo8DDyhune4jB1NWh93CA5KRv6lc/n7f+fqSVMu9t
7nFCMs8x07fVQd4M93ePdiwX+aBHHxxN40OfEDh5ZBEVHf+q3uoCtwIlGQLh3uVFLdGX0/xoDNZe
8ClxCTG4RlInwenVe+b4geoPP1YoV51GgW/VCwaUSI+9zvyu9O+S/qWW6/z2pJCRZZ7LvriMtqFc
qBjNrQlGIqcV8FdB5RgmeEPQyZfOp7pyAr6cE1cIIZP1K1seD4tKqp2ndYABEQcnM4j29w0pJN2d
qyDruGs44TCaRKKfVvZlQxnsK9OyiArCOqt6Ym0mxuY7jQODD+WCOVhrrY3XotwlaYFNcOQV7FV3
f/gvHT0b3TOyyYbCJMCECfoIXRL/z1hFCQWS+BBvBZEFm3LPiTHlF8WnFtCeK9CQTITNwbZoyGgX
ldhhEkVlI19Bfur0Z4o0D6gyqFoNGCpJksPCKF8EUXwVPn1pga5BG4RMg/4EcxoSDeoSrjK1Cf9d
h3KTWmlMDSrFDGEOludtr89ahzt39iTm5eX8nk1jRbNTwO+nLUL9A2k7dElp84yH72hFPWd8nc9v
adP/uEFFQG00R2MgeTVUTau3krP2CD1dcYupS7ZEKdvUDKgxF5lykvuIIu3GzVeVtvFvCOA2s/95
ZnAILCRrA+mJEM0yHgtMOWZ0w92SaqkHX3Sjm38k+uZl6AS8r86aK85uMIhwv+/maAyagyAO7BW6
c7ICQzVJHU1JnhnbTgGAHtwCJxjgyiKdhyKJBOd6+UbFACJqRsetSpYe0dOeU+hZpw/HTsm9+T1j
Qwe7Gr29nmmZVsS/ivDCLd7PA6z+6sVVAhHlzvSkhP2G0E2IBZShgYZRt+7q/DE9wppOWn6emDcn
sNjwQRIiy/H7/1c/yh7tMsPzguS9IvUnr9kW7I3vPNbWZDHSVJHhx9BRBFQDjU2ZOrcOLlb2OZx3
ldjg0KUwC1VFxZciDPpPFpGOqrDyat+dtqKbPLWDuKLN1D93EHrzRKNheAMf2m0eVe9k98YulNv7
9IbSJi3+M91wSPQKgjFHcqtiZ7RF2EYSLNRhoZ2YV9YNg454tx8fcx0Jl5YIhNFQBWhhjHAjFKdL
XFlWbpw1GA8PaaPqzywtZE4CRoy84CFMA/vkYUuRco+3AF/dimnbqkCmNKpdRedaRY6DqmtQKXAl
SERZAJoIZnRCzTYM5+vmfEtbn6zs4e1AkyWe7WzdQKOTqy3uBZfK7fl0nesE1CfCrUJegy74brWv
xNLbeNmc56KemkCinmB6Ip6ApAbc4kZ9PujXhQvk6IRtjI024WxduWeIsQQhM4EllwhRaOn4kjcZ
GPKJJ6OyJ5FiX5Yq8mgHzbMybqFeXf/FY6iicWz0I9/BYtPg2emSiZI+cQ+l5LXDzyZ8ZrgoDnst
yuPLmDlMrZUIQbfonloBU8VQ8PxcrtdEwr7PI9JQwnHN/PAR2x6mOysax8UDGOR5ZRwY0NzMAx68
y2smqnglZUkT88+XckkWpsLM83KbHpUiZ9V+UyjR1Uxb6I3/H/oW7t/EmqTAVn8MXb2KYcAuICua
/+/sPrOpr1EDW0SrQiDEp/5uKmcrqK+iuc5HikkZVzUYHYlGiLXMdMwEK1/zYlrF7D9iLWo6Nktx
1F6gcsZuZ//R4VruZzv25VLRq/IezDOSp6X537pFIuSupCiTCfh9RBVj5mPqQpvv/a67Vz6AZNve
LD0VVCXwQskzi1ZTX+7BauP0XhEaOobw4Nl18TD07CQZC6GmVdRGxrK1Ge5QlcEgq3a4gM4NiNNU
FiT2bl/0dDrGrN1Lp7Zzuk18rV38cfUsq5zWdIO+AeF8HgBS3jhDaQDYlVkI8MKvryz2KeW6gk42
MC2oTxKDYpADbGXVb16teQdGTdPOPztIwMNVurlFltnYmPqKFiUOc1/ccPE30q7oNgIMzJy6cA5f
lVhgyVPXVfL8NvzsTtT/zTl7IQlgwhZtdDk8zlGMH6Htz6JF4GS2UMGMRVkGfGFmgNdOsiT1q964
GxPQZkUplWqelsv7sqi0eR/fMidVtgja3+ALfOjJeu/nepaUgcI52V9vuJOBzmViZjcipXJp9i1y
QzppEsX43eF9UEe/v4N7BZkg+7SJZzCAey+1O+kYPzpWeRxkJ0DiBetF8swJZS9MsCpgcNgTB6jw
srVnB5C8iraYrdH33V7vY1YbJ6uHIxPEXD4Eh5zQ08csVzQstmZB/PeaClpO714TXpX1sewXGD6O
oIbtXWDzrgi8uVS/AZM85DFm2Ex2HDxQEx9Y3+b+9irP5bu75Qthlz17xBdsMaCCv9lm/nQMfV7V
z2yaRmpGMjcXFWC/q5zD7x+HtsXhNBsymqOGCedvJaPokY14dX8DAiKKNRtgXSdD2h4v+ul6Ukei
oPbAbtX1+PGz/9/sAXflLUlmFisZzozdKlmrPEDzhIh/JaqOlFIxGAXPQ7QIHLKUuboYFtr+gJ1N
CxURKC9xotQ4sSk/lmGmO8u6HHqgSWnLAtQxhQy7hadgt9SLOaop1gPOvWV2eIRzShOUrMbstLm7
5LpIp3QiQ58FEuOuU1FPNBy79lIBxI7EMY6ZTvQnaEQUrbP92YmL20CuBC/U8/uAfPDIpsKneple
YAmU53lu30pLrGO3EfR0cVTgeNgL22eaLJDLVh4Zo/7nMZEcU3OpfBXMNe0vqaWOKVl4u9ULjdt4
HXEE1TtEaZ6IvPUEmIwdxED5HElw6XTKLGitG66geeiRPMO+sy4J55+TD/ZDI2+/TV2WEAWhrXeq
Nx6jKjYBO88icGyO5xcab0kTPjmuqGLnAs2+S5LMTHcov/h8iXRhWn1jlKV8TujWK07V/hdqHceC
ZbdVEniBSIcgLsY+Z8+ciTsrj/fQTzKOwIlqKBxBAqty87/QMlEhfPUfsH4W3LHUY7dYSmr4CUdd
twaFWATca0iIUgw8EMO29iPF8lsEy+RBvAlRPAB+4FDXc4ugK+4j8nuXwU6cSLE5j1DsDIZB8mrc
xZfi6INQhtyCE9UB3uANkz5yAJ9ObLduv2nIWZ/XrimMv/WX2rOzKYLmI0TV6y/820EkKsw4l3JR
dI4tFfEMP/o439GRCPaXDLFcYkhEDpQe6xfWWQAKKSl+mNS8nIVWYza6BAYxq+vhg4Ztc/LO6RpT
IPhq3FSBWYh8X4oNlEnHVkWdIjlPgKF/qUGrtW+4o+JKQ8AWNp3oZ8ziqSNLexoRs4EOeCKBZX6r
KSkaDfdoJ6jRnVuOJMs3DZVwo0+fBdFOAhV0053fXHDCN9RpCXVRsOjub+D420AiBrlSg61oKBAb
vIt/EtW6U95DERY1UXbWYA3byX2QuHiPACbYGa3DTsnn253O+hZ+S4bQ6inpPGAJ3HsBysrZ2sbh
bPXy1Y/az97WcHaBdboUryXNPxI+YN0xfnRPo9NpASGu80wscAdT4um08BduxZ3eAwzny35QekBY
JBq39ysHU3KIUagVslahgZ0IwTpvZinc9dLMTRbr85VJVPy9WTEJ4G42S6YgYMPjKq8TAPdVvpIp
UaqcHlzlSb+9EtCunsUSbLTNUSzRmlG+NPxr2PlXLxPY1OdG4ReL1DH0L7+5/4iMDOkL3abxja9T
sByQJPktOPK+ABdEFMHOPxRMqioRj1KmyJRNiOjofGmUzSR7J5/z/W6GXIa9kG5bi6gvQ58cRS0z
NS1z8ZWYcdXb6KWBnm3RvZdb5Kyqios9gB64vF3DH0qw7AfFHmIh5yFdNkhcOq5dN2lDA88hEh/Q
rYP6p54KRJlEAG+nc4CRYDeRLyjWNV6t/SFjgX0GXW3C/SKcZMWgqPkfLB2PYVAZoLClfbFNku1p
q59TWNmFawmS/fFu/b1ftnzrRbCc3BqJF5D6f3LkIHJy9Sv7DfYElfkeqBjIeZmJLz2WTouih0GU
wldkW7iT+e4Ck5QWqWsxBKQmubNQD76p1dnj5N+H4jEYIDie49s6R6HhUQIkPm588CqybuaKuGUb
5vKyGN7/xP7OafC/I3tWkpK4/NMfAnmBg88A4x6cMANl+vpZtTbM7pbXtPRE8MNnVw+vyI/xvMrw
jhlzjYGGaoh/aqaWdiQYJia9KP9dV2oyUxyQTD1nJRi0UDJKqa3Iw0gypZvz+Op3qgXAWFV0ktBO
j9SYBvWYXi15hO5SejruuxUud9/EUxIo/KK9XNZcKB6zH4H9+Bu3PnXLeFZc81AtYDvM0ny9Uv39
3BkAbm9+yBb15WLU+2a681j7SDX3P4jHewMdYQjq1lh56FG158efayJXLAWQSIJCP+HIYMzxMs+D
s3ibNhfWvpDP8es32s4/t/lI2Gw+4m/pePFYv+j9gqDp4L2m4LsV9r+BcDgT2mfZL4nR7xXG6Mnn
NgGPLwGYMXZAsRPkaW+zpDwIn8gIrAiC/I0Bj6eRXco9K41W1pmK1Ww7/gHLrXICmv34YpL1RfQc
lVS8VfrR2wcyfkLjm/gx8CyOrgGq8PS6pYRiScztOpOfeXCs4nohDhUZ5MBoH9dWXCGbgr+Anyxo
69Q0kdEyJFWkWCcmDUQsGGAH4vbDNf1heLivRnQu1wgmX7qigtcyKQVgAg6Fq6nOpiuNckO1L5FP
zPLcBn5ulMydc4PfAarB77vw8oPuxCYWf5DoVYh8MT8HclxH74v3nfklwG/otV8mAOP36CIpHdXa
8EOHVPFeqzoeo51Kw16VgzIlOQMvfoZEJXjOPf3xjdMROTf4/tMVxBnmEhjat9GHEkJyXfLnrx4m
tZ7lUdE+NhBM6OZjquRBIhXfa72iys2IpJ9PD1E21AnaoiMAnNjLPD49S0zhyexz2UoyaHuAL928
o3V6dzC1+ZgJgS3rmWIdff5LIx1+cxsFbdbOH3EDiGGPqySmds5L7UtOrDs+DkKJ1dtQSxbzDMWS
2x/sR5CPEeVFn3cBMNHA8oalmZfRt9wEjS5LhXf9aQ+29WjSjL/ZXGVd5xA6RSP23Lh5BVAxmMPT
3zJF6urE5IPeyi4IJgf1in+2CsErTR18v+gdvDJyJ2/+j/ixve7Kce+JvYz6S1VDoEQqNG3mEnT3
PFG6906dI/y/VqwaDRuC/AJsN3eAh4E/GYv3i0t9iLsqeYRh018vYV/2X0C//q9rQHpdJHiWqZz0
BUNlJC2Rki95bLPAxVj/q9W8U4OLzKSNK9EZ4HkTn2CYuew3Y3GMRAd3nGWc7QYOK3GCPoxUQlNr
lqVa9PZ4dW5tMSux16K3Rz8OD855dNcfm3C5Y2IE59Rw9C9e39OUqKdt47anZ2QkeMh3KkvAYekh
efZ/NLG/u8pKUncgJn6VZOv7VecZBJpzdy1XtDLoIBg1v+Xep/31NKgIDlYzALGDxlZy7sqEGlPv
a2Pm6cEAknP5TEzBue8zBPR3rUQP9sSMN8yapvoFrUDYhxNybhHvYoAKdNX+wPdfZL1f0eSwgm+r
oB+DwL9QIcVuqeU0K72813oLIhpsUBDSBGUdnQKpIADmYjhPrJcnozqR5HXzSH1GfzfJJ9cvnFXr
wmEFJ6+c8g9vSjiGRUtqpzOMKPvdAvVV2/PocLqEe0EwQFdUnZPAGBZZgosnTIp9K8dOn07KhW+J
g4NqHdjEHCtFaJCuQkWpRk8ss21x8PfGIQFdDdJ/uFHRQMzibrbFYcpjuuGrqTqOOvjSDdO0Iiv6
1FL0RPYROAErq5Y+oDZQd5Q6QqT9AERzb0f9YiWfOcNwmQ/A5tilspzwVpLGqYKvw3J65f+W9pHE
V9ePaPNdTZkwVg7ZFc6BAmOD9VrtsDP4O5hD7p3LsWl8xS8E8qoaaponI4e1GMvcrJtlmiF8n5wl
hFc6OQMSNz+AUWb4kTVa+8FHz5fFdq9AqZE/70gAEsDZfSk+XsW8k7Hqq7Y8Cjrtv09ltcvgAyrn
YbHERRn+XJFRjM8GxNsbdyrNijFMkcqwZWQqNOH/RjBxXK/BV2a/NINB3hspA5tNb8DxZ3GiVYCr
+deRF8xKGz2ZSUYUOqX6SkuiLnh7S0hJN7rzWDuWBotTCpCtpwc10SOM0ds9O/gr2ZUkH2R1RU6I
nvjz5RGgOTYtdgnv6WQrqvPyS5zy+jSjv+wkxXxgPT5CFwd4HhLUBsHUKeGg0ZKtplK1GPOKo7Wj
b5QrxGzTUEfkaxqxGxiG5FIsbucWSEsnknBWqeh8ysKEXmWJB6PkRCsPdwrb43f2JSaj0ZxwGlSJ
yXUGHjl8jo4Xj3ogopP3Ec8iF0CWSm3WBlzxm1ztRPpH88i+9aAG2Xd620I8uJzZFIUugr0OvM5q
XFa4SwxAo2Jg/HZz9Vj0BCt2OVjT7aJiD+82sccEQ9x6UFoTQKHzT4WGbgjVDu06zEM4NxDgNGrz
9f5uUKAJg2CWYHT5FDFRsx/7oCvfNkK3hmlMMAJZGU4QcazmOwcx4KxJrNlfHFwgSp7QjV0lVSPN
c01XOKNXUjY7Xo/JTco2kxiNCilfaToobSDeGuUCh5ronyWlH0EwOOZ/X0AjaTC826U+IcttgCrE
GsOxug4xzX+sb2MNwtJDeicHQ3uc34pIgWkqBQlzReTtfaNiEddIut6XxFRNsY3ZfzccJ0PaCNpq
TQcPCSlQN3EPO1RRBjRD9xqkOLGJrdM2mNBqMNIGYMnNRGihDyIPdgB/RVsidFTtE5TahKWHxHwf
XD98qTMgi4skBlRDcJYGMU4Ab+EOxYu1Pg4nl9AbwYwFNhHyD1dpoogl5fX5h0UmuR09UE5bpCdl
7n/wRHGfj1Pez5gcbSWqtCIiYOhaZwVQ14f5BCNrYEQM7KgdfU8LtFO0jhJB9QzBXOAxTM5c2onY
9dDCqTSHSXukHiniDmM6vKZLZ2w7o03o70RMIc0Q5YP6IeJWg/gBpuqfEaDFedgb1yeDBITcP+f0
hKdoOPvwmCdK9VkyWUTtzPzb3iqjukDqmAGJZIn9MOpIe510GhPpAQd0WkSplNx/T0X4CuX/UXnq
md/2U1KcMjwpMDgXCPuv1GBs87PIXCOGPshsZCb+nrYgc78PGIbPOe3rqTVwQBtMCXmvfmUaTXWj
iLBDnWuMaW5wtadVlEqE8r1J1osRRIJLLb4okU0oPCypkqM0k4EP2ft1KT1K7sSSSp0h6SFVBCBS
Nkf2brKacAnbQdj9SmKD+mncyLuWbkhUvB02y/14fdU4Es/AVMT0BuUU9mJYlnohH8x93SjXhO8f
bkfmrEcVf3DgmJ3++yAiJAOcWc+GRoBU5Btex+lbuhEmvSsrCwa+luAwGrLe7bp2fqTnu3YGpqc7
3N4MZ4yqC6If2zX3fPs4VnCiEbjj8xSanhzZpIwLu688ZzvZOTr9r4ixuwDMUTBYzoJh4ZQJqh0T
yI8/JsgyjgTTHDriKl9dwo7ZQm+BrUx1z82Gw5M4DEo5LelxCjjeIiBe60/sjRlJhZaO7wScVTnz
tZFd9Eq1fcQpyx2noM29f6LPbHMM3MWPuVCZbpY0IPIQtRy5Y4j9yUwMZPF8p3TYC9pwD8B/waWG
CbOpH1cMde/4DxvTGE+ZxhPdsxh1yDu2hEBol1PKjMUvr0lKDpno0i5eNl3C3cFx3bJZ2G4Tn1c8
/sQo+BsBZgkYWM4fJeT0R1KQ8PSZkzIma1JC8O2wsEGrXoi+ipHJ1d4o0plQzE+5zIm3Y+Xlqqxv
7d0F6xuJRf51MP3cQhi+D/JZCsLCXdf6qcWHewyQoN9knUp29ut6q9Jw+1u4gni5Or54QOO/PDYP
/GzeXe/f3Cqj9FMqePuQ3dqe6R+YiBXiUkun2qOvy5KZUP2hvp4t9xCuJGI+FKBGS4kT9vzpCWyj
bxNxekBTn85FtsiSBEoHlghHh/ileMJ3fMfXQBeMA5zkNKJESXXGMsAn+0Asgktnwx6upTLtiMFr
KZSG5m+8YyOfl8tevUZJfH4/KEb3ZH6Lu+mSP3DxbhuzZpbg6EW+ygavwrySDfTVSAYJ5vKvsL/2
UDjKb38otJF2kMa2IUB6bzOc9SguKLYZoG2XWRQWndq3KXQnvt1tVnFQIOmbIC7QDJvax+nNv1Se
uyQGvEwILWEarqqONJYf+2ZWAfVpnn/8ajdtB7/ql92DH9NnZYiHtRZsRtU9WcgaFXnMptPLOF8W
Qrgt92HM6IDDhYgaTH5re48YRogYWJc8+8rJfwsVlyQzVIEzdNnOkuAy8xDW/20SYdmbr/94MUDD
3SGFgCHeJVNpMAADhVHx8gIKohs07FkgpZUDBszPGZROmIU3nek0E7+T1a6YKS8Fd7vHz76C23Co
T55Msu/DJ2aihWv8Pq5O01o6kjrmRL6i0a+X45w8jITsViEvWtSHxGTk1IPIrG6l1vc4jPIBJUBO
dpw5fPFOC0P4iPT3jFe442wIggxyJnK1AM+bm7J4ZiFueiBLgKWxRVJZrlMV79OLeYqzb0qgxw9W
0uvRex0TDFmB96J6fUDi6yqk0VMnLJTg+DQ0rOu5BTGA6d8lgPb+zlYuJDUuFti5cd5UwLkifNtT
G2GvEjQUZrT4mPt8q/27yIa+8nwpiNnyv7y32gxXdTOXjV2GJ+YIUKPux3pFMb90gk509KTA6lvT
xco16BoXSbMkTn06PvC/LIghcflJW9CS9h3+yezYi0YVyL+1Hsh0wBILLwDrMmXkPNMn+gkKXcKU
M7bdyxx/E56EwOiSWViokPvJUAjtRlAuQRvp8CM2aFf1TCzJXB8NWWsgrkUvUG+dACkTyLz90IGN
bp5kriZfjhDwz6P5u+2Wy00R8pOreVaBeU1eq0jKbccQdRwzgHMhkX9geheS37hA/2w7imHvqYaE
uhtWggqo6L3lAp/3cPyXXSe/dYLsZuWki1p0avkGQIPEXE5MItPskqzOdUprwJSXl1FlLEk5oLDW
5e1qfAEttejZiHkS6XljhKrYqXlZ1tYx2MnBFuKSmESFoj9XPT4Z/oUBHtUuhCP+5SLQO6GVXNPJ
XXAvhFAFZUJVH0O3JqvX/ikNvMbbo2IVmi/3C7XnjEPw5jxlUcbGyPl469rN3ML43QIwXhP7ZAoJ
zbebdbL16DMWprKLYr+U0Ib+K5555KOSUBEogNb77Mf7Rf4liI7y/pfjadRekKlU+4CK9LFBZyyP
OjgsuLuvIrVb6KQVAHyckVQzduvS6cflAOZ8iNLb036t1mEQXgXagnPozvJweUTD7Q6O25Vmow5E
2qyDZBuYwnjweCZcNmxmwvx4Xtki9uRU36UyhDZ9er4/J+XEL4dA3d+kolW+xSAPnwxNnfChLZgm
ILJkBqhNBuR5zdmTFYVLhm5kh8H1cbGE/6mQg0vRCEqoSI3fBDVuCDZgWvYcSsb9WHViMPnajOCw
tknmX7Qn62x/KGJgKWBMUF8OPxQAJ6ydpDJGsiFB1Nox6nt3t9IOUD2Kj5PIoKU9GewqR3fZcvsJ
XsYfQDQ4vy2085t3e6NPmmzHFXrziSIpVdXtSDa9nyL9G1uYrH0fk2iDwmD1T0f1qYGDEHarDh3Y
xhiJ9PjntzL5zPOYf1k4x/sRsgeOz0/ZeFPUwzVOCh3YE/bl1jEp4few0EAy2SvyJ1Ir4uJPYSAG
qRpjRfMXogT4HuQYcFCz1E8oO5P/c0Cg69b6dge70InscxWfyEeSh1DWYSEQ1niTHjKA9psbpgFm
3NY29yFx78NIkNvFfV27XrBSgUiVNdQghQYAcJyJngWXLHfMSE3Q8+xJL5iWTY0b5gLwG0cDvlfJ
4c0lRRRV2ziBatKRQE6IxxVn/AeoZI4p+7piDIiNdjWwqWbcQUsa8RHWnOY8/loyKHlIhgvxIwfn
9Bcyhx4fydC1SIubhECWvw97x5voLNqBz1Meow9wtbG31EiH9l11znkxXMrg701zvbwpLy2sl1rt
F2y6uv9ASbY4fA3nysZRTTtapbw85X8B2EhaSqssZurLlXrdzjREjBww17sZfKx0iUF+p8WMZ9MF
wtgO/ncx/zXV6ziqK0xH4Y2uB8G5C3r40OcXwFQ7yur4+IcZu4YAI6ldoJRTzkFGXjnIkH+7goKs
aj2NiE7cS/0tdOSOjyvVHDwu84xhZwT91R5v0NlBvb4wNQ8XatOLSHW52Jl31dkpoou0p8wUH676
TNNV5TFegPl90QvedEjsH16kG/DuW93ZhNdv6dW/GI9xD+a9KO0vLd1yVm3DlVMTglC2URx2XkYz
naeer/bp2ep0tuRdwb6VPohYPLQZYCQV4rBJgVZiEIYUIEPFsO1XLurnuONpT0MjZ8+tUfsUGu2D
KLAbjUcTgB0GskqQVCbyhPtmXIhRnWcV0gkAFxggwxwCLs98PiQfvXuJhc4Lti6qosNaN3XQzlq9
B9Wtkvie6sJ9cOMSkOn1k8cy809AxXs+3t6+uC4X4eSKKc2wzfrhJIO5gm9xaDSwFsX2iOX0XUpj
KEG1rVZo8CVuiBtCZcqYGUAKLqVpmjltlLkT9M8Xt0/5GaNOlDgHLo9vckyhttr+6rC7uN4oxUNk
1DPJ4z6zGvTROqi0a2p5NrsXvgUj6nTPDQFnbOsygVB8jwVm3dWnh34MBkP6/8udD1fwXhvlvOjO
ZgeABuorFF/UYJIuzELcgy5UKkNa2ltN1K0U6U/R6UCLa7ZapodofaHqnJ8/Nhvqxn44ZPh5ewqI
c5uvAuMzZM4Gg0ZYJgUH4R9b10MRLbzQNUBIJ8TEXWnDLpb48d6oOjOu7jhB7U49t0UYKaiK87j+
5+bsFWs7MkYtr0Zhl1QQC7LUFriFolSCp2GyaPhgwrsdZeHOa9zvvwaw+/QX9GKxBFC5P/fs0LY4
I7oS/FpTm5Ih9bbJqpEh3q7KGj1IdJc0e05bN/3vuPqXeP6JatV64Yeq2cs4cZ/Rpq4RGZAivAIp
rUF3WhssX9Bakc/cP5Muh5pbmM3ktQBjSlmhC0fa5HOTiuSYBFfnB6Z8REESnUqbvB+EQ9PBr+8V
PzbPEPXJp+t0fMaddTkvS7cuoYfnRTnNj8rhmloz4XYoENUq2QNfY6dJ1BFrO9YqmlephVNMc7tN
WDD9ys29afvXwXnLOBqUCNKaU7V0ubmMAbode3XLohe6NjyeXKUNVNsM463hj3xShmSx7yWUEp24
s3PBid3EaWbhJy4TTqo40dDmcuzO3S2zBxmGNenUBWFk+l6NiLSVsF1PmXDCJlhbFHTcxA3KfQHd
m2NFSq4ytMU3dtglLCv+bWttU1MRRJYwFZeTv7f9+oRPHEm+EUhYJ6po4fz56mfc1tZ070Q68hLk
JnPgnfTQu8TIEaaLaXZRFM7SHAsRj5vpVBJtL6w6gYZ+9Wv1u1rsufEYhc6Ft3rUg102SANIpKTB
D9kRfB0TKK2OnoeGnW0IQAybB6QhKOABg3mH1u8tli/HDfH3SoCwdDw3ICNmn9rP7456P49U1ROA
mBRplipuoKIa7lGVCryHZZDcIslcX8ui99Tx2ipX+KapHa1dm2j1dB+hSZWCkzoK1xPQNtL5lUqk
fIlxyLuDEVmrr0tdwerp7oKjrkZ9A39GMrJuzEhhWVNufacv3r7Iz8xM93/97bDvsbsddpUb/AtT
+b84VPOLlVTvpjeHUJn0gehj9ViJI6MwaQoHzTxNho8X33dOQOzf7TrTzOkqaxrAe3IEWcOcbUzz
HIS2YNDnayQ7uA3k0a5DFz+QiSOZlCMs9Rr5hd6HRo/bWOWarJxBgPJ77RsfABsp5l/HOwHPvelN
ess+1eDGPdg0Dp65LrVzalWNiB2EKDjWXjiUEGyQG9WAjTW12ISZTEaPYMnG5MvYJ8pHM3sX1z+C
I56KTGG0rruSxNoj7YuNvwnpW1K9IPipdfZhvtOAFiWHZtua8f04sLqNCDt/jcC5wnsPbikjydUE
wbCYOumDZL9Cy/SAJysEHq+1AihJ0hHLPrSVVrLGJ7GFqh0oKQswnu+vHXxAZz5UeJ16cuSUZraH
tOEAzC2qurPkTlKOLwHoufH4vi1mXBTKkJXzxKWY8dpCI8Mf3RF+m9JTWvDFhMOlO7zXhwCDaONL
Kubsv7d/qtdFNaXvTLBku9LvLWsKfxRObwIAxy98wF7uKrCQvn1rdgFbRkRkXBrl/jyX7cmHwQM8
V6mmhLKlbsMl+oF1K+BzGXYANc+/uz9CvM0EtVMyDCoZIjPYsClkNcdvZc+5O86C4Z2k8mv2gFaX
fRP7zCgPp4I6v5jYo8jTIvH3ht75oHPARSZ+Y8Tc3qPHIRLWf9oM1yDLgMusxsud+Si1HDaHOB3M
adp07wnNl78+zwuTVQOJENq6XbBg78HDtk4WRrm8toLm/YJK8LLUi5kVeBTvrOiaoLKkyBjWEtrX
4XY+3hFBvCN9oTUHThthZqsLl1rn455hwXhQ/ag1awqhhe9OQmXgQtAZESkCapOJyUH3mVbV0p1h
BoE8pVM1YFZJ7VjLm6QkPcHATrRIJBxgVNgzEuFq0bhssF62wdtFwgTjQ82BwuAwdg0Ctjc3GPJu
RkEfZcqhvC0zOa01e4Xz7qPMQ2PV3q/VkzxCdfLCSdDvQ4Y6bH0XjyqZrmpVToVNE3Ye9OZbmwrQ
CbYS3ZAoT3NM+69CbKl84Vti91ZOJE/WczMrIKTyhK8SBCf9y8jwq4jdhRIvukM5FzoOC3dMt3I6
1tg2+4L48fEtEhvUH0g9YzQKlmhK9nzp7TzxQTwzM23aq3IijOXu+TAHpyAE1oKUR6dL7rGDEnz6
0QpCsG3NY7OparKSRNnRqNiMUFPjsAhd/DWLcsCAMeyi7E3Pp+zmSELbXETY8TLxAHc/Nz64nCTW
y41D6O3wBV+YrCPQuaLi7GNBQke9yVPR0CtAaAI3SGskKiAWUEhaw5iP5wb+dYLPpkRmbldUb2iI
eLk0mTmnmhvK4CMAij8xz25LxvG+eawjtwEBASm5EoUg3lSZXRdi22srITVntFs6/yJBDEGkpUcO
TmO8N+yyldnoawDr+JUpwoQLqtirqDTCJyTJlvNpyRxApwHDLSTYswW6uArAqv8fN8yP5LhRYatc
fcwCIN90Ce9CxDFtPSm7/c4L40U+2Tqa6Ps2F8wpTH1TrqBsdUneYIrafBUZoOjU7O6rOaMFnWIA
hZZGKfICfBuzQU98i68g2N16Tjol/OI0jZW+eB/CEcVr4eb807CjtmnVMutrKe80obV9BdeW9TUo
RfCer6WgMp3fAwmbEdKz5+iWV50K0b/M9jIf1iHfpEWPX/WcPpliqlaZm4CxJj98QwcHJkxv3fDK
pVR7gHfrVhsb4hEoYLikZYZZWMV1GO1+6iXkPcuMKRGTqHKRfSiddqbd/MRD95zwzUW/YF4EZUst
whM3f0SQNf5HI/0SmvcaHJJfsU4OHPF888l8ejrIkwqq8PKEsxsIOpqThqYeLoUkJSltvJm0wdyA
Bf4dD5biGUSfOFaEYQhJPp3wCrV/+Z9xJFWmsCyMb3yH8ERDsu1IDITqHuaZwtqouKs0XRjO4WyW
+zxT38f1TnbkGOl5rHDoRDSSoImSWfjnDs/svw624gvPKwtHO3isV8MyhbEM0cAKA6X2ci/DPDOx
QgBn2mBGt4n8EnWshYYKUOjIf1jxdtc3CBd70Qi1luhN9WFQX253Vss6HTt6EDDiPf6DzAe0BcaM
uRJnuY5ESAbMWlrbpT7f3Mv1ckldPcsnsE7f7GcfelE1cJm0NPODdOcPyJSfNQrUhx+qdQIyC+sp
hPwbaKR4Z39DiyiZI44v8EK2f1F+UURu+GKatCAUToXBXetQMLp4Mus2FwtSRvJNNVGcJwSZw7oq
jBS5lgTy6Et9H1g5cuisdJ03GIJX+C1u/xhfP8hpauedeLtG55/34mAasIO8Hv2kkwMmFzQttVm8
zlO9Fph1vFQsLguEK+o2LhxtxHyUknj1WoRiSStXS0ItG8BgQI6guUQ1ecV9Wur2FAnT4wTuN/t+
mkfhAiqNq4UQNjWuxlhHrKWmpvDok6mE5fk/uw+bNbbd0wO5Ii946vJbIGOuwnUcEkdX+Z36Wr8p
o7/SmrJwFNkOY4xJhjZlW68W5KtS6LU13hdZq1vBMoPfxKVowEBld/tcg0OCOBPxUHjhxtxU/evR
EY4ggRVymLWdFIVDvUT9BOHn51KTwnrCCFVpxlHV6p/D2jIElDOW2Wy8QngQUjEi5R7LGY+VCRDe
vSsWR0Q+teoQuNEFVRcTJoHX2r/8A5XamEaBAGBMpmadmADdLVuhYwyERJwGCH2x/IQaugyX00jN
KBfvnTLCzCgqoZTfi3uJ0+A7YgUYfj+I5fZoS6Nv+lUlZ575TdZLh4+lyuUhMwD/KWDOMQnKc867
+y8W8r1IybwA7T7uoLBGl6IXVp8pL+Bugkg5/6lsK/336phAuJOxwQxf+PpjlvICD60T+wBZj/F6
Q1Gee1eUuMUEZ5SP1gWqpDt0NgL5BnmI3RneKvT792vfRYd5mqnkIc/dAWYtN5pgdEBDkA+0173S
EuBnN+tH1HKervDQbNKcxFtZx3Wl0PK8wZ8ly3KIKcoptfxSv8VQOHsrkSSlm6S0gvpV+nzk7jmP
dxf7yqb5DOnQEVTqUbyJLG/plQEZXg5/XlQh2UVhjAjZqs3lPvbssfcuteFek17cA3pxFqQo6IUD
I0JseNwhHHAcEPj2vVzKu/uZXHr85aFTkblwtMEN11Q9iQtdyiJs2kc/XyiYk+YyN0GxkGxsQGJu
kjU8Tokar13DqmaxLwrDvJfCKF5EVh63j/LONK02Uty3c1ye2FipM29pP9m4lbOlgKodC3pVttBp
jyxpe26yqS+nKlgV4V2CQc+It7reWNZ3qca+gvT4/9TiqHw77/kD2ozEQ6H1IvKYDLrz7QO1j1YJ
HLecDLDMocmFKpynmu9Gn6UbgZUnT9Z+XLHIW+4NQ3tpGLz4aGzFu3XDMJ81mgmb8cW7BUqyJn8V
5ICEu5wSOcOFycaTr+MPWjKmMrapstf+f+jxz+X8xbZeJLcvBrqdPv+cOM4Jl/7QA/riJKa2FXVp
qg4xCbs4i4nZprOfqk+5QThryzos4cANYij0A7U1bVwx9tvTDGuqJ96SElA+Tj/FqcYn44JfhuDk
nmjcHuD/CgcQqYF4a1JV3HDQpZttojSIcb4hnTwQ+bgT7dlKEaGHcnHjZc4i/Vh3+0TQvQqJF6W0
1Y4OAVROKBddhEUH++aFBum48sG0r3veLUcS40kKBYn8SqNoLpAtt50QHOEPSU4yMsU/NfT5NxsS
oxIa7Hycmi3Zuoj9qCidpdV+E8Sy/AJt/GWeODGMlh3ze0Ym6SZ3mzDrRkkOAi0CePcrDrSCFA49
psfqivoaicsUteBlNVR01Nru5IJ2KPtHmP+w7lnOI4YZqgwsA630Z97kYQhoqRgh3HHgM4Nvmvpn
03oQlzI/yPIA2FdozsF6+0uW7UDFjfXAIxN1hlODK9Kad8goWhrb25ZtFR2SgON4Dk4WDXM6gpah
wagKarFPlrmDTWu4ziO0VsnC17b+Haper/k2AKtdH8Mp6K0ie3V3S1aOY5jORBrudMhCUBBIZ+wA
pvwFVNqkOmb1e+tm6rZIbxyjIttfIe+ZSoL6lCBe0pnRmvxisO7+hMeUs4ijk2k2lHvlWQR+3/BP
qhSniAjHU71wYEwX1XERAg96CA9jG1UPwQH9lYdb03bSjABo2+EqSqttQL5mlGuaz7/qLYTXZHOi
EYkQ5nyLLEHS6KPYRsvIV3689mz38lhBxi8cYKXR/ZWlIjhSzzOTQ34Y59qxw4GPO4V6nt9GttnX
G/OQ6hMNxr0TukLUJyrozxyeqrn6f7fO2a+/gdty2pd0Nl0K0FKS2JeDA+beIWjY0Jds38EdUQHX
FxV71SXBpXZ/Kf6DbehD4/86E46T8c1jWs8bP3AVxrI0iWeEkihSlbvffybvzrOYI9rAMVSf0wqq
4WOUKfj5L81CvO2Osw2dNZPnruvSs+5Z0OiFT/luuTVNB4rHHxsXdUyk9R65UCoG9YBofw0TuJag
GYmExPLPEfkUTUQO77mURimbU9+X2yUv0bjk91ap+ptMxjpOz9s0uXr1vd9BjfNXGTTGCRFWe8/3
B2MJhwfz9leNkZfBr6UXApOwAyDiuKVCBsgvKTEQSJ6EtWJp0tC29Y/jcuKY7moS6qgBYpg4buC8
fSnmhLjb/0VGtVzp+VyR8Ou5RLHieRVpvQ4fSMidkuHHcz+1Eo65G9h9a+ZWQdbYGfs3UnPpzIaX
7F+69A8SlSiCrXJrXACqtq+v1Hr1LScDizYGs5Txt9EFufQfTJCVga2JA/ptra+R01q20WinBWU3
zthaj9ymjKm8rjKiFK796FtB8Jcpk/JhevR5rmHPNKGA9yp6dFAoxlSgCH4wDjivZi/8a6OAsKBM
PIE36XB6o/5JucI3sIxOXStGl/JVkwqZOOHo5edcX9IaycJ+Vv0ppeLsKjIDuNo+GEcODibLuTh1
oFXBr+ct5WdlhxkWsVFD/+K06eXBpjlarjwtHDAd8V65vmanH6uQ8A9LcZcT3we1kmm2tILaIfua
+Y9/DooMbi5/MNUmNv88QqmLIPEDj5qIxUmzh/avQVO9SRwjxmqQZ22ttr+BqpGezUMmqOa7N63A
4qvQEzOS2H6dH6CuddDWvoWcRucrsneKC8HhmQmOrJCrIUMYPKLiabz7L1YNUnQYn5KK7cI4QhhW
NsKQPyaOr9GhaEIFJgZnx85umbbYz45UlhBYPEA5bKovX9AxwQoP0GnWYrwm1Qxbows86Syae4nm
L0i85IZi7IEFVPTRk7dhjJGcdHJsnL8Ll9ksE/fxLgW70mbizhBlYXLNlAkrrYUV4Q5Y6zRT6WZ3
uR3i5o6RmhK40gKvNe8NjLOs7DyQuuailZbk7H96h/SFNiQ48Zf1Yfx+wkXGguDM/ifcruoY01e0
PdY+b2VPuNPfilNe/AvEWKcGjIw72NUwOlF+i5qxhHB5pV1S8d5c8Ncfk1Twlk5g8Yl+TmxbUifb
Q4CHDFKc7OSY08Phigv0scQvbNocyoYdppdSDUm+ccg8L867/kCJQqKam5f/mXI3yV2JsRYpcw9F
pMuM0JQHkw/OkQaw3W9FWFHST6QuWESYaSa0x5wLDOxcnjTil9y3ft0MfD/NvJyLGK0NOwlegl87
oytaKYzVdQjKrlyW8Xu4BGbpyHD/tuDa73b5RH+fhQYT4e/RU39Hugbbcn7HT5lc0BLtF87EXVhe
64GerMsPQ/tQFESrTVgF3dLQrLz3gJ4WQVO2SJIpbP5LKTjz1AZMNJCSh6HjTFwmGI5FMNuPMV0r
g0asFa406M2+bHnOyDIPXCP+Ln7M1RbzIc0rPfm9hCIQrA+jxyb/Cy93aEAQuUTIi5IyHyXdaxDL
v+NtjBeGX25C/IIDe3L+tE4vJrCIOIv5kCgJwLKhJYqRJM6JVSUXXlaGR3GooMBqO/CfOATumuT4
5ebfvfmUEz4d6NGILTi6XUSna6RS2QahK5akJ5bOPkeuv9cnzqtl5sA6dM5tB29z3rRm5MgaVH0v
stdmXjY2mGmBY4eMds+odkVsnPpKhCTdHE/KTYJsI9DSkh2PjIFeRV4ii5bOQ3H29q2nZwI41uJy
KrXypOlN4pt8GvRtO8aSePFcWcbwC2CLyh4S74iAEcG8o+A0K7EUIlHBD72IOiU1OoYUQJDsA8pN
OMitYeqAaAvo4IadGAsNWDvAQe5mNVMvW23xjPxoiFTUGrndvJYnJtc01aC6dQqkx5GoMW8/b+gX
HCe1SjCPS5NsB9ltyu6cduxbCZ+x4olSdEbPGwrBdcGMSB/ryLXZQLpItCvfPO3e5HrgJPVZHu0p
kl/0Gj3Fut0cPpG8Ph7Ffdu/x3Nwu78BP9s42D2EL/7s8r0pjbTS4YSRy1YnxEpzSXJIgCId/DMx
lMiI0ZlCM/CVeu36g9E6r9PzFtUhRE0CCOCWZ2fe+KIJG8IaZLwSCwhEu94u/yiukh2gXDTcim9R
uR8Yr/mpRbLIfzz5GYhx9XYKA6hfQNAAKre88s+BNSfTZ/2r0hr6NMNguYf1C1nVzxi/5sFIFlWs
AM6fhKvGmhSrE1Ikwew28inoTCbo0K19r0Dwx2ekBWG18vyG348zIRPxa0bVNPn7slnD1eEBZ1Gq
FrY7jzFoxLEltictUTY9QivK8VHPz357OH+kfN6mfXzX/Vim1QSaQcMexcUEboJp5FU4tQLWip0K
uCuaGcegp8v1NlLh1G1q7JoA0v94ZFH3e56jpKgli2TkMqPdD16ag0bxi2JiFflOHtK42qzCMP/J
Kv9AVFkUQ1bIIJRbr83ORa8vhwKwzMue11TlpzxruuxbOjQgxjrFYciG8O2SQWTtEfl1Ugz6pjos
DUYHDc9H1OqcXK+iQpukHP6mmzHiwmm8NN05u/zwW0r5COlNyYCVlQ6yr7bCY7UIVAtOa5Gg7Ii1
qPlJZWEXt7nGvlbxAQwMeDTFi6MGSTWSzkrwU2druxs99wb0RrbCbUvYsuGyUbLKXam5UIrDs6rO
xqdcmSzT/Sf4Llk5mXGEo2de79ciQxlKc/dluSpdLhKewKbG41gIQkhOz/pCln+egbw7CftMf+wq
JnxkUVQC3gXZaNAk3YgPc7vY34Vh81pyUFe/6IjnxcdFXBqED4ol+nAkAj5HBXVJJX5tneDuYuC6
Vnj1OgS4YCFiDkneLR+wWpP6Y/+vSbOeA7bTYgwMj3ITk0RnjJFXkSIz2qaJtXapiOv5zLKCJPRF
B3SLAdFY3eXSdWeufpocjMwVA0h3220N2GDd48qdAatta0E8gB3QPXE+h2NNIBp6sOzgdVxM20sx
ZLU1QCUB+n7sIGuaB64/fkZMBD/I8jNYciKBGBiLag1uYOKa/jzHo+iIf9ZJfQ0BurMw2ztfeKlA
vcK9eaT+9oL01XCYLEI0rI6DLSrb4btMXjYSrefJBx/Dswf3CTLvbL0HfFQwqofwxPmAuV3b6AF3
9VxMPaObo5vGD1+iYXGNIVVMCfAAXJrvAx8Qo+s1dLWAhlCpmHuhM5KyMAIeqY5Lb7AH9IPug1l9
qW2RuNcTscNDGF2A8vCdvSPN7AZiDFSlJ8Df7oQy52JuPEcVCSfep+hAA6kgckPkBi59dI3RjOig
Y87lGYFsUwJvA1O0kCSewbjNYiRBzXZmvewayZ5G0lJxu+Oyvb+Ze7PCxhZ8KAZ44MaiHyBMzDE1
TCjYH4dz6ungjkJ2INMLHCXuJG2GTWgibREtR1EIOg3XPGSVOdUewpfD09GVbgMjQCEAE7JG6ebj
0fkuxvGwfG/bkYoNqPQTevn4RmylU+XmvWnOhzj9RQaptI2jj3EA1rkEZg0MqSy8B3sLBm2A8SYc
hBvkMikrtA+AbKVQPON9rdIPJ0XNt14BJrNM0EyNhWXX7HGpo55Cpj7fgC5dOYq0c9WUnHvQyuOL
O4VE+4S5WCHHraPHvq4Snvw7h0rLytyW7994ELtrRQYCF4tPUKyGAQYkPM8eFmN5NtGtIi7O4BgT
otk9qBwb+Q2+StGx3n1d6PuKD0mzQ7Y0asEN2QndGmtu/VcwGRmXIf0KceIXW27BwybWkkok1/Qi
RZKm8Yr/QQ6OZbba1IKtK49DE1qTc26ihfftSuVMUMx0hCEBJ0pq6POWRh4EUz15xuB8jBTJOt9y
RhM5wPL0UjyyLqHNDpd0O7iAGfSsHIyhSYauflbHD7RX4wCAkYd6uPbCJDuJmeBanvxQb80bmLsP
+zxn2iJCILK23mdQ7UAoMNpIvZKS3U6LpzysjNFCzf/ZmIGKMwNLj0BThpTBdMYiOB4qQWdbzJCC
sSWwvli6dVqkM8uxoL9sFiC6SKgICjREr/QbxmraDqqiKta+x0O8FMHe5v2BPxMO8DV9KL9kAFUz
Tlx84gCKXn9ZZhST1ctiuaNY06pcOYrocMk4jSff9/F0Refx7O/P9X9dwP3V7CVa+j/csNLzPBW9
aUDwjxEh9FKk4gX/lgdxXffQdFOFImIRDmdIhOKU5DXf9kfKJBEVWLPSwj6WJY5kU567x9+kcYQZ
D3jI2uTarVFFs4mX6nI4MMcZbtgIQpFHc/MZ8z2qCArjiyPExMilSYQ1gQ7GzFY852s8xUixOWFE
9+0Qs/UpYyIf1V+TZmYpM5L8OuQ9dTjVZb6xYDcS9qyO0+zmxkxoIXLVROua1HbXML0dH2F2iwbC
QQxbPsMGJmzdKbLqoxckY+BtTSefvZe040k4D2wO/GVA+O2PH9C1F5s500ZQKWmTZ1AOar7k0U14
PD4mxdmGKckQWufU43RmI0ruhPdMMHOUbXcshBIq9vGy5iBEIPAV3fKI8oVXxR/6rHs0v/5bxDZX
s2hyMmpWUWXN1fE3UEl9zVfTIfJV4EW1NrJkpQRGfv902jZ1+w9ydNWLRv9Pxd3pLtpTYSTRTJA4
c+QdxXYf6xSCStdnEugXlnfsgU3E+ZK4BK+I6Tcj9QuOfY+zx/A4sRO9vxglVdgAd4bVmNWgG3iv
oyqzn41M5RuIXkjYZRoU6+Z1I1aV4eSdk6vRx+3E/25944b0RjXeE/WjAh38mjtIoqc17wA5HU2z
49Gze/kbJDUKCWrzVuGD8aGpNbW+rutCsWDLAp9g7f51pZty2olAHPSiaSChGPbp1AWMIPCC7wBD
Z8H8DwnN/KqKvwv1KmhbOlYmICCZzx53/H3xcSZC4EnAZkYfaR5qO/vqkL1dc0CSmyGtcUG7s6hN
pbPH7Eif2VJ3NLAYrZFQ/PCjx9emEqZMW3ucr/+Ne/mG/OznvYZHgMPjdJPAGABE3uZv+W+FsI07
7m1/5gnJXCTrB59qU/XVlDqNQ/5ew9VjO15czoe5RN0DPmKDT38w+2qtl7DcMRYieAg833blsvWv
HIC4fNLkslecov4PWvtmUOcnHt/7oSdqIX1imVu27AiYn3gZiyuNm9zNSRgB1wfXMCTGDaDYRU2p
CnLwB7ON4BXSuZ7x5598uQ5hW0LBhJ3fk2bQ/cL2SoZXm4BZHUAwIEMr6LmCbQkQsbFrFfiyhKuU
FdUIGCcJRyQNMRQTfEyzCr1l0M4Zl9i0adaLkNvU4wKmbcDsbTcfM5PMNCloMPgHWm5OWKzNyYn2
Sz6IZ5N/rZP6w60r57v7/rh4vn7C5dg768RAv8P4AjYL0hLv4oNmRSbf931xfPeYvM3S2tKWLbYt
S1yE/aNxsKXtqKsnSoyKt4N3I8eW+PBxsi3eYUaWnT83Jl7jNzNm//cZiexqVBkI2DENExZJ+eUF
Flbh697q0G/fKwlJd7iSfMC7ssC4NgEHQIaLQBWvdTZhu6Zb+ice7RLwvj5uUsWrWPWn9Dawj5u4
nlaN1GmEfW6365dZ5uR/wGhrDNfo96hktrRs5opiD6Ddr8GsatEdb6N/9snNQfE+1m+KG2p79hzj
y+rk68k8sgWXodTsfneKRzvP+tAVk7xlDH4iTpZogR2MKEfz5gxgbdcDNDf7vM+NaZZMJaEW9UlS
VdCSDRSABtZYsJ50cF5vPfsYbVaWIWIXYIYPisani81hWy3FEYcxs2mqoPxWr7deUqy0tL1CG7ev
amOACkRH8c0gn1rsmo3KzUOeI7q6BTMStY8ycb4OebJtNkL8GruqNBasBYFk9MxcL0oXvkL5lZky
6PlvYBhVqgU32GzXCw9nY9qcwsBFMa8h8/Xax7m3w5WYMrnAD77Ht6gIsZfdSlCHKYAGHJ9lIpxn
fAYW5ao/oTTYLyH6jbAMX/jr8cJ4aCy8hlZ4WlMqIy8XNdpl1TVDGW2+2ZNwplrWcTLuLMjTI20u
Wd+lh7uGm62zzI3EgeNGVzJj4G6SOG7+Gdq8ybED7yG5WjdTO3qt5vJ3PHBaVQcXRht4gy4qHul+
GtuJ/2fewnu/kjIzxqb60pQjAMnxpdElzFJL5iFb7ngJPHdeMcBMpo6jWn2uP6Xs0vmngDJ0pTZG
iZPGcxHX2DsBJm2aNbFEIy7vBZuTPHgmTJcnQEKwgNFFrFYwFLstXCE4w7eNBJDsTuEQli1xjOG8
Fhq/lVxcfj26couk+mgpbAQes3UUuulfx4SNdoBNGBourwU1sGGBbqapDqDGCYd+QOazpz9Up/zd
4AgkzGH3WYIEQg9sTfJeZxwJOpEBS3hBBeYm1mpiYf1ZuiFRANm7/5q4LgRgsLI5+bY95iEuN94w
cFZBpPzOxH1qVJjtaYzWHO+X4wFHS5ok8LSf3HtoHMBN/lN5QEgtaqbrdyfwYLpWHFF43VudvWzc
kIF0QRNSZExcQBjCcPDtlS3W/tcKmMLOYow062d5X1KuYhZ9eSHnQ6+PL/aYYjZz5Qz2D3ytVSRm
n5SQa9ReFrpHSJTC/+h6Hy0QYJCwtTCXX4ka8SLDPzh6ZyPU1ly4E+9Hu7fQWfFdUfFZbQq7lwaj
7mmm9yuKiE5hJY8D9pM6Sbu/lpZJkoGMq6TbsWBOTbdxrdhSrX4JiJz1huxnQFcst+MSc826BIqg
gFwnK0B4e7N+DSZdQDDeePFWDzOLAQjtaVasjr8OQQjOUxwfGaybQqHFqcZs+LfGz4Ow8acI+9Pd
UUihM5CK9D2/oXX7ggTs0XFLUa7FAIIT0IlBSSDRiiRD5NSkhXbURlMBhr02hjyJOHlg7YZVuqNr
4zijXJB408KKdqD4qWkejClTvSauO0kvPDaP95QshxqeO5BOihC9cZTdvQMwLsyTj4NQxTz+K9Ll
+PkeERjBxHp9g8Oldy0eTcY9NXpyejoGMHup1AYaLNUwGUf6TfOKoR0DMWeTQUyfA9gqnhGJ6L1G
aez0hujttI/WIZCvy2GCFjOACtZrq8TgCBZkTHZWlFu3TBqSiAeFb48l69DP5wl3pPhq4b0m3zS2
AffsO/0HSq1gd9e8y7NiT4tfNtbXjgZUDmrwp8lCU8Iet8DDsQDxK23heVvIhKJ3OXZpYBiX6X3l
cfiKp63mAu9jGkJ6v+IF4JW3mR9un0npxialScVkXRNVevnxhTWHnetj7H0yHPgwkwDDTkS3mt9t
VNJtmCBVcQ0kCoHfjLuNbQ6cfNIBB7kKGdDUSlG1Z6B7qqP3ARtF1iQb4fWnf4iLXZ4eko1mcBMl
KKSnIFP9gUVB1x13dwaGPdBAHU0SQ6mjCfEJLxtkFmFBUvYOEYedv+QwJe37x2UwmMmBc/tCSXyl
1/rBClwfz4c5EgM7rNzvCgBHm7SqGz48FrMbUDTwedfIZjSU6vvOiA7O187BsrTmA5b6ACl0QYuW
5vU4KQMTmamuexfCKHEijn82g3Qzjssg68ImXiNWllfc13JD4Y2uSfRLbhrXZ8kAvTvPw1tunTUB
oBCts1AJ7mWHgLvAyWDAoh2UCcV7uMkf1Ne1YHYmLY3mOn74rgEHsujRmACZHCPXwuOxm7Xq9dSM
WVYfXwlpYW4xZ9I2jkbclwXH5K520SgVHSzSc1hvUHxcazkFDrLg9hpZZmrnWuvGgUtwaa18ATuP
ui1WFG/2/B7dCl/+sJLIfQb8UqhDe9+P9ccOopv0X3nvWqnhAAoKbpykLC1SSuaDe/7N78XdP0Do
kUvyI+B+2GlyO+oqVJJ5YHvNkwaam8jCyVc56jDqaI7hSE8JhsRs9Mg5liniDLo7MQkbTOegKbz8
cmCJM2PG28xkL98LG2YxJrl+JLQ/QTef+dtkHFrw3Eo0aurDWnZLyR9yp/knrR6ROOtn3jD+0YlP
ysGAsSXXa6glfeKmT3igAf51wSXgMD7YBbCi+jgkX7x1iHZysnYjcXjO5p0ViP/iryfcL390tj/2
KMENCIF/w01tqIY5ur4+/33UGLkREQqqW+Q2+yIv7fHHsWkr0fGuH2J8qy3bqOvUbPDtDM4RQxWn
9FkkoxBk8CVq/qGb9+hCFZREOGhtL0cFmZgZx8584b6BRvCO3O5FNBo1JXq//VcCelqGjzPf88EK
mYlN/Rg3l+Ils1uSFFgUTAtli2z2vysybI4BVXWFeQs8biNuX2z7VLwT6MtX56KACdrPijJu3qAq
sOEYkNxRWLgpBjbY8TYLy5igUMLFqJxuWJ+ok46XLgjfBglErBFdc4EL6dvcNgUf1kF3owPRvKXh
8xwCAPWn/qvua8D0DOjSRL6mB3T3O/AqQEbEr4tqlwYGm23Jnwi9waMkXjXxU9mUY5f6pFcRcoBD
DTOp8/yTEq2i1FELARNQ/tOKmjYN8tTUJ2MY5ZHyz6g0DJNR0IYBVitELmmY2XdIteKrhNIiDCgt
0/f3kI3ciOGfpNCclUN7jZN1jrzKnYVX6UlsAEhK0UA0Vi181gAdjP1Uz03X6LvwCQs/lJ0JzIvH
as+5J8XyYspf80oW/JzuSrhIn9no2OZS8kdjsaOGAP9S+iT/kXLsUF/16f14tBnWaRLn163akz8J
98GH2b4Nr+Ipziw4m/oJNlb0P0DKFEWioQnASbeAxiQmAXEIEYqIw1JFkQI2KVDOOdlk9xOu9vrg
qa7OOkg2OjMNi47dsLOiNf4XkZkV6AT8fuGBpnx1vRf5PoCyrAE2tWp1QRXXAP3dCRZncOqNKRUS
ePt6gL8apeY5H1eWl8znwCz5/X+uiNkOXc+sxmC+Fa90b3rUzFXcVm04l79qpaAPT43Y/sFOL0qf
5M0qrbdpCzOkAMXHBLcUhPQxmSen5czq5/SyyK00HA96kP8HNmexNocy/jafq5SsfJIYJnMqAVWy
N7U48vEOFcUNxJYxNG9e+uj8av5Htf9/GOQxCWXG4kO/5qY6fzHYuM2xzQTNFBlerlVagtcwqUjG
Dq6M1CQuqHJ3VyzAIk0vGLLpxP7OhCNVZjFAxJAf241OtYVXn3IFr+VyklJizWY9IT4kFlHS1UX0
ekvs3PSkLsitaYkFwDGM5S37Gdog60veDf5+SHDP/28wdmizVXjo5ZMh2HRcV6Gk36U/Hx+UgxUs
ureuv9A6nLXhgVl9NWQtdeooQcjHsUZWwPj9fkV/YvkRSTEkuitj+1BEvSJvMOrzNDbzIYahiIHI
ZhAnI+UwIcK//dsy3sPHcMbLoJOa2pAH5oeFzAbToc5jvVUDa84dmJDGoAqCB0Yl3Oz4Sgnm4MNZ
KVDu6fgxD/bs4/V1F7CG3yH3Iv9i9yM42NiJNosjW8g77h7WQ7n5Ix/tX3KvZjlNr1hT1WEaCKAT
6u9y2MetGLYVgl6ttmerX8qSJAxT3zHJJH2ytoSOpPFZbHpfJqliZAxI8YQ5Md/lt85qYJFoG3OR
1cjNvb+hQGf6Y3/AYCj16/i4dOxTDJs4ca6sG6BVQ1k4To2R8JnszJOf0VtmnF+D9+AGT45JjNSM
pZSJaXcKWgrh5C/aSE9fBE/TyvEoNEuOPNtGFgVJzbCOvZsMt5ldzLx10FM3LU+J6MDGEFLWvZsM
JYEHJbDK4vgXFxqfjI7x1c2q5ZltW4L543TFaIjOU3b1Fd4J5FE+xLNFOMkWvk7VRWoOAON2ZrSm
C6sZKku6K9kEqG52yziQ2LZ3kom5I2WFPJNVTL8Zd30WGy+uC4YqXzQORoRz4WB88r9/cF01nuAZ
wGiONCZxanL5dM4BCRVldb/yZ6qTJz+630qWCH+2aa+jeeBs/sZjhDeUb8BT1aAzFVIbVhSGOt/2
4JbGcRgeKJpBidPH6kFcYJLxY0a0cs2DvHunoQuenrNL6JP43a7/aO9FaSPjSSWqT6KikPetJGB3
PXHyugq0duNQKHpicDeKDniwXlUG8a2g8E5Ff1onTmFniR2bqsqVPfwAzVmsGFW1KAyPO5Cxi0Yb
WXqtMLoh2h7zOicKjk9DiwW95ARCWVSlsXQ8mQ/12IgkcNhAFoxLvDERYGOyh+GtgLI1KVZjG5Zi
uKb4EDhQW9Qh3rJ2ix6VNmA53YgIunwZH5R6pegivucMcF0snmzfLqmFVpcxrV3+ASuKNf09+8Qv
lxwEQaUcIalYALzgLJNwBjQQU3MKXpBBdLuagF1IGjnErALM45rSVybvYEShOcsoeXagvBSjsunc
KzT/dGsesY+oWW98F6Qwz1FdEhuXh1V6GT/1IXc9OIj3VNwt8kKPvqxiTBZsrguTwR0YfZCh3Sx6
Qh4N05otm4AdRYbiUB21dVy8gRRQJW1PkFDNpOvz0cec8yhHGnkeAAR6gKJPPOkJRi0XomG1+aqe
5eHp0wnY4ywP1OYN1iA3WnuRWZQg8c10C0ILnRxsAc/w/oluuGnb+WOBi4eJhQlOZ7MZJGLpZDs9
LQGtFfksFra7/U8q0qEj3Eunmet/Ozw7m5p2BZA662Ow63o3rEQzNKsL40w+w0IbtwN/dr0Q3Df7
GPu0mvDl+DvV2z9oimpWwDpUVNYj6EfTWMYA2LP30WHKGPWMKBYFUTibD7cNLxiYfk5YngbXT71y
v5nI+ZNpZnVnCOVQxWrElawI9ADYMTaEgbaZ/agrzkOKK6+kHQEoDYij2sqMoGo71KJKCur9Puc7
6A3ixYegNBOWAFRN4OLrtisEkg3dpzRFbnR3ds2/zH/vvCNiY+SCNR/IqIl1Z5ZPkA896+oxhqJu
9DSwvl9xqASPdfBMIRwEiNFafPXaZYZkkfSQ3LFO30X/AREXCaWRabdD7U45WomsDtct9+PUbXeA
zXqOm/Jw2y5J5BzghncZEk5MU/SQAVBstjxASoJffZu3bRsIx4aS/lPScpfwVYu0Nv3X7AESx5at
3/UfOPtM/d6kBWAgmEGXurpl1xkZFv5d1t9etQAlAxeMvQ9jPZNIC2IPkiBrXDt9bqr2duksBXR2
imSxKLx+FmdNZj0haWwVTKmOJ6AHKUJKPWw4FaLUNd2eZK/XDpQow7C/fL630EXSQBEJsf7xeryA
91Gs0I7ScrVAP9FACdioIRH2nfFN8dDLenX4ohs4othneRlnBnvmqjonpab2Fp4m0XBuiR8uKLhb
8y8a2z+e8Dpo2JryRkyU3Sw25TK6/RpzcmxV4JkQNTkjLTXgu47Dqnrkrc2UNhw/842N+VsDAASN
nDQNEbcCBBBlTpwJl+Y5eJwYQWag1PTUAFpsG2nRJf5Q/ckdrY2IGfX+QWBNtRTa5+ajEDbtZRul
Y6rxZ49n2iMIst2n2w5J+4t2uMCfkizdJq2LINQTeHGmcqIMANL1v3rKc7sP2qtII3Cy5j5Elwgd
4GinSqWjLjLdoetBJSMalogAfObabYowxS4rKfvEF9+vW3uk3TZ/EtHVHIaO4jGxnEferOWpypv9
2x5y9H718DXVuiv7MpdmRu8FEoHwlL510vHwWdSdvUI0UF1CC7v6KNREguZpxGgc7fjBdNRvlGvJ
RzF9rFIMpkafpez8xesTVIhUyDDpgWmf/94gc1uXr3aoOIzTkwayX4e9UX7733p0rwmDP33YQAbM
fFvCcaMuz+e0je1xFTf59aL+LsC2OOg60yAKvBqnr1nmIYCrAFgRVYQg5CGN827DeHj8uQShzxtz
EPJvSdYQgM7f/qbdzWMLalE6G28RkwqtSw2XNCew1iaYdRja2nGac1JShn6G6DDOHN88K44LzXY+
2YhNNXkBJhYP+lm817phTr4EBHL1eWoHfpsq5YR78m8Roi3Lwa2fEezF++HMjfn8Y/ZYUzjg/UNo
2+O5IHDtLe2yQZh0rMcWjsRi/TbPUyn9nPzpBA8dVWDqLE2WQaajTGxAqQb+d2skLY2hwSAusNQd
FNjxLy8JkdK0fSHMyyI3wmGHtwzWfMK3fCrgMgcxLDhlIfTC5wVTIPL0o0JSDzX9+0nub/5IW5KY
0ap61gcDKvjNcVQPCZpLRkwsk3rWoaUvOCb9zx00YBAdM0ve277l64KjFDSPmhZrikGB9xTNyj6B
nKay7pC3j9kT636LJrIzuDmC4mfZZtgt0UR/FpYE/Q7qQyVv/jwNyi9TpxWAmKnJdocBJT8PEOPd
/LNmpeCBTgnVIvZN5bdmd0vVDm3Am2R2FT/ZQK213gG81b9W92DkvTYB9buHltawBOpLfguuzXMg
yxwSOLxaw9NPYrQJn+83l21LAkCHWIcb19ruBrLGcRfLQlwYOSh/Tk1SANg96G/gbY8C9V+V7EWC
mTIZcW7rqTeTstLSEFGLaWQCIgARanlrz7VM4ex41KcED7vlx6LDazcEo/1jLt75KHv30LRalKz0
dD67savC4rKZwrmjaM+hzXdHMh4N8TJDhhV86KfOFkXvlTTfqUYs43z06Qy/tomTp6lJJQmC98qc
XHdFSCdPPB87A8uUocqRg63iJw3Zhl+6sEXfbIfA33o34xizqZvSjlQryMsL4f+wA3LqaIr3TDL/
B/HojhEguzlOFXMFgPZRQ53OiVvWh1NtEJz4/Cn3e9OPYbwM41MHImQz0JgLV1RKtjNRvjXUEkX7
MlwAJxmAcLJQBYDm/kRQR7E3jPBpOn/CX5zUNy74+Jar8d9ekBog+dl0Ai19hV9Q1QCXgMRYgdvu
VI3sZ7axp3wCH3BdaujnM8MERfXg/mBFbOumxQ/vM/I++CAuIc30x5d0rRMvWhQAyXKobr4zfh26
ML1SUe7f3NRJmYl3q1W432F1yCNnGtY1l1GwVrY5NUKcYtXYWCggTlocpR7ptbYPhE6KR10rCqJW
M7PDQK0OdQnyOWrrAmTDr7TNg6rfc6FwRSV3C8H/vkz40fRFHOiCdb2aLADZU8QsFSrKlVk7IDzC
j1mBDYyLL+W0didwFDQpDROxYF5cbgpr+DCx+rrbSnGR4P2qDeEEZO6eKb2RSUVDZzxv0Hi1izWE
PY8ui1TDhYS5Zb1Vn9xA4D+ReZZWiJn937sa4g+EJsBfcB6UkwxhwE5sf5mMkyv6Iu7NygTwxKm/
Td/p5U07gY/NA5klgfnz9aWZnaUWh82sgQOYICtXhyj5zInP/NTU5AkLZRcPNfHXqK769k8s9/kJ
f3Zj5GJSsNLh6SvXG14EJS8KKejkAbsgObG68F6eFuTqNRFGRUoO5WcZBneInIW1eDs2NqG0Fc2Y
E4tMiTKqjL/Za/t6oNfu+xdWdyPZQNZkqDGrJpnelqXSdFA/tckG4CSSMGfrla1Gu7dKwBwimGsz
FJPuP5GQWpIk2wVUoDLRJl0cvOt5NsQ1Ky7pieuWchs3ayo03C4QuYcovAT9xO6797hY89OOYSah
uffWIYYeCOLukjtgZVUK2dweH7e4jgmQ148qUU4dak8dU+GOz9WHmWCUi3ubMyCwGF+TDhsGPIPt
BjUnR9SVT5fr0qYirv2NtAk9eEzgyR2kl5QKE+fEPOcUYhmTES3poTpGmDdyJHq4qjl5cMhXw4Ax
eSmE/lmrZjZmf+2QEYWE3xIb9t8lXIzsayrFCbFmZ5FrGS1xTfCLYyDEWbi8c1HPqZeHY8eCK6rw
vDDj3zSibzDtMnDzgQQ9dhFBxNkvjG4M5mPi83XTWGiGlS8oYsGdG/Xs5vkmFC41maiBtflXkJAx
9VRSOAnkA9jcja5H11X4GpRcETsTXeJi+nbL4HbjKMrn7m79BE8wVrA7hi7RUaUte0KAjt6Lq+iR
LAb/71WSFosbV9wZHOmzI40X49hJycMOMC2BjhU6nV55Zb1hztEg9+MorbC0G2YCeC0gv/XMAk4M
HYBT5n8jCroiy5MgFPGaKjHLJqW8S4ycKsxZ8CGpA+Sib3k4j3SHGfl5v87KVHDIiCBOFEVRdNyV
ZyaXRihL4oCHHEGumlI6gdkOuJARzyyU/nXFqeFq2Rogpqdz9nPsqrMjbSMFtz4DSpACF6QUbZ8s
mmIeLSZCxHUQkGmmt7x4B93E3KtnEEn/7KMsoFZaJFMIek44MfDYNXodry0Is0qeInUJYtsnFaVd
a0R0WRA+vT69UDQLqJQZSmFlPCOBmxvA3VG5zO/InY1+wEnWd2+xWec6NmMCXXLL7/M0fSeXz3Nl
ZuggiNFcRDXDrVfk6QtbWhveCiQb7vrGPAVAbbf5mvDySfY9Z5hvg26fVBrymjOQ0YfCbV2PhktE
MkWIISCLhmCo0hOz82YGuFaFQUf7GDAOHdKwnkStdTbhreE8HlkG9Jkwtmy8Iradain/YQJ/ZMBU
tJ6oHkFOu4wDmwB03IaltwSaz9Vwf8x4Rd3iElaoUO/IBta/OgN6bxcteKWsSR3ZXhZMXpURuTWw
mNthXnjC7oWihFC2itL+aFwDvPFi6kGkW0ubkL0s4XZU7g2GKY4S98EiNY9wAxNktqy4ij5TFJLn
MS5GaX8YdeVW6m7xVw1Odw/j4Vhso3r2tX8jmCRK7ex5lSS54gb7wi4vEt0eeOkeYmjdrFXTBWGd
oxD6vBlEeOvHbd4j0BmVI5vk4zwkBGR0h7S/w4GidXfIxO5fJi9uTKoZ7yDhMkHdKRlkTozqq4xs
lWjIW26/6OW4Xruwyt5zpF24bgXUXFLo25WsNvmcqNP7mdOAMueNCJr858Gs+7L8HrSAR28S+XiS
1lxMiw7Wk1EY+fQ+7bLe1f8IIwldT8NouXwC3xRMpnswt4Z6RU0JcSPMF21jsZZ+bMiSpdnDk7PA
3EEMBnsF8C4iUFtAtPhtWIu98Q4/3wk6oJlaCCMDJMewC/80GxWz7vyDTSaWtKKrRBLwp16LlUbT
ae8CrL5uLdRuhXOU7Rsyv6Pkl2SocyGAgMwz3NXQhrj5BcXsWP2SGRZg9qwSCzlpNY8ibUD7DXKm
WFiUnEVslz06FrhMZa130c8y7IF7UVxb+RTIPfQOP1uapH1e7npaH++s17muAcA+UzCqmZ982bbJ
Lp5NJckZVPPE/o7TWtvvg6dqsEylk5dtsWERfMHQ3ij1XZx6YwBlNyQY+4GRNQXQrOHJqHZ/v5X2
lR0K78EgbcUNYZIQ9BoGFZChaAVBOGV8NfcAKLi8lqaOS0u0ZHJMda/XTHlnda/jDxpZ3oSWelzQ
a5T6RMHbitR2v3e0bDXIvXYV8OQNQNDoGE1L/6Kplq3Tc2hjoE4F0+RT/0rXIkIpKv85nbjW1otA
oPYlmOYClDsAiMhKjgRGcw3LlUBnmzq75E+Y0fQvZ9cL9wymqWyl69L5QfvuKgO6YZaYhL+EbwD4
75ZMCxWmRuSeXVerkk5Qp7+3i4mbPQndW4EPxUfgeoW5qxN7eXrHjbjRhwP2HikJPrwIAk6cIrKY
1aOdZhqsTDqjHuLSVq4lTtE3S2W/Jy7b9UFeT3LAnA+iNQZpFf1L8qPh5ElvdpoNFhx69kUy7ozI
INZL0Ac/ZZUzk3lRg5EKy/PMvdW7o8pGLd4m+pooYyjhmMQ7IrvtscvkxMq51eS960QrLRwY4MRJ
KZ2ihBHyK+4ACTEk6XYvlypKSHsJxbUMAqiZgIMEpd3R0vRmiQ6QGc+evn6KGbV50XduR5HlNxzT
j9vulwu593zUISNcm14b5dbaV5RGGHiRF9QMJTjFY26Dt5icIL9iaTzCQw+RG6YaVlbSBETsVfx3
6TyfrkpEAay8/n7qbUTf+js6OkOBDpq+RQVxxVmznaTeCBp5qBtUx+YEJrATAeOR9NpbU69AcQ7J
q41AGcVOh3dIS6rFVkzPcpNvSsWJOhLX7kufLYnJemGyW0qTOxqRkXhy7QmXSAjyXlDeM+sUBS5i
RcdsRt7jBly8DJcPCV8sSO3NEKp8FkgWctJj1kj+P1kuaA01eG3nAvkc0LhoupBS7gfz6zawZ1Cp
vVDzYsqMJQBy1cdRtlMq0gkIm4y52NByPLNbqL6ijkg7r1VSbTzKFfHdOflLxqP4oa1W6X8n87+0
GQ/cyS5ws63QnMM3QLEQGtgPNen/rdJzDHSF5+fPmAsznLpLT3rfK7awJACPSrT5bVclNW8mecHX
pPPSOYTIKxvKZApNHMdl6+Sll9Yoey0lDACej/+lMNNy+JxAoMxI55uk3q+bdv4xeIlFXUcMd9n2
BZQQSrt/1uTdYebLqXZppdkjDHxinhVrNh428uHODXHqh9vSb3kvWX1B8OSPfYS2/jiEgmccT4nd
n/dyzZ+/qC7F08ei/CFL6T16X/04k7EPJ2vYBZXd6JwOcTSkyE9dN5ltp4cgJM4DlvptTpM9PkFX
QxCjsUm2ScEPbAzT2cJxzqe1fxTB+TCv763g5upnBoQ4+0dZ9FmMM2uss7iv1QRIGaTQYY9MbFkR
jU9PIKBYa0RckBOM0WYekpkpbZcvpzqi5ofewtUxslnhnlh49rTLJbCK6xRMVE0Zve89jo6LIhKf
uX8XmmJ7o6rqdEXsE3la2C/cSsSNoMacrcC16S1Hr0sRjDPHdifFCtOx7T059MM0FhDJgnLY5cAJ
ALSyUM7LkXAXPx7Iaou2zyO3Pyg3MKjuInKXjEkvY5J9X3rXGba0xJjSmFBhQUkqNYl7pZVhJrAn
zsb1842mheREvLTp57IJWqQxN2isX1gpKYvv6E8xjq1z8XGU99PXIBB63v0UlX7HPkwBFZHrWh0k
dvTQoZFaHIjTfxviKbzU34F+DBHqK2+l5iF9dW8HgzIk3AY7GtglHwxrIKs0Q4uKKsL5BP4Ug0zm
dsloCeKDs4XuBbDpoJoNqrvft1f2ruFIy64l5oPbWs3Sf5ce1pLWb6G1ciIDfkc/StJb2Orbq03Z
1evuGQBu7Tkazaa0DcAKQauasuxAmFIXoWMR6Ey93PAiQ0ZliThQWFWw7z62InCOSCy4hvFZ3p5h
2odUNN0fqttUCoVwBi7gKKCqZtK9p83SHT7M7mkgKXaO1xUfE8I1SozM8VBeXGclQDF1gwlIyh+C
3S7relWaTD9/hzhPHwskgkp+V/0M9MKojMh3wCTtvMZOx7+7QIn792jmiNEoVbBNln1081D1OVWP
dSVnEp+pOo+x9I/2uGB9vqXn0MkLsPS0BeD82S63DQytlQxn/mTTVoE/sFjE7mBbMHDLPb3Wn8Dn
tUMmZ5LnNGRvBwag9T2pYXwWSe5vVLcSyuxcp80YFgywwDScVtY50TeaWAf+JleJvPMdnD0k3kFl
44z1plekmRtAXhJOGikAOqDOEYNluVDqgHwR5DtgBPEufqTgIwfB8xTlw/1mEIq43FHrdo16ycTO
a9u6hyOJAjGGUsBeqTBK9pu85OzapN6pv+aHWdjPAcntgqyiYHXh8lFbKA0dqvWcBLnvNM6xpwfA
e6oh8vSOx2+AUoJcnYWNsgflwZTUynegjV37frTxPqCulWXAzH06q3k2WKnrjvkZwwYgUbbhxva0
8uazvDxbSDVZFzPbZgSMCy99Lj88PLRG3RKZgdlDpTGAC+mE+Txc8qYbNJikSQ8qXrAY2kCY8TSY
hIMJmQ+kNK6RpPafDfeICxcqglj4ovL9uPDWcTb3f68M4XJyKEVm4LhslNRuPOXqqp58UHlalV8K
VmV7dqAf6H/+GVJ/oBPaFETko+wfSPnoqSpvrwv/2pVQyhEVyq2IW4RmqJXcNDVuVf3I3kyXa2Sm
HisIlhubH5stHEPUmTWFEqzvNH0FL0z7KPr3gYDrEaIWFsmU7J+juCawn+lee8IcxJF9hkZsqbJ5
h4hUqpPDVsuKnTO8h+QjhLxB8OszvpnRNYk9xwGverENdCGWuJDYaz0UFNRGJBCaeCwJkUgppgN8
OOiAUHkK/OFIFrItgmysIIe/OSfdWVSIzPihw6U+xbJJ4p2vE3T/TPAjhJV4Pn3TgLPma0RcU7PO
zYHZRCvjHGl0iG5PMyivIW7p7piA6udVoaS+zmWP8gEL/Fxt6FCPQoUF85Rvd543WxGmh2KsmsdW
sETwYdSM8XSdebTc89VTkhOEPCApSwJJ+BclemodbVERhQAsvVpQSCYbyyPsQtEnGaX0jwpMt3+R
39v8zkr6MN1tCHG+gBjz+cjEqoI+LhTsvXGgI/Q97t93u6WnZyv2AV+tSUa5Go74UOcoeQKiWZkA
3UMY+9bmiVwDc5/YOh15OBJyicxfQ4Ln5ZbTGrw5RSvbNnhMHwVJq4kkd1yb5QPSz0FNDpUzHtAz
U1m/UHWtYxru4IF2UXPVHiSK7UxstUSF9jS1vArjUtgg4B8S2yOrcDslP6kvRJieoQPi+cd1siaI
S1VKO6PI1NBBX1rdrFfSIqSZ2OgfzYAw66PHT1Qgt2XwqfoI9mJvx6N/8yhcXyI+/5EFveR6ui2a
9j0dy9j8QVOumEFrN/yREzzBzJCc/fX269jhHDus7mwwM6/+CHyWeic/u4qGnB4H0aFIspT2v5/L
I6eDzi/2QC1JE5hP/xlmAQaAHMKlNJXT/rtkwh1Rg6aA7tlV/Ik+yXhzNn3DlrdFu1hPsB19dZta
/yhORilIXnBCaXeokhIaukwTJ5+jcr0+b6KFgbvl7g1WQjs0+4F02kxr7pU0+x5rbqhf1nZMYHNc
2tEoCmhqitrhxDyiUvd5Dvm1ufXjMLu7wkkc4K5iPZ0gGdpLl2qkhkk6Kdw99j6XDoLb1WV8jufW
t0JCUppI7DMnztzb/DpRN92h9s4pKZCtdkhEEYXTcsF/qf8O/dNoWW9DKFy2qSi+QPRKdq96YQKZ
VBein0n3v8a/BCUsIb4i7H83rFHepAKndZViStNEakIZzn6lTkVLBwHDdU7OezIV5gKWSjLcwc9g
B/I1DWOi5gGm/wk9ZjHNjLEWR/rCjSKQqrbIYV2SumAB/0SDREGGRhb0p1HUFApqK0zX/dD08O+o
6DwZ0CJEOgITimFjr5WYerbQnx5ufaAElGkAIzX3fNXVy5zUoC9oGI7tZU1YR6vqHAx6vi+nLs44
pE4umuuB05SLaMzdUgOsESxhe7SbNQIK7bNfSVwSpS/fmn7uWFXHKgUkk5fpzX/SvXwi/QymRk7m
Jc4NzcJC67cLr0og68zZoiFJ7QMnRupoMCLV7p8DC0p0pcLMzwCPSJr1vUtmErJOQ+p/BUNluFou
D6dMSET1BZto/soQVlnkOkcOmjUpNjcKKckqiBwRiqvEVpBnh1oEsGlMEVACq8B/xnnZtHPGll9Y
DEughUae93ksA1yynXOC7zD4EnYmE9zaZxjurY5dUjlOrHJNDQG4OSDofxFkSedC9To0KjXthim8
SRs6PRETzAponFtlqmtOVMighnHM+ZJAY+NArVUnUj+NGS7g01ps09H0LB/YijMBpeo6ChLLSrGq
1K/2wKuvqW2M69S132U/KiG7/PWxEQ4B7/y5KwWFbsc5yifyVoRK9jSzMTjrXLVTmTXn4HM1c5h9
rm7TQ8ORBK0JFVYwkcFCZ9zFvYT6Xunt263Jmk6Q5xpdwkt+0Eo8xFKYuLI8jPYUNnMX1xoRLjdm
JwqV+QvmypXTFNfQuDpFaEWi3I3hE/Kv9WH8m52WtT7lRObKmu8R37zGEDgI4pTzyjps62tcLGeT
FZhbd0qYhdeUBThXlKoMS53O12uK+Qurs+J7feLMmsLlbgTsHxrjpTPi9hefAloC/mGIEt01wA4/
UZo9zls+vQChh9PMyQpl0qzVlurST21fpw/HrMLqGRrTklLA4eevRv+OEo6uWfnxpULKyD/52P9o
rRruGCfNKGr0Hg7uUSU85YjvDFF/wYf0F2CiSiz1uYbKp35NRKvxTYEBJypLKOOwg9I/sjCUG061
9CkZMWG+bQjne5zAmfloV+gglVTpB3NITVwdGxKmvToCCfrBijQ1sVXiH5vBhTOK8s8wkBFh4Mb/
TnvWivLZjmTQ99/WlufRvgig3Tekl5F53U+62cOrxz0KilCqMKSxzmSW9OdRs7mQ4fGciYpgxh6w
/ZX7Fr9LRbI6Hc+bGUXkVWCn+bKvdf5UwrMvpRWmWnv9nn3GpzdEDarkp8o7qwtKFb4LPfTZNkQN
H3vsrnAz+dCHw+kMP32jgo3Kt45+bUpzNbOD+lZS8t0MdtdRoNq+fQCza1392hpfDzkI92ZjO6Zg
vr3thJYavkHI00lQL2w8CfhD7fHGHbbyyzU0KSnW+oA0yROp4LaUcXH83HVbxqy5O9+T2Q+k0Lx7
gBXzVxEgCRoneSj5teQQhhMD5mKfQOJeNzaCK7Z3wyuMP83yPCRIS+swva99DBOSdf833p2nhZzc
cOjBtKwdnzDEpW+H7OTIcsLMbw2mUwMX7QamMauFNOqCNCsldd1PI2FLhQlq/Y5J9DTaFKmWyeE2
AaBrnB9RLIS3JeUc5+5lMXnE3ryk2SIAL5aKBKl0yKKt3Nb7ktoT1iJbnbgRbUAxzHwrcbE16GnJ
Y7uQf4TusWaUeQiqqRxOuHK0uU82znlpBGGcRfYQcu6VSQtOQqiuAFbPT2GDKGGQlV2QO74BKUak
tRBOCM59G0AjsrZ4Az5KjEBVJE8qz2uv7Og9SdkKX+/nWE9f1p7enXoY3DjzPBwwW0sC4vOZ5QQY
uwwq6NNDhpLEDADnx4QR32gpnh0FepxU9ienwNUxNgZxxFTmvzYjx0wJdv3I8JnBtNmtQbRNRswf
PNmjvImBYO/+mFY1GxTEB4Iz56WNjNnVdAdS+7aWGUqOtZlZEjkKh5FUC6LLZQPRYs0p5Gd6Uhl+
goRq38OLI6EPhokfyxZlwrh/FreEQyu05APMrGA9gnrWtTdRQ8CbsovnkCzCwl9fQeFgjf40gLAF
9ZvukGCueS6AatTui6jyi/CqPzDh/3MZWzGctpF2SJV7zzQMaBAFJ9klRB928hLxAA4LP9H6XwGk
pIvs2hq9biLM8964ozDIH/ZOr04ifIjdoeL8dBKIwoM8oxVFD/23ao+yCqWEA5Qr2NyJyz9y8ZBQ
DhE7yjbgkS7BnzGmaE7yh9XdV+WTAKrz7Qjz3qkfZ4ZP0x7LjX0Z4qRvGRjU6HDVMaZm+jiyKjV9
2suTF2hwPGbCYDrD6oKcbCt5AKzdEPEcCkQI8Q4x662Q7eehmqu/7HD3Lw2Ygkya2lfa0pRhErm1
E8eBalAJ0E9/qrTx6et+lzwTdhy2tKHC3oWcSnZZJzhJ2pyvSeSCPw7P8FNptzPIH0KSNW8jmSXR
1BR7yKlKkzPHq6o6Bnbie7C1HKqa/4OB5a5Ll3YgOn21iUhYRwMMATEVPsYkfBypND73INhj0ION
HHnPkpIeYyJb0jXew8kc9En59bSj1mI5Uy5CUp+LS6+kf4K51ZzQKmAh8rqQqikBKIAwAU+gynWo
+AsLM1BhjYvnkzreSxV2Rr6VTmoenQGW+NvVONcQosVb0k+LGUHp37XdS+v0SzexX7ih0unEB6dE
C8l3Xc/MqlWphTTBXkS1qynVOufAWlMTLyCjU44+5zP78p32yZr8IEzQV2e05U8J5DnMHaY11Ll8
GixVZJI4E37DYMr2941rFC2zNabm+XAlas11dFBOH4P+qry9bokZiO6hyFe22YLTe0Qm96mKaEoV
TxMtKLsJgSCnS67BwNrdZsafI5pDmDgsUBDEx+U+NiL4t7xoL+wpzfvrtzWylJXArVb3w34FwoZH
n+fVv7wWL2kTjzQWbtH6t08gQolAgnv1PcVgxvDhnY9JoFqWPg7d1JeQBILL/HzYlQVkXvw2Pmht
k27eNolDLwLwjlHclBcmAl/5ffiwr9LGCys0S+aoNKEKeEVS6yXSIsVL9r/L5VqkRIM4xForn1f+
/rc5HM3AoorO+I8wv3x5KMmk2eBlqS3HWVtcCiwIkgBvHicWxKmFuo1JgzeKzaYbGEG3bTX5PPm4
RFEzqZzz1ZOUbGJqPS51anvEm0o0S91R7KU3nRBCOo3t73xFZwFtBlv1oe0zrZTVapdei2yIDaKu
JNl+K2MQzN4XfPDVzEiQpSX+/c+RmtjYgNRGdyG2jLkDnFbxL0zHSalnVwQJAs+4EDVz35078ORG
drWcRnsKwUsX1znxVbTsemuNrSrKOwK4d/MKw5gN7UM56VRML6hgLEv9w4H81JVNNWEmJz1z4jab
/5mL7Gotxfp8q+4wXp2fxue6rY3/CzvOZDtNte2eluTw/iIlZ0xxAYAZBavcPwuO7ZeKmwRE1r0r
TV/ZzLHa0u4OsHuRzxjCcO5JCD3FzzqQj8y5nf8yc1AFhFpNaGBhj4Vtzk6g+BEFKFjt723sQFgz
ILUgZxVRvvZKtATyDWM5NDlZStcq+kJ42yokL53wPAKJ+P1arUmwMwwHk+2ZNCqNG0qNcwKpxAdq
U9Zi235ATvrEzmebgWn4w0EtSLhFVEYuFTdk7gLTvcouFfFRkLjNyn0CZH8Kikc6YsV3clmZbYB7
I6suW6JRMl1VOJDPvju7bUNNedUw8JWBLvWWb890JA18nsnr2NBtmo7/FYilFXKh1nYQ4w+tYmtI
GM6nMW7Yd0C+pQYo0CzKJAJkkUJ23Uxxz6EASjrZpQm8y3Nd+z3cnc323LBBlO9C5QRrMk5diGZ4
8DJSz3LZYimqODbrDpI4xhUQRJu8KzkEO6HTXgH2kYifH/LZ8RYn71bdsHk776xAA2/wJlg5EZfI
X8ZDYcKf2S0sJ0vQZ82nqBsmf0d6bWP53ROQCHQRtSSkN/EjPFHZ/dlJPlDd6KIpgXajcvzceQJI
xv1kYC3jiGrhGhQPG+HGAUPxvFXchubs4deZeXxXrHlrhszu60CfhYomIwVjto2tmgwWdaXrjhsc
w8GV0wyl7EktoLz5I75uQ2rGvH/4jHGvtkxv7NA5jS+y374yiJU5mdDA6zCGSoPLvCowSZ/EjAgA
0t56AkZTpowsSarsenVam6fQfK2Eqm1n7i9SzB5MGgYcdzu3bazSxySOdJOtO53KlI14JCOFvDOX
IrHexMP0Lltx8ONBQX9CHqAFzkUxhXvsB7kUdD1MDpMjUHBkILEnXY9NgjGDioXLnX2CFJlPqfab
iI8YyjE3AavlvtbR6iHRgPcsazBBoQ95j+2V5INWle1Dz8ZAAqD+/mKhXDaVMlkib2R13VWNvhML
5lr21HiQv80r2xZbBC6Tf3cSAIRsJUqPjI4MKUkXxCmL1hHXrquXbPp4rfdzUJ0VUKuU7M8nM+9Z
s7TqufX7vJNWDbIGtkq80Rs4Pd/lbk0ogt3XIpdg3KFxqgV39dKvcNgBOCz9LjQ0AVxPhzIwX05w
Y4CCHDPcSa63QJ6+o3TQhKM554C/n5EKQKXitPIFAPuPqPEVX1zoSGxoGx0Kk2d/dkW4IiOuQt9W
PIiQv0BTvkXJSZjTyJKnejKhG4sxyqUsjTenAtBUHZEF2Te9qhgT80Tef0/jBKF2e8MTUtzyOCuB
n0yU5XRTXBucRGw8QT1yGysMK2AVmJpXNRxFOp2Io7xPFQ9R5vp96dR61On9ScNtqEuXXk+/ePpT
WHcPDWClNP4zfZoauYdO4meS2wsvo3DtNeJodPBWo1oomvyTPsAuu3sdXnd5d+DiigMESsLnuaCR
oR700ra6kYBCTiRd/5pWRqg8U40Cvzm38tjeEff/wSD64nytTAqA5U3N4CC42s9GP2Re3DUXJOj0
JrjM4oGAzZkbQ/bNgNBhkGMdXtwdGdeeZwb9IVWqGDlTo8r+5E1OT2PnIsmRSULTsJP3gBSnzCEQ
jT+cWWXTQ87LBbM6n9D0MiaRxGo5tuvV3vTebEIxES4NOpPIbea7Pp5Z0zJnRV4enD5+taEVQ6IT
xDcvtFgAbvC1aHuX2tKl9VDE2oXCCKmgLET+pjQLWX7Xprf1WMZQ/0DySM59iV0pwFzhMlN2WJw7
uMezec3puwID24i08Z1ZCSpWPcjEMwRS5y83KtPqn8Trvmt3T3WQC1Nhb+fbB1LVUpZZyxXemJpl
G/HmGHEKm/hzAqXnWzINboeSjq7IN6eP6LLsfDPP8x5KqdmYUj4h8AkcXdN7AbjD/LEU1t9G1y9x
S71WJiCFzMu1oZi4CoBx95HTgD0c7I3+u3ATIeOaehVxqybZZg84Dx9RIr0HI5mzOoLgenaH5OEP
R0EqF9y4jJDxredNSaX38qyQbY7l4tVzNNLM4AA1IvTHPnnCx7iu0RRdWvvFA/O1vdkDByKN8m4g
jseuaxyyorfZnO/pD7tZwJi40nbe091Y9esZgOBu7wjOWs9CQD5Qfgajn0WMokR2NNfu8DdXS6Am
ByHpTRaP99fdzrFGWojfso7Z72eg7eZS/u12MBZHMjfaLtrDJrpJv50gPovcYbl4hcDdPjUw3j2z
nKu24NEGSvGhBFuyk3/c6c7MKNVV27AU657EE6td478TZ16WjL08I7mHiN0b+qsZmRwC3Tqh2buJ
oHOZ0vp9rZd1hsenOVTSJaB7PsIJCg7We15KE+jaQ9PO54BmlstsgTp4GlMQ1LeS93d6YpUGBfPf
22BtIpMzVOlX7KBtjibfGtv8pc4sLgmH3i3+tyFk6vnNkAomvjgGiTuB633bsuZArVlwXHQrnh+a
4FZ7Ct3Yk5jyZNXLYLjPh8Z9w6Hk9p0b7FXstdZRgxGfdUa/U/D2S4zSX4UzvIYpIAw4bg8+riGJ
5NF5kw2qqtlz8x8DkWXbxzniZOBwry4p4cACJs/9sJfCpw6RKuGc7bpY6dDBcowx6BxKcRXGRN10
/r51wfUjsgU6B1qoQOvIdBixApUcuM80TQuMYIoUEHLdDypv8qa3effJUuPGaiGxOEbBbsAKxtFt
VZ5obhqak0RmqzucO51aEaOT1H9nXyvMVlKf9R3b8RvzgqHvwLKpKIv8NreY2c46wY3ILy0ULRuJ
/3lii6W3ZDDaSTsnYLsKw03OsZquL8MhvyFHPWt0vxoS08gjCgyGE0FD0wKGi4PitwWadefHSSda
DhvTSeLEZeKzYFBuwdcQqrS2ReGMwkYaxKOHvTgGI/t98r8bfAaMIgIWrU+lAhs1YJE9wveUfhqI
kMyAk5veJ0+sq4wdXVbyj3YucayPV2Pn+LU07Cq4xUDZ5labTSHJDXjQEUCUfFjMttBuwauqbH67
UyVa+HiebVeRGEL6pZKg6sUwGuQT2LWhISDYYgwiSdiECom+TpIi0Hqoy/lgcz/amgpxkJo/ogrS
7hYi8qLi3lTINn7QERRHdvXj79BpU5ZdTGcMrrZkqZoz58sKeYskb7g9DsiviNSc+NOzzfMwT2/g
DqzSPACy95m0MZA8KyUAhfkZjb/9ui6OwEFhewFwYIxgpk0tdLjPZYCu0iakLjTXDRwx7Sv5gxru
D1k7xBBKO3fj40THRjRrudgaXmP2zglv3GEobZIipejSDI9HX80iNlTHR3FxW4v6OOUd5bpfLu6g
edcigX4QNEOpEStDDkyp/F7bRuMV01ce+9G7R50+xQpT899l701dzHD6CFdQnIp1cBcxN95TJiW2
Oh9kHhuZ5nqN8tj4aCh/Bko8feD3028Aqxsz6FEjfxWtFMPSdlaWec8TC+zARR4S49Dv+HJ8AhKL
g2zH/emFvlJg/dkXYfREMVnS6FeFO8vFOjxvpthy00CO6al1IZjXzHV+8o332LJbfURAHZyOxG/T
0zW2lvxv6DFAFqYOV62eaujVOO+a9+/S41luGm5D5f0lOKAxW+/+6LAMlncNJr7gv617KaKBE0cf
3cvNUT2FUaxJw0d9w6hPtGOe9QRQA+ivn2qlXdMZmZUmC5Z/oH2A1zSli9JPx7qzsvAbP6xV8v3f
Uz46ELOpF17YoRzeYDlnOMRX1d6aKOXbZ3KTkfaahpgf9P6dCOTaFTcDMs1HieW1ppa55Eo6nq8q
bTAOBSf9WUzPH3yiUaQeL2TuGgqhjr2oGhr/WOB/3zahjOA19fTK4TFMDX+URKWEgv+17vXpfPE4
e+VCWjN9SPkSgI9g652ehYKYzHW01OnWMQujKDiK9r/rfVRwDkXhXxoqptZsHMTe8LVibta6X7qN
iy5jT7H109ly53KAUsgg1WYd+/nqwiR4NnfKjScR9xphYeeVxG9khEjzL4ZUmuvlg4SwDLbSxpoH
gcTnqcOKZLUSfL5LGbhOh1n84kB/C7AZEDRhH0WhKV05DBDmWPkMwtElrXexW/GTzaxM5KK2hfXw
IbXZNlj809Hr74t/9bCTNGSqGT8r5bGZIPyfxy7LAVXxKjbVEtLXfA8OIsHbUwWDFCWw0Oq9LT85
Ya1diW7ecrFhjCx5NqUgQ8iVNLadnUgV/g9LsH/BKkXWtTOYHf/Z9BKbaL9z9soorM4JeOwgW6+D
tiR+uA517sp78JzdT13bOPgw5TLRti16gCErxNVfHL+U8d2AL9QmeJ0LClb2J019hFnSFbgEOhI4
ohgN0jRPIQBeI3TVbapcMcjG1IdRGIBlaMYyuNYgxQVO0ktshcrFmey33yP1kg7KxwWzRLfQiqe8
RSNDVxW5IzPLwmX5znuuAOJ6v1MgCOfXwdEqFbPfFhYniDofFEeEqnzL8fUw3Z9WZu0JwybfJAHo
OYkbyEm+1dtAlFK5IZgtSxN2Yy1vZBF3bNLASTOyRALMuYqeUenekXooBi3IjoO+o40Zfiho2BRG
Pfb7uxS5BFRwAQXSEsrQzqOrfsjY3dGiQVvjEB1uD6YediUp2NX7L6iSZJ4XGF03eZHx6bv3shYC
q9893HH4/u/Bk6pwlzJA/MMl03P+Rzt0WX7LL+mK6S2aJqYrz3ZaxgMF6+bDANiNS/iF+pKvUeiz
W5gD9KkfruH01fNjqKSn9eiShC9M0IeYCDZkGF0DevcvgXoCWAQP6HuAUWHDz+zrxWvTw9b2Z/5p
I3v3ff8M0OjtQQTnDoJjba8N7Cc9SSnQqsxlR12gtH9hd6ohV9sMzLIedkHh7mJepx9H/Lp+3vOK
WRlYXSj1AaTP4MOkYW1yxSnObDgPz8g5ViT3wqM0TBzQfFddW8vdED1OPmiaKrIpOJYgZgaTuAQz
MKfjjEte2dw+xrgYh4pj9MreiJn74DDn2QurCaOZ3UKP0ASpopnA7M7ylyq1XU3u/qnv9ba04lC8
ft3TohB9nMaDgGTGKzNyILTT/Ao8XfckN3zYQ6Z7VrwEVeRxSLEmlu9jxa26b72Qj5X2GpIgw1fL
zRDkBmqTSCtXCgckJ3XANPWU0d0LyVzJcQWAAIKSae8OR86YkxVmpXDBIT1pzfGNaVVhb66jG2Em
zVSKl8J1T6CUU3MvtOmK8QjCJ2dY76ZEuq2PoxvbX3vEJsZ8DfW/Wp3xKS0DLmBlYT0zeOC3RL07
nc++3Pd6Skicht0McyfSxf7sUkVJP4gPKbIcWG8CATSlipi4v1VHrBbv7KcjYsAmTlT1yWnfPQ6y
i8YimHv5fDxOhhxFo+YYh8JA7yPbmKtA2eCScEzb+Xcnw0AvS7vG3zLB+0uhoN5fJtOkPH0ZCzqj
rsfXHqWAaIaecQtmcIsgH1sozLxQImnx57LFCA9Tlus925ZDEX5EVOS82X6Xr/i4kyhv0KJRby2V
bvs7bXD/GFHtFimQTKcWV59nvEUw621CLCQR4mr8xWZPFpRnmaCgMD+lB6/0PiCoXSMMG+4dRKVw
Xx6WDTiW3dMfxmDm94UVOdaaR7sLgrs+NM6IJ/tdSt/Md24Kq3gdd0dOXGjTa0UtfP90SFkJr4rC
9VT76tNCCNUyib4+dopkksuycbTHiijS3RgyIyczpTiEI5JLkQ7cyBFo0Wuf5Ve5mAtqaDiJ7/Ps
j/gJM+vZ1Jy5eAlq0zdVrReZwyjMovJkP2P2swsueJroVuU8qx0o6KUn0q/z+fluQ2csibPD6jlx
LQKuGy6PWT1D3DDcIPqxpHAEBodovrt3P+j0OURCO26G0YAMUDOQaq29a86dBl3sAI+I2Q3n0+Y9
G2vPCA4a+PLxZhf1bc8fNZiwTsZtqVBl8n3IdLaKY+OZC9umQfdUenoW39g4YS3KRgd0iTHV/dbS
fXs51BUVa32kTyTqnNiMBrR3iVT+guXPAaIjKDx+AKsLaxT2ZtgdNKYMUaqkPKFpE52Nl7jyMO9P
ZF9lwXOVldW6DJ7hViqsX5ZSiwGqPbcdSemF8B2xsWomnpt98WREW5mk+Knez8gmC7kpd1Oq2pT9
M4Nt5Vu7h2hRZIH170Ns9Y9QmZ3tf9Yx3gWwJtY94Mmf++zxIJV6jV+HicFhUYqthkhgdA20z6Gn
nvoMIEC1cWBez+rMFwyf7/3otdmGXaAwc1WOGcmWkHTL0wFuavnEaSc+5OZR3gsVCXaVhT1W3wAf
c43bWAu4YWJiJgCKzY2aakO6dhUSs9DeAojMjEsRtXAmdxrrnOsypVZH7NEjyLHJ9S3nQdWS8Kfq
4LfRZeIfoi8NR5HWy38UBooztbjLtws25GjDgb9DcARpCVnuDFQoCf6kwgOV3eZKWaXVjyrpPVPL
3q6f8rpwtZnTEgiovwrIGaNRjPp/iEfolD7VSOmFSW/Yjzg5U4cPwmHtMS6+Y8Y7hZ36wI+9h/BC
bj3BPV7S5SYxoH0ZntkUnI+lVypsM3jPLQW1pdkIFksI4d4o8X6TDNuFyed/hV/cZKrZs3RR/9cl
IhMvZ+swqYrhzVUjkwKk80lseKByZL5s3qsmhij6imxlDxbrFm7905abt6R5ypNQSsGFcc/BcbZu
eeKAhFQed/jvvODvcZ5CRB+Gm5YwCKfbYhTwS+jopP7P4XyPZ5HHtDOgOyfAnfTURjAPiSIgBp1Z
3WkN5u9RLbflQXbBEWxOQsmPs4CONRzjvTRB14azttQASWofVlOi9Ejp8QJksxYhlajnBOP/HZ9i
87vpqCSQZGyaHpMojpfzR4eV4Flo4SzfabpzoeEk6sDzx29chMEi7pwpUZOZLBlie0JF+FM2GE5Z
9a0z+K/cH7vo/cW2v52+u42rH57jqjt5s7TfpnJkUY4AinAPWClyBbTKDRJbx9WUF2wCNoYCUyqo
Ohl3l89yaaIPJv6ICveaHwXpowjr9sowNT8a/+pMiBCr8i8ISFDvTefAXV56QoGyKuTZ6cUzTVp+
RtMfXh6T6XTzmHoqnl36l6HDkj4zVi6CT8H3JazOHhncHx5KscXDN2BFJzMxflfmcg2ZicHpHe2B
rG5Lp0ydXCjV80QyibWB7yejlbEgRWZLLRcvcEqMwbNeGCxW+yvG/O+mWEhUoPM0jNDxIAE/uz69
oAxzlux6bBs5r++eAuLq9ApeLu+B4CYgemA3hPJzARqOKZBRX5iYErcviZkO/YupOvOqzGrni4Vz
IUZENo054ykSFCnas/0jkxh2BMNUlVt3ktBxg0sqbtYwffsutBnt89QmNGb3eZFum/Nj4iCUfD7P
GEnN+m5ojpVK5REP05YWi8GeqN6rTiygqcuW7ILjjgW8LwWUmF31Dtx3Dhbm2T4UGUJEpGkSTfA4
nEXfFbyF/4N+VFs42/Dg85fXPOijG2lpKFYzLel3mNhqTVtULBmKsQew/FvqgGqi143HbI9ujyw4
0U/1DBsYoIQyPJv2UmPOMgbW1evlKSCnKp9MmxDrpOvzWBe9U1akLlW3n33t2FgoFkbl+YQkYexP
5NFIZ5U75EC0aNohwYegYE4taInNH3CqpcN96heZo8FgWrqq9WU79NqAM5SqY6zu5GaJ3pFuJ2OP
7ojpx7oIJYotxFXKJZIoeMR6G+FVSjaOsrxUJf5Rzp/qa7/719BJ2Ve/qlyce547J3Q+mGbztx8F
eVgGKHsctzTbqS4qNOYXsrc2Q3QMKlzPaycB+KtjjMntZtsiJddD2E/Db13GPb9b+lY2klizEdZp
ip6yUH+LEWjx55kv85WmlrxpMDXo6C8na+Fw/rqHBIIH0pmX9JXHVQ6gbwco2IOgAC2Oyf+hvNzb
EB2v7/XC2sO2qIRbFr32Ev5rR4SE1lw7eEHHesLsVi4NraMbeCY7cZhb8b6rkrsQ8saxG6Xknfsz
NVgj7Ir/DGrrbxD19dVbZShPN/55waNJZFvzCwX54oVR0V0j3WLqFkNKFOPmrW/Pei/Lb6YjmanE
3vxSkr7siHlbyQL8Lu2m4Mj5Xq+ZTZ4ePhd03nw/OWlGIUnHBZ0WNUa6FTlpBQIEWoFEOa8FNT1Q
Zr/TiJJMAtBfxL9ZIjvkww1d3hYzgm9PKE3ltaJwH62vvStRZrVlyfgcOc1/ZFBRwuYE0/JblYaI
u45jGOcBLlkdPCMjDIomnLAXZ9UlIy9fbNu5zPO0EcxeKwiXLeifChoCG2AmEJQ2FLCwXOXxIlyT
8AXNLQ4jsyw1+q6wFuHxNJOwMPa1DbnX0c/rwP38thQncirJ2cSa6v6AIwdl1G01u2VtqdlCCWzS
wwZvDJ7TEEGMQNCSa8n9z7RmmlF9fQcY7z4CvGDZuwpaAk8qUzCePNNb3OogMxJjgMuf1x2MHdOa
GjuizDiP13diV7fGSsTUnyrUBWs8eEHEsVGBbQ7FPpTx1e2YF9LppQir8Sh8sr+BsOJSbjUzsiNN
X1Uufg02UM27jSP1j9PezfBk4vZ6Cx2g2AhsteRRixLutI3OLkqKKRd3/98XuJU4I4DH3dgRLaHA
F58yn4igj21g3my2CtMnVeD0jTnPije9aVRmKdvgnt0qOdta+x3rDsqPFjJE1q3KfUNJmoasbCeb
A6eXweBXlvkfW/4zysopNGTFHFtobIKorItiIgdhdOzU3de0NmEuZoWif+O6WmwmBYlN+fuAnWPj
N9QaB359c7qGb4kEDSp9GsuCG2xvVVIRRa/Wwn7B6lknfd8QSuJtgllGGQSP3gIZpA83wx/bhxxK
QVbACfkNL1/x7BDN9JJFrbEzhKrgNozFlL8jJOaOQQ5CeL0WCRjlSxoNx8LrFRdg0Z3LjQwsDEXx
ZMKpMF6YLyKYSvkBMQObcml68Mvp1jPQ4rYLLQrH146m1kaalQSybif7U7est2JBuDaPfgRSQNgb
uRlKP2gsO0h5ZOtSQS78aHyqZCJqGVdNPKI06ZKGARmsdsR6L252Yl8yfWVMTwmzSPPMLm/DZHhC
fXJ5n4LwMHuqiNaaTqxrwlWW5c6Vi1hhQ9AvEDM018WIRkClC1ZJ7XV5hC513/lbMA1iV6EKs582
2t2rEu57roeMLY1sCVhQap5e17/+u/gmU23YmzW0azDdy1nZSnrTgTo9YVkt0Z6bBxDRRBAANWd2
wm5vhaF/n96FDyCPYDgd6RY/gD4VTsKGyGe+8giIKuycEQR/Q7DNFEpJ8/T2OWz2d9mCsN9UYYO/
TD/8nAn7znLhwDqzWwwIHjMbKlibIVfEpjOOLluPGyoVxMOCwtFCCJ0WFzNrhQxv+A1Bp7x88zjj
ch67HDA1hesZYI77xxc3TJK6gW3RJh6884IgI2f3X4dZimZbHJvkF0amddqB+M3fVfM7qdRQFaXh
JlmEClva6cBkvgfi6mV0RCsePn0B054a9JMMK8INEdMfvlVbISLsDkBMQ3RZjtiIbtQ1qaCVmVaa
cur+rtwHY72uHf0fbTHRSSiOK2hQlnIWuhK8Wi3kDkRt27lTS39AQ2VSnjW9lGtNZWIGzayhNM/J
urvROwdHVDFgK9QM9lT8WjP/ftuQev+HPMLn8T9/BF6LZ10WCWp1MDJHaI6ZvAd6CqAd36Y5//BA
wXHrA3KF69i0nDXDGRapBdiH7EMORdsPr5kDY3D+sWIG1FI8RSTJRrCOmAzr1E5YjqgXxIfmi+AP
6IgQL24G0r87T6DvdCnf7GWvt8eRp8nExzR7v+z5fI/VulI/kG2IMv0ywom4STDWweWnOdLSbTJp
tzPGmyMtcP+om3NqpKC/0AaIzL84gZjADQqhQi2O3k9aIA1TvMVdQfoUbzCW3puN/hVNlAcWUfX8
T915UTc4/cJzOB8WKVjP5Ua9eIqZQP4DWKrKR6nTS/oHOT0I2BX/iYV/5YYZFCCX8O/ekICRsQFK
MOXqpUmfXs9LtqNPVQELpsOwU79bnlDyUMqDN3F6M1SnbRXcOfBSeVpCc/wde57A5ZSAtXUs5EK7
C4oBPX0Uhc2dZcg2c4wFC5jjKlHjekruW5I9Tg5zXPXdru61KpFtCBhtw0QaCKj+Ond/SDGFFn8U
dx+ZCcWw/o6Uu0JXQjoxanFOQ7zPfC1ImlfFLCscdcEd8APhtK+uWMRxRrYPxzCOeKO884Enxi7S
m2ViszNM6aLo5pYi9rMblDZjcgTKFShtf5B9X5eYqiD01B8s5VTnepgHbpeKVQo7yDg6f2ORFScP
9wlf+e/rIWfvl8jUqmPT5cHYs3xWKnv06D3s4xeZIeJajEcXVPFHgWGBCe451yVT0dBvTTuViQOl
7kcYEmGd9BsVwKEgzKxKQQ972kVSmv0ROc0mnVLR8+Mhd8GRc9seDiuEGiYZqL4h5NUSrD2twKdP
4MICuD8XPsoiuUrrMvrVvtnF5aeLCPmLvi85iphe64/VieBVUt3FrYjLk0SFiy5I7i7WztQklp5l
86TD3WAXNbd2hg3Umn6HaGN2rFFoGeishpV/rfs5JLshkSgcgHVDFk70/CCjdMc2XFIm3rzYOjUJ
F12hHe3FTEACyDpKpUrSecGKwd0ciGQYs0NCWor4xi+xLDZ/WT7Er48NSVrxZGqMzHgkQ0WpYMo7
FVQXtlgRNpx5PgumznUH5vu+gLTZO4uwxxuxGCm5Yy5BEaFxt+Vg1oVDwuLYr4olucoyq9odA+EH
IqyAvFmdkzBPGieY7lBsllOzY8fQOKm1ZGA0kfU3oaM0b+HMOXS+fhDuIygi5ugx5HPIG4KiWmNw
vcmJQuxOve8+S6yhDlEusj2X8tEnd1G7RpxCJ2JZA6Bgr5p9DtiRIQmAJG4v8i7Y4IEQp9cg6lXd
03PTc0VQFBhTHYj0zVcZOve+J7NPoMElRRRDcM+D16pm8fU7SGHVsl3XDbR7ebNenEDBOjD6Vc1f
IKlSqu6sEIHMr+JZ+/xDXG8XPjL6QeVPQFp15TJ2kJwh9Co+X+LHrDMOC7Ej8+VOlyzvZ+UEcGtY
sQ5vBhD9+jV6oNQtOYJj+V7RJ11m7dALSLtdkScCnAB4M/agV5ABIIYLWwPPFyRbGZF8kv0QweRA
+kGETC57S/9QT4UMsmJWv/aieYUSOLZyOgNu1P5VTjG5uu/FBiHz8fjZSgIEAz0SUTa5GKKNJmJU
nlXl9lusxQZcf6/9asJSdtDSsMjmI9sjAM6AL57estGDEkCZQgTiEbIoJs2VburBP68tmhmSzPfH
UwQXlKFptuwHBiSBTk+/a44i/C9GFpX4iNp+q55pCyA7Wifm3zOhMowtRLeeBn1woezFsP4l2sjy
DaHbwySrf10XxM4+A33M0mKtPDgTT4Hjnhm9sfiTi4/J3dU6NgCmGo7krKygadZ0VECT7WfwCP6j
qUcWxQP9uANMAUw/+50fx36BG/1tmLLcG7X7+9D4Rim2krcQTAzrE7img+0eyPidpS+JFBHcNiY7
c3C4fQh9yccxSR2LOj4wUAefvUJjnTjvnJ6S3+B2rcqaoOT9B2LGZGQxF/94iJOsIL/xgSRPl7tw
SNxWIGplGN4Mlw1MkE1lnZOp2R8+xfvSaLcW1BQkmBfFrR/fvL2DNNl688eVOo/y/luBRufRx5+P
/FU4ae33smoRS+tV77NSICChAfMGz7OAuSQeDttJ/0xs/fQb81K0nuZ5zcmqMLMyvqWXDF8HSIt8
ly6XkJ642Luq4LFqT4tWmcKvMGg6HhcLRDbBikWmcnRUYtwJn96UPEDXmZOMz73jO3f5FN5zrEUU
AXOUAzNKc9PY2vtV2fRjdOWmqZKne2DMg4iEOMyg3b6mqf4raXT+mWITwr17r1CmlIVB0R0Shq/Y
ojsUyYldmrlLm7PvN8PcJh2jUsG4lx1YwqpHDHGCmVRoVL6V0xNKOfL7TD4q/QREDnJp1P0srYPX
o8a3mE30ewBJxSLITpSpOxYlqC+2dN5/9rUcCRf4L4SskjhrWZmQnZUUEj39W5oE2C9ugqrDMDl/
nkiXtk0Uk4f+v8b3gnnyobduABWhRUVkrPUtLNQ5mRZinY3csuyVuxlkQM82QSqc6/kcVhu2JjKM
hz0MvjN0i0hrEi0ZNIaAODBF0MQlxq0KCR9gjO8pA6PZo0fQyrKsPDUGB4CgwBDYMKjSk++K2MXw
VT9vfJwplasQAH9wmuqQcvjBlQYf8F4B7Gx5iyulxD3VFSWzgiw9hzKH499nDUs1VdraX3qCGO6m
RPDPPMC1mc01M/fXxl85TycqQKBBiRVY7AOeaOOdZC6G0PwiSoODGgWn3OG/dCZNblaVEiWOsgXl
FUhyrtSF12Zyn/ADhtAncbT5ODkNcwfcVWZI+gf/5tUArcf0mbpyH4hZdsGA271hqe335+XvjbAj
f0Y1cA05R1x1oG/XuEHitgI5BwtfVJQAyZDMXOcJlqV8aUX1MDpbW7me2cxfm/8Y3S1u0btTv9lC
bily2HbWgpAg1QGJWgiZPAnNJKj80uBeDNAOm6SCItBihZwSn3+TsVeGJb6Xl9uBC8ODQ4ScwLAr
wyOY+mV9ZgUxuuX8qXn/t8bcWPRLv5BmNbR7x3KNBZRAR9eeGn/UAxbFb1Ec9fTmwOcqUG6zceI2
1u4g5aX8TF02Z/D9AT79qzDrYNZigSKFwq+ISSIHWjNEG/Gvt/maTTOdA9Lb2uy/jQjLMjfjVA7a
NHvWAeeln+T03uzqcBrTmqSRGUQSx0LU1th1cHjJBczpAUzpdZQSosYuIjPTAUulKdKAwjKp3ACZ
a1+KsKxVl0nETmJqkB2A639JDI+0Qrd9fUJQCC8C2HE7pT91H4WjpIu3uM9K4Y/JauGBTzIdTg6j
F/3BWvHDr2YAP01pq7mp94fWUixS5maJpDfvujq1ZX+KjY+FiyKOj3zus9cCsKyboZOpGFsZ7Ssm
kU8y+HlUavcoBoXFUdpByFqcE/Jr584J/QuyAX0JtHsPD3RpHYirxNvEwkyyVvHTztFbnfU3ZwW3
mCfZEsiDmuyHLtjrUWTBnKOpE/MbiEkgIIEZFoXIfY2nGAu7oguH7En/trvLo44P63Cu9ZknJ0SQ
UZI7iaY7Z2E+ppU7QbKn1vtbVUShFQUt33EXbAx/gDUizvbpgII2Tp57mk5DeXGDgKrhm4jCeWlX
GkvraQcT5+UinefduSSheMWQukuS28Si/DgJG0YMViqRS31gVu/okNnK/Rm+y7zC6oO9pBpRjtLm
kP7TWMrZSHufLR1A5w3E4pUd3FnXnLevHMHnR1WAY0Ii0HWkZ8tUiyg2L9BGVwZFmAppp5nBtlru
DTR5Af9X6vFoyo/6EDHo2+oP43i8vT6TeWSkbMfzOfH3qWe5JBkpjcgBX23/xpfL0+WQ7lmCRXNT
9qf7wjE1lCJ8ceaIlti4IS5sOQqyNRDo/A9gyEvaaHys5YZxipcSv39G3TdDjj4hYwZMb9l70fMI
b+8gSgYAWKa6dTIPqd4a5fgcjG4FBCPLtX99G6/bxq25HpS9GaNzUhrji3HjFDe5WRVSUn/YEva2
CYszFfdMO3I5Uy8HtPBkjXQ2RWHA6noarPipm5PcUSAz8GEoFbovhLhfUMOnJhmGA/14gvghXawX
kY90KKhrt98xK11046KTEwDDWiAs3+VyulUkaVWsYNM/Oq6tj9b9UJUfyt1IUm0OybguYVe1IcFQ
guUAHgRj1zSfkrSMD+hmMV7fyKEKqf2sK5O96tMPfKSag//v2webVLDJ7+DiilV6f1Z2chB8uXqW
2ZgNPGk3H2dw6mRjf5OnAhB1xSdHemT05lBRjWLpDpk91efjszbijhXHylYudL/zXcQwSSpFhNqQ
nJRanhbVskr5mMd20gJ6tQiScRA+fSs+O9f23msFYMykPKDCAFsxiD4qMyNy2UbQEFVmRyBpGnat
+Ybpt+CTba6bq8tFyuzqUHeN9Du/xDyNDiqsW5J5zV/UM0P4ED2/I6+q1w/l0F8D1z8zqZKWZocQ
nAd8QRIruwDn+FRH8f1N/BpJyML/NVb7H7M4lB75v16CZG1SstI5YvF6cYPXsaW+ZN2Q6p8ARMmp
zUop+S0OjJtK8sqMywbjZUyLrSgMpnZJaJyKRAYiSXyYbo2+qK/6EnjzoV4LsT7RREsdTBbvf2zL
exE+4Ko4UYs02TnJQjlmGNI650ilyxJJUPr9volpKtU6ts0IQSgHMWBWCv945tbWBppSB3yaadTl
JdQ58loJdObjG93Kg7pQvb8paFYsBNWUEB+jRdn/lJS2t66go1iGX1KMbRgt8i5nsS5LoJz32ppd
6JC3Bf9SRiPMa15SntzPSC+CrfR3tLxKr5iN6H48xr/rqPbv+nehOMvp8ATO638MQIi+ekqi5wI1
fLHoHL1gD3fjCmBCkLr0ol4w4h+Nidj/nFPz4Z9a9FZblYlTA2k+4sI6g/dHkZsOmVAR/apf+CS4
PTmiTOMEq7HTzcqdeDqVzu01iiOm58Ki8GR0jnvOLcqaeFiDKcMCyJeXbo6mkp/5esN46Hr9stiX
gvM1fwxcVFCFaic9i20z7Oit3tsBR+c4BJrG1N3tm78nYji53MM1DKxp4dwWlASQK4x6gQGxKMfg
6f0LZj7NRONgpD2hwe/aFkMfPa6JUOy0rPi+KUFcEiccHYJ0m5OS0SuOyAHjdpRmR1N6opiShmIm
B1CbP498y/Wnc1KQnJkAm7U69gIiTRMV/2HBPGBeZ9PzcTOfl8AWXFOR1AoTk8EMSuIxTvrRakzk
plc8yrioX2WwmPwKXusAQRMO/MoFwb9CXFxbtKx16VuRuGEBBWmPC9jNJzdb5FdDw7CFD98M+Bg3
INw5666T7pAXDbArGuLAdW0p3sj6JubB/s8vzQ230zvsQatPcWc0txRlNXzbS2BaJQHo94PkYPH9
6Z6iVyMcxwAcFNKo7gXHZk3ZIv2KpsWS0uzJ4L3VePN1WLi9RY9pzWZ5o0+lrFgKG/jgborRsLvU
WiYfm/sSwfJhg7gyCbE1X4hQgmyTxfvvEKbk6OaVRD9rzZ1AsEAsgAbiRThOFrcEieG0Yi9EkH0a
61RoIXi7xiDEObJa2nGJwcaV8f931g7PMej+HqDKg6f/BLla3Zh6gXwXqAD1vKyDVmMLgjO8drsC
LArIOCDoB2y6dmJNOhf1NYKxBiFbYWuTP0iEMqAqDPHNdXBPWGJq0LTLeVzWngJqoQe/CIdWirWO
BmQxjvU/Vk83paSc7FBNz6Qwzq4qYBDAwwrAYr0XGTqjQ20l0I5N8qRN7EzfEQhcwTWXMyCTeWGf
Oxq01qBkXnMdeMsjfCsrcYZTOAcT/VJTBADBDKHZFxDFko27mp67JRQc8B+zIWIX0Q6R87+wTxK/
GT6m5dRN0VjhN3BPEdzykmeFVRCLKMv8/YBz/T7c/wvA683m1/uXrsxwvlv1nG1hSH1zjRlAStwn
HFneLdAIr/rZl/CM56MbCrjvVfUj96RTtLaUjdfm36Ytsv3wBrd5POinvCb3SJ0I03eSM1MThu3j
y7Val65Za94/O6AquZWf0P313LjQiDH2KpzJnGoFioXJeTrT2iwcYnMsE7qV3wMTJv6VAOBslkRF
FgesyQvmqEMdesflK8NTBnJ5OQknSE7DXBzo92SZHdijwGbx/z9BZRUSoQsREJAXQfIj8URxSUde
3HwpqQRJIVpntmJ9HJ0sLalA30K+y6m5e9KwNDnqarUVo/d3Il29n9uZA7fao89AMQiWU2/ByeP2
Cmi9X06iucH0aJILignnZcq8BtoK8aYEcTMOucPW2poB/xtputpyShq3BO6oWeU9zthi2Wd0Tt3m
K1eLf29Gio8wg16XOY8/7Y2f8v2I11Fl3qRPi0q0n3Pr8zI+nrQa3hPlEO31UfNFrISThz1tew6l
PBRZgL64vMWtaIu/01BRytlADokvLlgGlsUXLkPwD6etyQSXF20xzIc/5/rLqXepiSV9xmL7P1y2
6+qO4zJcuCTFhRbvCEywFULegOJEQF8FFHJkuMhcAuyaF4rEz8ltekvznvuN9NgQzDT4K8QS9XQ/
GDGIVH4T8kYSIrVJJVBTugSIjQw1/xJYL/FjeXJO6bFCP0chFjIMM6Z2KWMZdH6ssYToNcm6C6Hm
Oh/dyMYIXTWgHVjviDtPK6mE6mzmtyNBlKlFGMA46MyQzeIgYWzLDoKXUsMhJ1ZO+p18H5JF5DLm
Rdo3c/gHVbTl9BetsuMgyUqW3lyhWc8gvB5Ob3oWLipy2NCgYqJqZshYRUBbx8KGG6whITwYUiGZ
IqHKBK+w9C9sWlO6edGeV5nJanD0lBNMudIsjxI+CpgCLu3Nlca866q61HQLRPcTaamR9JKIESYY
c14x0xFU6sT5dOV/ZpXZeWssJxurDLArRz9oBDzeHqTSzKWhBo9/UrNEuXg5ugfiLv+LtfGydjjg
2k9djHOiKMW4LD0bIlURQHx+Uud19lKr6wIkF/lg8+V3mOqFEZiLgJw2GWs1H/iyUlUBC0ARYT5F
mvSRb7Nl/iMY8AXqXTFwXgTm95i4risAIyKK17gTK7v1kBa7b4uT+g2q3bVym8ixP/+X8UAa+XLg
lR/ya/6Qy4qVBiG2y/2uSJ0S8o8TXI74QDtrpn+mTjADCdGVIdegt1XPIA4BASQ5QyBFqKRr/u+R
JFs4JmLWXemwd/UmLDLboYhtb0Ui7mMLi2z5aC+w0HOtnbJT9ky3FbvhCeYSMSffxFTUghDoqhzP
YRlWejHvLzZ0+O2XFTYJRZrv1tkGMUFXEntrJzTuohatrdDiyNoHb0/Lauopd5RVYDT/zHOpyvKR
OPsOGK64d3dtQFnQTtlPKUsK2fTzN/x+Y22dbzrmNixRSuYF07YQYjJlA36j6uSaRR1teZAPoILd
QrPlRKVGtAJW2F09foj1lgw+SEGW+EIOee+kEq+kFEarMIbYgfwYc1W8WM8SfVfJABPSylqi4D0e
zZ3K0cebLLtEAuxy+2Nl9ztDFq0WNeCeF2YhFXXjiAOzLa04KhxAYORXW5kSPVLoZfz/3qqqwA2o
i4HZyOk2l/Y/OQhEEo5V5z+CYcWYerKfRu1NU1K/zzxW6U3VVuO/DoqSS+9voPxBhzu2WfKTij7d
Efvk1STdTfyi34Cj5yzEgN0lwYd07H9hDdk2wZ5UqrVME9d5B30aqxUsaKyFsVOb+tSaTNB8gnVx
GJGQlCXU6pzsk+f0BkwSzPbIn9EO2ppNjOFw4qqOFoWGwY/LI6bBd3jTzqAqQb87LE9A3OnRAPfy
XszY+GMXNGImEV9u2kPX/yQkIZpISKNmadsbzil0epFhsJIwhLR/JWUibOJLDeYx+yX8l2SC7esz
1bn9aOLH9dSMusvifQCGIyPSuKuOm1pOsQ7SEIm5oLVv3YoAWz3SOiPUuYDb7fKKuOGE+gvo3Z1N
Tuud19tYuE6O1TXB0nz/xPSK5gXcHgFNmV75VQexpkHCQrSh12uha10k1ih73hJ8XSMqWS6HCujJ
jqi8fVXkbjox3wmx5/83SjPXEDGMeMDbCp+PF6mmUPB0fkZxsiLPkj5sgSqvLIHbsSP4FzIrfUKz
kwixPWPtweWLtkN0T210Gfmj8ah2xYQsM1UEA0hwoV9nZ4UnZoaySRGaSBw8DGMRs84gj6dtYsnS
KnrBshFPnyS4kOZDuuMDGaz4I40HdZehkN6nHG29Adpji2yQtBWoER//POI/VOWHFCAA3Q9X+cPU
4sg8HDvFFCuU398sGq6kD1sqA88aKDW4/7uWc4Txl8PzGY2eljfr23XEDH7+9rxGBqOn2XsBvT8v
gb+/dZQkxzW7yug9epkVmigq4RtlVS52kjugC75K3atY17s0GsvxXvI8gklPae2f7IuAWJAUQWPM
i3B19II0dKAb5L46cA57CzI0LOm2xCr21oV4A+oOlpfRwsTFXyolInMNSRv/kgEcYdAacyI/NuVs
R9jC+6u9f8lXYjtHv8DCaVBzGMR1x1PZIbgBWaQy3G2V8jliYE5ff8Js7U5P0ZXi2u0tJ1DjBEb/
OpHyCcU5TvEA/DQO3VSWFjZVjKIYcKwOrIBCZdXdNgE7m7HnGlHv+JNDtW3l55/AJ1X0UKdt3POM
vF2DVwIVC8PBl0aN+AN6Pym1OE086C6k3DZOq6JqOkjB95YlnkSqMFmpgPyluF6uhgDKv9GSGweU
MNECwrVAjbKk0OR9gttqOKg9fFxIe+t8IELKONCVXsnp1cD7XCiWVGJmfegGN52d24vTlAyrcsMm
bbOACKQrKpwEOeAcAVCVttSniNohHnnjjeTuhA1Yo4KLBXdCbu+TZyHG10oiWnSoiuNQ6WmsTt0e
8/62WNH4Vc67M+PcuKn2MwlzM4n69Phd6iz8vFCK5KB0zpKTpSJSrAotrcPjj/z8Pm8JXE0xV7XV
6Kb8EU8LFMQUAhd1Am2Uz6SjX2pqsqxQ43WsHa64NQzt3aReqyw1sAmnd/DzbQnUL4a2h6Wp1BQQ
lh9IDu7AgN1Tk9eghS8PedhJ+seSLghkRLv7Sc7sadnav++nD7XSGUOSTbDrH30FaD6hHn3GGCSI
4lh1bnE5Qe6HDsVuXQ1zcWNB9qCgpWwbGuxnW8QyMbRcNqQyes32xZreMnO1CQoM7mIf+R5NOy8i
YoOSnjKI8GLAc6dWzJVoP9kuU2wgMrhKsWFF1eNUd4LeVbf9InAsMy+hGpVktXzUFOQjUpd6ON0v
wU61uETLlg23BVOTE8itAVtQSltKOfaRhELz28LZte9+GB6Pm9FuxDzDWA8Go/Hh8S5IR82jrT+o
AMDQ8Q0GdQnL+E87HGFjmZ7HH0xb2giCAvssOeySiKZFe9duN1jjShgKJ8RFdVQj7+n2FYMVi3KD
JATzQ/ta5w2Oqj/68PbZJhVWYYTON5Ramg+UkWSnP0Bv6DDtnLyKiobG1vGHeNBWcPZpm7JyKr3X
JfmqyGKo4cXi8QN30/9ir0clyZvDg56tGJ7GTLlmxjA3XIZdsvxG1BfPqvgxHxvEi1NCzNJ1cggv
aZCOsR1D4TQ/R6LpTh1Qj0ZyxYt/JNR9C6fMO04DoZ8E/odBKDWzj2SfU+t6jUDSawA+R4cysVF9
iTRF+iHtx7kj1WH4h87jfjfgFVUDHsYzPwQhMDznnRX71GitTORTr/X6lFh4XyXdMZUNhMz/srnK
IMGJaRqtYGJwvRedGnnM5BHfU/55KCS00hZaOa193P4uKnEt98f7nKNsqHk9bc1wzkRj1V8SKnzL
tcYofdofv/f8tcgGSfQDboi2OdmsLqe6tn42JQk/atJ2USUy8bRR9Wdse3w9EWyP7IgX0UvtwRwf
pp6ds7owtIMJoomq3pwhLeSIG2ABPo+J/1EMt3ZprK/Sij3Sbwc7CHd4gjqJKt02g6GGT7rP1Ymq
VCzHLTglypM8Ytx4UDVpQ5zUIbvLnm4d0gWwt1Hjvfp1aeO2KtufSwbyJGfflX8xk6uXFaghCob+
9baEFRWS8KvNKdG4e3DlQGOOGZCzs6Vpl764dq2z3MDKrwNgo1UdrhiVYHV2Hmt7LXNO7KUq9Rq8
2EOfzO2MtvUS+1tTcY80RnNWnGwptJwzKyDUYycT2YMrtoKNcWIPVTCIMUQDyX7vzkAvj5O67bbv
PoyVAMvPVfGtkHds5YO7B2yBHnmQjf5UhPzo/tydYUg+l11QkbcybRlLyk9aw8ybGOs1KAXQW+hN
+y6n6wvxTP3XUOGykjScikbprxxl7KiE+aDZXmtwYW+f/vH97jUEgIRo+MdfjUByi4BIYZyTKS9F
uL0aMGcAbeZN4AIela0HMrv0uZEKzusyt+feUiHFtkpW6lfvO7ZS9s2GV7VLeHqAP1pcfWSAxo0g
qkJl8ncA+LgtZMick8nJfDQ3UcvFGBsMiwxK3c1v70yFeHDUmF4ZIz3hNW0xxQeKAPqjBKwzYQ7h
vC8Vtd9T52qiO3xFlVIfzn+4iBMx1G5I9RETHYd9cHL7QgN43qolmr6SUTb5MRK7bDi/xCqq7P/u
rYZYrdGyorMyeojbS3y/A6KhGXdMQzCineJXk2m5ErY7GhT9Kb3btZ8/SvC56oITloVFheB6R409
QKtRK1pKoTqrMkIigtj+84PyOKvWrRi/4FrWbSjhR2DdBf3/3OfNIvvxcsXwrDIImcJYNAmDcOK0
96WOptCMR5/jmoiKIbaXy3ssKePOjqR0u1vVkjTKJ1D99n3mSmrd28MK45GhCeHI5JrrQmBq6u5N
T7Ux3hFB5prxe/h50YSIbGCmAR+1HREnyitko2JMwXD587T/fce/pdm2NWDNT+CazQf5KzBv3i9W
1x2h9a3uGBAUh5y+d/8pikv5NwJ2MfbMNo0rMwplOMgw3KPyCY6Igb5ruwerET2cgzWp3dtii8RK
HK7fTlsmIRHP0nUzF4P1Jg9OJxilGT+aLqJoRX7KOPNDdK6wOkpMogMYN7V34UgTrUyH9EF0z1FN
muIHE042KdsORVfyveB1aYcrnwYOG9ypyttvc3R1O45shwVAgGoIjKmdGsTdAr6GcdOM5XAfHvRR
hm1GY1CNt2Sy4q3H4IjSDcupPymB9WDNaMHl/4f9sTwUK8LluDU7Q1ZwxdbVGxBL6CW2Ktv/3yNq
ln8EpiRfjTaY9ZhPqodQbZoLXhqcNyNw8kYpTY4ms/8xBVGQVPHA6H9/imE57XDuehN/cGp6TdSW
YTYvQGBcH2FW/Gyns8m7ShG0Gnlcxj7Mc5qZSgUQhffi1hRQPcAXU7Q0QTlIvqzQoLFyU3eg/QDX
+FJkh6W3TaTnP1uf2PdwDDWgVzmMQwFSkl0uSwQgPrpm5tLhlhanztsygBvqZOQJJuQaoP0d7UbP
zfCD/dIidd1BMPK3JSPpQnaVcuIGVfTibZ5ScMlWw4Xq1+f1AsgZ0UepBy96e9u/L67Ih21rNy7B
A8iYex870NmnKev51tYiG8LywPatqBFBaEpzVmIon4+Fyii/K+IOCJjUQdqDOpFxSHAw0014/zT5
fSGL3+Y2cWbjOgyXhzq4zu4NsWD/3w/cw+P8TF8+l+fj+hscRim7Qo0Qvt6PlkmbkzljKyqKPWsB
ug552VKD+VzVVG5IKKXHYcF0gXIIafMLXUj5XRYn4OK59YdCWV2AWmAHSAzRAFmyYatIpbh0grea
Dc/Jz8F2pc8oXUnhCOTQiAW/ktpQk2IeVh0ArnDSpKt9RI4VWDq/3Mx0BnLNH0ICXxWk1PB9Z83m
GCySZJIHSiZxJD8Fb4/JC0r2LPtgoe6hRhRETLl9p8uoY1YBGhgVPve7Rq3EKCl12c00OEGx/CXW
eLVNPKUjSaicsCsUXRYdLMQjny4XurX5zkXjjf5RgObKmpb2saNTCBo7WFvW5nlQZqf81tjKkcyd
vSJPWnBjB8GVTNy4DnTofbuqy2LUvdyCneC7OVXEOZ5HCvVVEYzdX1HiDvnNjZUSzvrAQwKlb2Ln
FRe6jZ3tR0QP4Hu7XNx4ks2IH2Z4KyoAvu3g5dHm73s/Vg9PUcpMPOXKw1VqoDYERieIikhGp3T6
FAZku7avPTgzjMji3Oesbp76swCDBI54vhEvuYlyyC6VZWa/sgN2e6TfF3G/AgSphOuQOAIQA7DU
ht52tZCqQpbCgcp5dwY2lQ/ex8m2jIIP/e9veo/E6dMxVxNDFOZywwpx0Sw1v2tS78/e3PzaxDsW
8sagbOvqb86tZenKtNPM51KWr3L/D7x15sXz3IcS2oE5rTK9pl/IChikW4syL8VTsOHbo3UbYmfs
Ljs9Z08i4oX8NEHG03jgs8e3xCb7ETrBQnhHXJ5hRyXKEC8K+VfuswIOPAb3g8yuNeeVicKfVn8k
Q02HOcB9aaY/7yqT4TLigqIClEHz+QOUdb/DuTNPy8p8l4ICPrx5+sNJdizifG2vqt3JMQ2OIVDA
oThlzvru8Z10rBtQ7ybldJXRpE3sx1OXAvkGukInJs7TJa6sO9WDUVXaShIzX0u4TWLtZfVq2dEn
iwFI/rFl+vlHueF2MRGATR0aXS7XrvPFmm2wqmYv906A0BzanFrhhmnrt61s8VwK+Jt6Symzmmw2
AdgMQClNGjN3d+Sk0HftpUiLNxjiXt2QzvnwNkEJyorN1kbJe7XkQSIPLHX+zvQwBCJDFkDh1n+U
vjEHVZ7Zo/EX137HQCdndIc3Xv8CrV+4vMIiJnxfT8E689lleBATZET3kKUqJpr6NgK53QOIDGur
eaxJVgOlJePpVNAP4XS9YMWAUbPxibAbu50dvUkgB0j07JPqdFYk1YwPPim6NxWtK08EMSL8vdHJ
IPi7QslfJbW1CbD3zBwd7NqZAQ2RakXOR/njIlcxqK4k6uGnVuNhhiiHI/kPkeTeBmjcygLPujZ2
d91LiHU2uaZmSRMlG7GSh+6HRgfxgOOgf3pbEPy39bC3fQUxoOFtSCOWV/nGCR+XMgOP+sC1kVQw
uKOd3emlaSvoXIXRpKD7Pguo8HZJa+AKx133v+IMX+nL6hcVgi3CCbmOdOJDcHf4k1adm/xs4eV7
eic3UVE1LOIgVc9arlftIGgWj816Cg59QY77YHUu86SNnKDXOxUbo4nSc6kezaaQDXutf1DT0jzA
cxIXGVOU5pepYJeWzkzh4IBTUQmOseYXDqPGVgVsesjwRiNnBOvnfGRFP2iVqj5E+lkt14VEc6cp
U9bBxPeSFKB+JxUuIE2MBCS3c+o4Wh7RnBjTUryu5eF1hcj2+e7D+L/8jXEbphlk3g5nh0TSzA5k
TQq+M2kkg5oOuntKAI2kooPavDwwNSxyBWeQ6gYFO4qUUkxbe6H4fXxf87ot+6cKAJ3MyVMkoO/9
gyNP9tdclcvjzw/xEpnZmUbrZWBie0hGridmD1H+MNWddB2hmfMwaVnCwRiPkB1YDCi8siQUshnp
KsISdA77yOWoQiaGG/yktCIJzj4KbmEr2b1GCBiSCHolJZN1Fw7B6O5GM6RXLwBKzcgRq3PazsfQ
m3fC4PsjxKdJzvBuP9wGwtbGHDar4u9IRf3+r4Q+P6Db8ibgv2nVt0cqkaAEe6+MMfVlf+INHSVL
le8spk23KWBUPBljBL0vjZpAwv2VTlDS+MhMXpPSz3C3iUeZdGXAZpWkYUlMwwWHfoHIV/lnjj9+
iEkYke7JvsaVTcJg589G3VdIHhLH7RnwrXAGY2FECZWRfBgnixGgwWob0bUd6g3w+sOBH/lNkZ9J
eEaDpAMtF0A6BZ4CPmT7fgMIZ9NE2IuXFEwFCjgH9SDnAPxzLbEvwIFWgPutk7pVXLuLfZYPgifa
PrZ3D6tqAQgyYGMQH+VAwoZjs2oblbtJFx+egPJDepOmnQoJz10QLL8EXW3loy06smR33DUyy1Ye
TE5ResJzp50A4pln7Rrs9lNjV8e3E0bIJZRP3DT8zwf4VoTl+dmk0+vR26QTV4Nw+wP+no/wx7YW
yUFYO2hyFK2ZonGI6d4q6z+SeekpxrO4GoCzfLbcjwwkJugkthY1mqAPmkFmPWhiVqhkDHT59u0b
JyVR2Gbf7fTaiZtfwxMbf/4MD1DD/F++o7AR98AjqzzdGbqbSX7W17t7TVnJUNJSuWL1vruWr86v
AjTCwchBXFSPXs0l9Hs47MjtmiATYGaE94nB5gadz3/SAAj/8yuYsE821D2LE3brxpkX4qr+Z5jS
vVWyTRwz8uefLT3pl2mr8fs5AyAvDbJ5rTlf87GAxOwQJfGGmigzWURi5nio2XDFx1b/qZDTjcbL
F7GMmzOqkhH4pbesvl+GqiJqLnCqzmNJWpX2tZO1z5GUuLI10Jq/RnnlsnfwDDq2miMn+BvpNAH0
5uZYxRisxySG+5/wQ+71Ut/SVbseesog2qDiFWJOQ2Bzro/cY17r/+/tchi6yKfPpJIdGYMxKzqs
qN7SDUIST2pvSWVesD1dWySHwdoLhRaaQwco8I2IY9ad2rOs3z7mJz00vqONe9jKST0Hed8iIRuc
m/hftWWhhxNcAwf0aReYXBbsnhxMjhMl13CrIJpBWKCMzyUGYxl9aiwk67ehniONJVBptGSrbs3C
AcSO9y6OZ02UFJaYtGo0gJZJCPUtG3vQiO7NgtDHeAhz6lvJgbfITx0CoLf5L5Gf9E3Tp+JNU+S0
baMMUtdQcPIkUw1fSf80OEmx+TnY6Vxn/MR+9EkRmflMj2BIUkPLCouBI1Xz1g/M5dhfxeCfg4sJ
xcdzX5AknS8dnlOiBQj9B0H9w3yDdpowD19BhupfkdfUFqliXH3FP36PbZfyx7fv9XHnZyufj0ww
/a7hP9aR/ctySxBuBtLB+QgN1SjZuIedrWN2iDr6RbU1Ui1G+iDx4czTUkMwk1syGyJCkOjho9r7
mY0kYqeGeZQbbqgfovFhZzKLd7RP6G0NK4F1/obFVu3YDc/NJOtcpmoQcqieVrLr6utwC6w0z902
zBdOg+EB6wTKLOobhc4LnBgElovqVQbWN3gmhuD31M4X7sPsXjPMr2hVzesqbBYi5xOctxnl5S9Q
afMUUyhJonZmbUer2j+wnU/yuX7YEEn0w/JM03GilwYmsWURDazdQDRp/jlEyiUiB32UUOPjhQn7
jG9peoOJwv/zW5YqzD8sobq2rl7VIIZ3FEpqN3XStCLknQT+bKmSkBpBveS2yXXXU4Z/rRA+Fa5w
yDcxukOIAmLyFc07ICOx8QuP/xKndVbBSJHKHwFnJQAtztAQNQdg78TDko19NcyesZjKB35TZEVR
PsWbKrl/IipfT6jtiG+Zryi+f/B/jlXEdtFIn9fEaL+l2T1GyOjM0lQQ87NhL6xTrxW0D4RnF8GG
azPIPKYOT5t3QAifwP0ZLRAyceIkXUFGrXo+zVRKrdiYREkEuxGXCzlGvIuulfVtk6nrDI+2/VOI
LWfJgCkcp5hHHvYuOpo2vo6A93kQIG4m6/+cDtfkhF4U3K0u3kf+uFPYfsJ8DRQve5wW+oCrmDrg
RD6c0uemlcEk1Os8tS8loZe1sArlkmfbt1ZemX2H4qnBr9mY5qELpEFOA1RM1Uq79YH/jlyLdMX+
x19uVGdeYxuUrNoR4N+47vZGHWxyutPg274Xy1EcjNDw2oa/GdjfcqfJxTWsVIelp8NVAz7o/Qrg
0GZwWNo8MA+L4XXpfOq2RfZh4xVMjYj3xcVkSvnXxBiXcPYyCVdfS6//TFOlNCecf/R803e0r5Kg
nbhxurKXqpBDDQc48LqF/hVT7HjemJJRnY9cL+yDx7X7zaGFYe4idGuvTKGrCV9aHXu+U+hWse7e
OgX16/jvVnjnMJiOa57ayZwpgepLmPhTnYsYHZWqKUhfXxh8Cu8GU/aE25WxiPh7apE931ogh8rc
wIbpCJa94y2waDIHyBeDPiQNSi1QYYnvhRY3q2+c/8+cHxfWZ9Q3F7HzPoHjMI2sDXNqG7eAOLB1
6O6HI7Hc81qdKQeA3lAzpfq8rYypZEEZpWNpEt3/4LmMokEvGA8pAlJO9jQbt027RDNfQNDZAi21
u3QXNWmibxu6rIUudxVORxTTtvigVvk/EMYs34SmnWGt9BN/9y0pTTAvvHsl/qcBhfiRJeDiikDi
zz5L47dNs+zX47DTQh4UA/EKE14gK5bndTirVaaNH+vyyJ8NIuTAa0CZRV2PF+sSbAwsQ4y6/ENP
e2WDz1k33EmI0Yp0WOgdASMg+GNA9Cn6vuRMB+bVkQ9Xo9p5cwLlvbjxJT6OunsY7yPjLlqOI4vu
vQH7Gt1xgMHHlqZSEcG2mbAOQfEpkuu3p0ImhVGpNR0y9KQcH2q57PMbf37ocOb/nfqU2ifkk2fX
Vy/7KSmA9sO8rWKo3FOMXJYYG3P5b1NveCGNCz1TlYQvbYxAtK9RltVSPNrzrJPYR4SOZrP9zX12
6FEtGTh2yqHJCY0gIukAL1Pa9a2EH1jldfkiQxPGsGD7ZomsjwS5zUH5ayzpU9DYezffV8Z9K37w
oniklTYTbDBd37dtu3sqj6eL2MnjDUeiW/SmZ0C9D1Snlllsgz6fZ+uFWm7reFzzGO1JXAYhMA1P
USSesyTD9K4TdsKJMEj4pew82EEeHb8PNSIw3o+W0Kyu1X2ITEXxZ2Qo2nIKAKB2WoAF/xgWu0jw
Y9BlWCdplcIjP8AbAq+XHZpjDISrWVMmkXp1gumLSOvwvetLpd3gD7h3AcRsZejeHj2MUE7nVQTN
XJ4e72T+MLZmU2ULg74lhCPTJFZo5pmGJx+Rq1OxQdPDKSySME8aZeCLuGq44hjISpgy6GcATQdU
hCvVLgS5b6hZmadwJm7fRh2Nd0474VGzqkKNoHXtR7FCNmlE/O7BBik3QcX5s21gmKHTu4aRKziu
+mSNB70sBMwYiGO2MvTNIR8NvDiFUPNoP3MBGwNRUzyPpr7sRpNE652UhPvcXqpjGC5A0WiI0lSK
AUwsJckQ5PM8qIU3HGyi0sGWOZ/p6f5XDHl2Kft7EokJBdcNtjwBaaMqvvlaVTKXywGHdXDV5QOU
MopC/X97eJkXLcjwRdPEXMV9TsjoYjcgrFMG7NrE9pNwb3vGS1WH4NBVcHV9bcup7M14xOCoHnHF
DtPLUAkJTT1OFtUBJCsKsCTgmiddHWd6V76vLH/TV6PmhuSD+JgjM9Gah5T2j7WmDPAWIPJt2oAA
Eck5cXoCHOf+jsoCP1Fg+ClbmS0CvQqN6AkrQrj661PeYKRHfTSwyY5PW/q9BCvCcqgaEOx0391h
bFt4qwiFd5Qu+eNMDj1/m+1YGPYLTbQ6znDJw6wqDgTmjmCHTHgylgwYhlCRMikATz3XhbZEpTmR
L1GVnaDERnaPHbB4u61BEoULnu4b+4c70O62KDTfSTYh8YT8eZYobELQgWU8TEDCTKn4fnUZHFr3
J1ltTocsvpoRoF0J88xlclsFeuQquMG8X3rk4lfZdKeXGmdyfNj3PqS96Vj/37JQ+yNRyzOM0H2y
Qo7mNGx+cBB02AAG5aKfmaLm2wHjvsBvhMRd/9zFzk8tD55zXIYThrOC3s3AuwRerioMvfUbY+L8
TdAIoCKmq4T9a+NelhQ2vmitJHwjoFbF2A0MYxv0HUuU7gXbjOeob/faq5ygUsEpkcTendtEQLeQ
94uWofbca4CGNBTRZVwe5D/HUB0Tpj2qvZLIzUryU3oxoKys//pxwHzfoeS9ZixLSp7WJTnnOH84
xYEN4UgL5HlusOynvYIwOmAlMUEnsBpoJtvLbmGAFpWBUSAqe7u3ZyMRl7y1kFaRCVF4HQTGIalm
eGPmApJYrUURSk0Q/IWlOoed4KAw5ztxlSQXSr3C1IRucAdJNDwrwFqU+JtLNDO3StuBBlmMdIXL
rFej8gRVnPdfKRzX8u3M6OSOrJn9hNepE04XSfIXHrkRGKPBcR0T8D9V6sw9T66WyJjmW5JtYZZz
SvLGEpcPXO8bW0+s5W4myswAWalgfuzhW9Czo9ulnC/dmxY4XXGxhRVQHPa1fFC/xSykSeYk122G
v8PIb8zqdN05ikmndtbBhjfRyPAzzK2aEz4L+YCLuByNFNtOtYBwpvnvuwjO0kfytNGrSihdm2Km
wcHKz34uIPFQ9crTKC3E4Lbe8v64YTwFOlXqrX8QXjDkd685cr4zHsEEwtPZDs3xSojaX9X/vipx
09zEuzRM0QxZD34kHoOJW056JnzUYSwe8CIFMeJpJYKO3dyuPl8DGN8S/QGSMsKGPC3nH8YUOooi
Vt9d3hMupCOQk73U0TrfM5Ood2PlygciiDnqACKXluUss5Cv29B8zhXix4hrIn6fGHHFkW2ZzNLs
SrtJxVAEeWdSAN4RUKJZq+4mcNR8bUNSASDwxHCIGi4OSA6Lai2U8Tklhr+Qs3INCnMnIHSzLL4u
wKb303OXvyNVwNdCsuSmL4SOP/d73ttXvCurrJNpp1trNKVM+YpcsfU3CIKKmQownRjgt12cF7bI
L8/i7RQK/jQHJjt0RBGeVztHpaLQ22ckkUS10jUvoS1ti+K0RRO9MMPz6A2VT+PRpaYhupGUMUsG
vMqR7nrrargUyJbJSEaKxLJz1OUItxw47Lwi4YVwhqgfYNPi5szuXyPc6fZZjI5HmjM/aQfmkdgm
6mFtyfXGzepXiPRcLc/rXN2Yog/rw9FhO7JgT0ZslHV8dJDliT+fIWPyqdf/RY3hNWjADo0kKXt+
OmnlGNEzxQkAE+3uADccxBJCPjSacnODZOYNaXR+/NdztXa6FPhEkfq3Xind8xj8SZPopgYvS+Rf
sa1/U2CdhcgGdx39jC0Qda8bwS+9hwdKgby0X0x6YRwOvWkgXgUgGuTKB+kWasMXkJxe77dFY6ma
UTk5rLB6g161yUSsAo/wVSo9XL2Pmd7Qj3LJXXSi8IORhNf8OWoOdtuORJj+IIGngpbtEWm+yL6+
NINjXwKyq/2CFvDGDcsqwU1KfJzJ72VOjhbXBKND67vtYtWVGuX1qUPrVVYUGzOwX2BqNUIG8krc
u+loE2c6JG11K/aoLzlX4guTn47lia8oV4T8Q6qAKNi68+p06I17nHRnZbnxP/sw9EqUZY8Cs3no
DbhvJel3gqjhO5mRlbCw5JRUnaz7g/ibpTBeMMweKFzbwJZdaJBeo+6h3n01Kh/Q5yAq31BUp87M
9KczKyVJeAjNehDIkUgd3jRQxl59lzDZ99Z3K37SmKHfGGReKxW7D1fsSezi73VcMGDHA+NuaSih
mfwMNaF10C77mzEs7hF2H4SCm4FMO217lQykTtJXy7vOnfwTaGcNx04g+yVGxcN0RM875KsixVJl
GosZ5EnhJRiUUBGKNrgp31SzjgcEdM9SasEjvyu4nPMMis4n4aV6zz2FIuXcrvWWAh24+8Are/8S
UlvwZ64FzULYKPrjSlxWSNbt6ouovcX6g5pA77aqon5VA2cMYX+QxxzkECyUwckd+qALng0pktQD
OyWovX7dd5sIxQH2aKLQeYjnD1GP4gD5D9GrIfbHoJhpKyAnUjF8YDnZxXyc8raLumPcxskvkjog
qpHMGtkdGtjqiGiYDNGnhA5jwy3nCwB26jruCNVm1+XwpX4gjPyuU+HsOsCxxvPE+n+je81EZ4kQ
PrvdjPN3J0rfVbkdlWr5Zws5cegDc1EUfDymuRQZjsUhBwfvOXUqJmklKSeQHBhnqFq8p0dFNVAr
y2515g5i1BzeJiPZCyXTptIxJmLF4/3PbQQ7uvtFEjkdVZqbx1sNOhZ3bayTKjsL5ZQsYfAwxCPb
XCzCfmCST48xvDC4/szFCoIbOhOth86AdLTnlnU86fO3ZV3dLsyxjEvBntQ43SYroSjeSHNZDKGK
1wKRoBMYtKRwme64roCKDbmIucoqEYMs/1Fkxikx79MSy9lfRLu788G0HG9vBAzMdYrEnL4i5C01
5MhmMsWlr7hIw7qIN2i8laz25BD+9ScaeooyfQEalsd9C++hS+5oN2HcTHg+12jzp2hmtbGS98Eb
zyspkQz69qSf3zLd6eDvaKzmjX8mZoBDefGmEnyW0pDT2+sW3mM0sm2o8u9VOm1+q8EQJ88TxilE
c03PBBOgcqUm0+wk+bPaH1h0lUiAL7aU7BQV2PewI8hSitkq0FFcOv9qL72AHlv7JbwZIJ8lozOy
zPKlMEv0i4PLOkZvOyt+EOPblEl7bZLYsA+fII+qvy0mQiJZTCmNYmB8Y2mAN9OoFZmJAM6q8zlh
JR87zrUmoI5eeY0ljjHz9GQF5UutVSA/f5HsITVRIGfJ76OyzDsV3SzBrFmO7hXiXY6yQFo6MYAa
RTRSEe8oq83vS0XkyQOxAi2fSjvQYdwqRhqiVWCnA/U83BB4jgy/iAm4Qefu9v5JhZ5duBZIgzrA
5kCOc9d7fV3EbXhiKi6sN3mcQqyPW0pD74rPTZzBWyUYdqyPvQ44JV1QvyJrWYNcBQu4JCyvABRE
ngoyTCHRH5XjRkYE9w6Qrgk4B124wHOglyl9i5qIPcAxo98QL5uT8G1oBP9Q/PHSGcA698graxTt
Mb+ZYMckta2cf7kketHVPIhqGNZXbVIV0LG/zmIxiSooxAwUrw22DykSM1qH3c/O8IOSpZzeHQXw
6aaeNJrv+4bPQUXpE3iSRIznikCav1OAOri/3O6bmeyE9yM4xX1riC1PKw0m1nZQqOHSz/OU9oq1
XvT8QMp5HkQdswh3r2WeY0CBn5QU4dqLZtH72K3D4J7hCP3p6fyhD91o56nuBlVLtjhYcqUJdjVW
4z6aAO4dfFrO/Uj2QtcbBVY0wc2yp+3KOc7tYtWfoeNV10ZhOClMThz1/VX4LH4QqPx+3f0EC6UG
nFLrEVtBcYzFE2liyrkXz0XTfN/391obMMT7b4CiI3DJh+Ck4Ng1+HIA4jsmN1xLGUdeFpLPRCHU
JPkrzltum9XRSs0hMn3EQ5LCZCOHqAcFpWG/v/fQ4Yl9SQe9e/o61mmpg2tzUkw+IvrWdyGi8sfG
N9iIc+IR28mZk/cOrL9sviM7RCgMZlXYOY+v8eR3tD3Pnmm3i0iGzAaqR9cpPfmp8t03Q4wAGrzz
NKA8AmHRCTqTDW9H7UOF9tN85WgKy+cfMUmy24se1peUFc8thGWUYwQtxZE/onqGY8OlHRrhcP0E
R4L7eQgsWwK7ZxkNC/BDJwTo7du7rO05sEMS1i0fEsl6YJL4O9u92R458j0oiRowgSRFdfXCRErp
s4GbZR3ni8mUmkUtodtRtogbOcxCRIbrIXQpdlQgYNUTvHxfO55Lv+0Kwj8Woba5ZXpPRHugMKIq
m3Em17gnq3EkTOU2Ssxf0q1QT3QThUhU1q4SiNaYDykIQsdzTpBsC+z7IO2ZGGkLf7R+tbG6NSPE
25GbP1pFFR+8aSIhCcrmK3V7LqvVSaRaueDUtLgjI3unfsHfstLZpYoruIeAU8vqdDdW7MAiFSiU
OKx28mtLD4l8tMJ1Hx428ua7NWpUhj7OQvD78aCqvq6+mmTIr0iHwpLwd0mIfyXlAtNx4J4m13Js
kUNcX1CC6EcI1XWFuhY7+O29IXalLn7kP9lVMKGXYHv4/X8986wcrHYlnrlLF2msUOgSnDxWlqEi
rSTdeATl4Stpd8szFEm6S/0839pOS/2b6CPUZhDURcFounE819d1ZCJHa8uYgR0TXefF6PQzSwoy
qu+B63WhX6GxG2W4TvJFe/+KPxfyCXPFfkxcedRIJFRrqljkOu0a9h4cftl427St9LUSt3JF9OX5
6du2RCLLdssaqnEwipbYPptfve/r4PYyXMrcdjVe7R3eZMiv03694zOTnTDzOM3yfxiYSUGZFCu2
yhnzqvOq8pPxFuib16LgMsbwTAOVWAT33cda+6Ynm9J2YBni/DVwEV1Eq0Xz3gQcdW6cToo97d8A
CI4z93PSx/07EjcJUdyA7rCQyFDijffm+YUa9MigDMUY+SmRFPBmyBu8Ba9xfvFzWtegnHVPNpC9
zmcldd9bkHgc3Cq8dufY4ucooCSyU+uLcg34RzaSFBrWdeLiOn498d5QnM4aNfBL0fHj4Xo+FPI/
kD6JmyRD6qW0uy1faWVfRXQLe7UNrT0AcBgyyBabAyn078Ksry5/zc0iS/ZLY9QOZtzFbEAsWW8f
OGYBiH10sQwCiNW6rJs9VS9Ly82o3aHZWGfx/yhtJR1rU022sT6i7vqMyBMkViaPnywff3ip58Rr
/Mo7lCa8z1WLXlUwHh+Rei7ZYrmM/8hxn9PHFdTBuPuTN+dmWUN0HXv+1Q9SeKI+H5iKKnZvw4c6
aukAeoVQYCm5408Gslp8Cgm1i36zjJEoAlkvjKl2Z4MNoz7ufwY3cQkOQsyOrOA5F8WvmBY0xbYx
cgFKujNKAjpqubhJPTBRsSKbbZkGKoQHezzyFhdngnvLDlJwi4L6yOPqom258l6wM48VovyJNJ/Y
JvVVs93p84rtzNSWUUQaYIpOC1bcWRjzJ1sjRIpmkSN8IfaVO6vEgd1zGIWRr+yS6zvCsyWYfZEy
Av/l2lghhWVgJf5tjQnlh/zGJZWi5X9ea+ZZLshGQm5my4gUzmqgXWgWWYeZSN56TdWydDYOnkHz
BzKtUYseoG4KqiK/wqKZ5WHLRJ9N/F2Uz6gxcrllPZGNIqDovZvY/uqmb7nI0Zs45rzuvenYk5IR
ALJWhp83x1TbYm4TzIgzOGf4A22OBfIiVyUkoesMHnJs/Od9+eU1LPBS6zGGMLGCpXngp2j9og0e
gDELOajcekrrRRBNsvqoBBzP+Dh2w11/2d8wiOu1oArYPKPw6qyVieZ5Bk87DJSLu1z1Z6y2TfRB
ofOlqyurczz65nYHFmYEjHW7kY1gYEwKVBHl92NX0E4EQdRasXZsNq3oXJbwB2URriRS394m4PWv
EeagvUVOw7t9L+zA8WyV+VCEcrgFqGYMAHCB7CuGKEdlSM97o11TjexQ21TukUbWxrScP7QwwdWd
UpeU6YHf/UJYwDmlACYhBBURLqVrpBJOwhvtITrU3gY0iwV7/UMMFJoeqIwVYzgPfLbotXlIDvYH
jj2EdzqEvOrwW72DFgT+Oxo6NvDiFdtRDq36xqz9VcMctko8Qyshi88Of03M5RSMElA96pEuVksq
yJdCjL4WL3Iw79XPvfGzCss1gYno9R/9NSRut8PDLKrYOh+9wLIWwrwFM/fF7m/BUJRgb9uG17y5
LDgwO56OVzxAG5gUK2oy2ZcSyCF+qKTQj4RAg4auPVckV+IkubwCmRpI8soZaOetjt27Qmb1WMY4
1YasueODGpP1PDBcKGPygT+qFy0NWgUwBoHPCrcoFNey5TMXeS3/8QcbDJS8ZdN85orq6SUJN1SQ
GoSEtPIKkK9X1eOhNnxUJndqgqfrOPuZlz2QiLuRgxGPZxtcydvdaWiSGewMEK0RuCmK3RM/dgZL
6mclfiyNoM/bu+otjcyXR26bWU6nLs0pk/7O80o8qpqJjPnobtigB45sf7IuHVCPotQ65Vd/iqKx
npQSyI+xwpOpaRpXlyj3ZOwlpIyf78nl3GNU8GFjvrihPpbMS/i19tZT7gUUerV8B427VGKOYQSN
bcZBaPImLrHaEsbpIYBTK0Yp12vk/qsPcH24V45n+63ZxxCpGdrUziYYC9zMpzKBSlA6UVpk8iwa
Ju8oekpuxAXOGwgUE6w0OIEYP3qQy8uW3yL1amGo4mhjPFbKSJSUeVahsXOlrgylJPrPt2sfa8Zp
COrb1rVOoEcmxVePNOgqzbNkGoI13bsZuJCzoxTUiDSOEvaThg8ym8FwgvZ1uG2xdc2eyCitkyKI
LQuOaR05L8Cej8qxQiLFdInQCEi3DNBJxVzYZ5bdmRRnmKlX1WQ5YachVcbCufOFy8fD6oxvuK6l
omdq6fYXC14qPDaiuhTjUnaUMdnWqereK9MP3mUNmCx4sPeKdQwREo6pOAYn7wpyf05eOgdGeNw4
CA363d7RKAHyOGbSznerLFtU/b4cIBTuMzqvI4sXDiZUmxpUji2TIzX6oean0xmDzPpNRp59QgBd
rPiRC94o+1/nbRUjtAnvQkSL92AzAy7K9J9avx36xrI7e0ekui+5SOyVHeHUlROptOXufXfFP6Aj
42uFL4JmD/54sL8i1yQAaW9plc/saQkslT3JVVrOp5OSF5nzI2p5HdFYChOtF1dmmowcjq9oDgFJ
gYR1UFBPJRaKqYvN0SuZFQ3+gVRcpQaj8F2vLIjBXS5k5l/rbMwcSQeIUReDwUqbFLAan+pL1Tsh
YXTrnlR3j6evubVDmJM/Ldg0v+/rSlEYDuTPmJvf3II9WqFfVCZA3L92cpYeV9TnrKmFMqZ3C+Jk
WGk4mH0//TPT0Mtl3NnGAAST8TRRFQesfRcyBKIZADh2vqFUX3zWT5Z4Mi3O9sTu4EzSjRZ6BM80
5wOXWhGCXk/8I0/xyWniG8jl4RuIhBfDmHyOzOwbCu/nKKpAWT6fOdt4zwLTcebw3YRWuP2oSTAL
xXNnRjtWm8E+Aoj6jmsE9jFB6IgbYg7ceqaMJDh3PLwFEmDQGzzAelBO5zI/7B3U+jnCOa93xOh/
DU3hZz/0aShQea+q7wFeLpYME67ks3i3ry/EVp0deyQ5wnnOD8mPeWAbHLjfi+GF6GHKljVMQzQe
RcXqQ28/OaPz0In/4U4kw3owqUAq6WX7Mokdbl0PEIMWMzMtokfaW8e0XYHANWWK3uB2y6NTFj2e
Kf4f7CKOzovUnl5JwonSDopTZMtyjB790vTdH3uNpLi1aJAt3AST+pT2dHEqutecifqz8zrulhS5
TkQ5Hvs2/sJNa/ND/hs+M+DEBu1cqLkJXI5eTEb2uNL2kcaqgOWeO9qQ9nS6kbzYKnpNVvLOZcPX
i58kBdG38XxeJUq2bsx+XgcSdEQ3RARDrakpqdkp/BRNT1ZtJYRhcYi8+LH4i7cvSPT5BIYBAAfi
GTgzuUEnDsYT92qtuTMXWYjoBXttRa5dgVpSEGz96yRNLo2DdRVhcNgrtnQc5bWM4ZjPQ3n3l/UP
zI7hnsnth52u06n9MG+W1WkUBcm/sDpyUwFyZ1+jnWqR+GkSGfYAcXX02zsOEmLl1TFziv4DkzSA
Airqb7E0RYZSFcSCkEH6OLZAqugRP57rPXIZU+th7Xh9sZO9eyzlBsRUw+6Vl6JPUdobmoeHc05C
nhHe6j5bTh7gPTby36zuOnDO9jNm5xlxlaBS/HzP8Wvbgk+L/8u358s8PK3Lma174L9mjwZLQTgl
Z+KHxwFNwEOYtfgFl8SwGveymJM7g97qYU0DPblasZxGvKuWBQdZiOABDMVxstMq/SeotENamDVa
j4WLtY4J1Mbr7NbhJJQ/h6ntOYj/y1cxxoUNKKlREDgGR8Cqpzutc/Wp1lCzhPdZqyPFWOnbD/HZ
hLpGx5VsLjupp/LHz2jbimZ0rhS2l2RjVAqd0mY5tmH0o1Qs63ddwyoSmXB3UDS2XymkcdxSx+P/
r5tQYIv7qLqVc+vnoyuKutDa4s0PMwZkT2vaxk17ymezEgzLHo1WJy0rPQnE5krkUOTlgjeYRZpO
w9QIG6MoYlRs8z9i8+d6T9ri542u6hQR827Vm/UoTPRt9kmfs+QhZ5Czxcd4oy6vxvW7HtFmiIfA
15yWItOqJ0aVJz3YXa4EYcRSPShBavvSGGe4FfOarup30Egg8KfLIWOHQvu22iqsjj///495O689
U0frbQ0laNHBNSGmNzSBQgzKZkdXY1j3vCpN/g4MuRR/+v8CD9oDy0PmYI9ROeqwhBvgxh+sVuhQ
e+boo/1vu3B1L0G7mop2ueNdVms+wIU/ppZF/KdDjhNjFw76hhCDbSp+tXdqjlmwo28JzH9htdQw
SqGDC0CKzyoO7goqTiN8nC1/QsYa+eoH8qSUTc5lHAl+V8GhxH/7b+c+ReItRtXqNvp/Yrad9z/4
F5+p0Zn34tyfrtmxhlrUVCkrDa89Vkm/w/g9wJ0MrR4Ic6hPgRoAYxaE2F0VTpaBTUOHt7yG3cOE
0MNBsDk+Pd0HopvHTVdqX1OUGAEaFlQKbd7GqfwhQiHVOwVEGdIt65Uc3LP1Oj0abpC0ORkQQxnv
JINmpVBtQsGRk2PeOSf5DnR2GtXZPYeVAo3ZSwM+xDoKEJsPwOftlMEG382AhlKYTsPu3xEKO7j5
N+1iN/cZzEcfPk+7guc9b1PZAZf0t1+oDerDpkJJeCokFb5qXu4KfywtTQ9RZIBJVK3i+o5B7vf/
YIBeg+2of3iVxBQHGXz9xM5LoO68+OoamGU9v0/eQZgQOr13U/3ymiuEAvMy2DC7U/7hfiRxIfR4
ETdVWyst6XyU22biU1iHfV6v/06WBj4vJXPvD6681Mst9rIx02rsHoutQURh8+IZ+pNEytkR+6IB
rLKc0rFuD75ezofFxnwsrYY5mSmKBYOl24FC1GQm1sFIaGDYFWiZ+lWNNHhJ8A/P52fsITxJ4bx1
gCmKnLuRgtscWnBlz5D8Gv4n+cd4f875sjvQwsjISTTlp6Ncp33acQohc1OBLvSbdtXUhbeqIuTn
BfDtmL9kwQ/CKky1EAh4Xvcm4Vel4GbUdyv/9M8rbDRm2a3igPXOjs9Doi0zFitXp0cnbKG6WIzl
Rtv9yrN1O4uw2yoDEVilq2HvIx8MwzpDfG7joreeEG4ajgarNXMyhEPA4FiNEJhlPukuA7ufFXf+
Fu7vzDF+rO9JVu+AdWtYkqH6MeiJbLc28dbbLOpVJs3CBi0uHA6t3EINW1V/esde+6oWC1a68wqt
nRaGIeJhOI884wghngVmyH30/W15IzCQSszAWb2UbhlK3XClTZQt27E73seWpCdBq9NhRP2Gpx5h
SC5xk9nDtKgYV/DM9gkQNr87B86D8G/afCUmdnB6G5nYPxLQ0zYSb1a0W0EOANGm4AYhi6ggdBIq
hLF7Uz36Nrugb24/hzlVGoqLJ571Kvfjqzk7L9VJRkeukNI09QR/yG3754qd80iiDMw2NIWNv9EC
sgSqin0hzvtbiYWg2QJ5kuyeXayoGyd8CE8PPjDAQceaAG1BQz3GhVr8C2WkncKrxp5Urk8gq4fU
ML3Th6mMAhTYakk43KMwbogTAieEKW8h0mhlM7hazfqR7/3enihQ7H92Df8Y368QJwjIJg76NJnp
aA17xAAIT5w1AXQpIYsAetBdKGCwK49hadcw+12GLyY1RIxkL9xXw8XJUsZy5WRwwY82DIY8UUYG
A2AWNnNauZjD9f25RrJKajiEqot72G9lG04+ntUA10Qo1/vpQF9zYVz2DjshdROyLsa+IBMLycBe
X5Om+y/VuMqjQk3RgL51UpE/tjrnZFO6sAYNPKVX5BK2XY1M7H4Mq1cawcn3en2OiemluqPmZAHv
4xtHk9+X+cf0IibgE65I9KA68JyhTbcBBaieAXmM730M6Kxx4fErytScsK4/vujxXYizO5kvwUY9
dagd+ZRIiF5fCXysbvHxIhmkf8VrNSZ+ihrhmH9/filnBDyCJu6m0lvlliCSf7BOeNmzP9Ap5iTJ
zSCgmn/0ygX/5xPmJyz+bfpnOQzj8459lUg3viz9zE+WBE9WDgF7b4iVvPG/zXo/S5AthQD+Gyv7
TOJUaH6om4vkD805bzKYbV2Anxm/DGRtfIOhCI+Dh4ZXlVeKw83FIX57CHJsr+PIS/EipEaoy57o
yEf5ydQH8gunsqCXPKluyPDRyzAuqLJnpubLw7sVnUDsx3i9wwHc9dOgYR5I3a563OATTNo37FCu
lMcJiEv1VwhEPS4Jlhd7YgNysIRhAQx1pOO5GdGOD0YPthjMBG3VkkulNjLbc4QU7iJTjffsPJuF
L/ie19vumHcItIRHu1jSs5O8z6ZS4/XcAbGQ2I3oQvCzlt6qlQKof2yrCJ8d9JocYRYQQyya+89J
OcRQTJWU9ynYClezVDRA2oKbWaU++4kJopnwAZdtiilEggzIAl+iyoXvmgmHTI4Oa6ycMIUruVNL
IVQ6HowHbK1yzBdRZ7O/56Y/JMt2EOku1SWKOMomUZlkZZRiS/PmBv5IvxRuejjCF8n+5BKrM3as
l/KeM7xYXvHOoEi2Ex2m3/yxsZ+NKuNaWj5Ff6jb0d4PW5KLmYFkvbyFuqYIl7aq8t16xfu9wK3o
bxvzmuWO0oIDwuCqvANvpM4x6x0qt6cd9K4QMD8FX2dHEirTwM2eLLwQwBNVIhy5efrNsYz/OEdb
hVhLBwwWtuaoVJgQg4pKPSXmB1+rjWp4f5FX2697TUYFfzI090Qp0EHURrZ+Fz8fJCbP7DNTa0Si
dsmEHoTs0iAaUW1fHUWC+Qq3ew2XnfX33Qme18b5WPiJz2ZfM6/uY6JPq61rSGwDZqm1BudB1kuB
aB4D+VnRmvbZWskT6cYZAyUKQw+Vx1j8LR17lzACTAW71Rcsj3Vw/Cx3jW3KIOyBhFEK5pbfYDY6
yWNXzwbEOztrFCoCY+6MmpK/7iwfGwzkx4MQ/uhTyqy36hpbPSp1ndgTc9h1ozBdMtW046lqPjvX
B5ig6bT9TV9GEywHer7TXLYObJ/9J3KpSOud31EuJSCdRLS9XB09dN/fRRDFmf+dadV9zsbeLGGd
xKFUW7pRq9n+OVs2NItijewklV1mrgPoH011q4sR8SHypSL8OrrJ4OFcdVfvQ/w6sxxHD6nSF3+I
qWoPNRFPfhkI6wbVxyiJIHgjUxINNMLK/foB1cBTsOP7IpXgUXkJh+Eq4o6y5ynAPX7AFD/PpIfu
DuTWtQg9uwcakll7ubYq1832i8AMXGXvNJkaM7DIQT1zDn2tUEyL6vQ3mQ/3x0Znv4Fno7yGAolG
XosxJ0wZDqq4tFcRNVFhXQB9imtska9u7ByRfmgKQ6PxldRZ6XlMcWGY7DW3hjI86u6scq4v/m8k
Eq+92RvOjQOd+zzEgdRSKPIwFSL//euHWIwEWWl4tvQdZSMd/VQLXFgGPJUeAuEiI5i/S6iXvnXe
Cgru4NHYNZDJxt57b2Hyqbz5WG+m7+55Wxj8zFHFAxyt3QKVhG1JlovAclsIZb/1ryiewjTRWepf
wMjWAklEbH8aFsnLzsHlNCV1uhG0Xg5gIKMEDBQeEmw4WclRUcH8965ebMuw6y8wRkR1N3E8sTPq
wRSxppF/Qv+LFSLD5xk6D/Spn406wbKLv7EvBDeNeOfxc3gZcr95xlHTAXa+8s+OcFRmSqu1Dei2
rKiA6k8T3JKzVW8U5fTal0emyTGWtYRiQLb4HFrqpNXdNggt7FnsKXupFf3oaWBsP1D6hElz7J7i
d/2C8pcGZpmkAfY/mpRq3xzZ1Hsm+HLLTciLCjr2aT0C3aE5uzAQCaJRPWatLCt9s3dwS1ZDO7Sc
KBuHvxM6ZFVpEEqMYaM6GZo8XNr9daL4iAwqtnk579zkyXhw/puJ380hGcJyN2I94BG8lvFnavNb
3mH+4gOYUU1T2v54xFsN9SpJeaPry044n2nkv4bhGNgKrKV35LfGcLXrnJT9urZNOITQlAzhK6Yg
qjA3IezeszCMs2DytfxqwPgJQZ407pMnzBGr+0gBKKHoWrCDfq0N0zC0XsoHsmXR5cQ4Mo7e8kf8
zHgCnJJiR4s57pT3MKUu5lskyP/jw8PEN1V+uUINNEWQriaSpRiml1l4toZ/0rrIJH5+nyFJWn2Q
NJAe3UuqJ1O86NR8hhq0OvhtynOU4/Y8TmlmfWROVQM6xicryFTAJRP35qMcZ3+q8GzBYB5UzWuV
Mk/fOxMwpd+xKZJ9CEjnfKqH1SXTVzUNrvHyhMajjLyFKCqWsEitoVspn57Hz7asUdaZpiXzmj7Q
pvS0cGah6gnTmLQTXhOeomjfjmlXFzjs83kwdMMMbfzayI+pTjOWScip8RGg+ha5LSUcWogcDvLj
PylmAh/UA3wzEmD8JwPD2BfLps55WQTBDoZy/je/lyQYwLdSOQFBMHzNYz/z9Yu6NL+Dv35VnTDT
J+HiMJZq4RY64aE4lfXrOqbeuQJyw8202T9Iu6IUDpDiwXDH71R06aQgXvCGAPNCzUvrkCFSgn4l
ZOCgHSYx21fGs5Udp7kr1jOeBwCRkRfRn/n5khx+VtODGn6xIm5FtVDvG1AJ5BxDuuPks7vY+hCh
TgNhKdmEvbDq5onF0+b+AxOho5Li4oHUUXrQX6nQF6KjyUEVuPcJy5XwX22QNuNHLYh74Tiov6i5
ifABplzeGPj7G+SWctrV1qw8m5L9EQMBrhBCzmlkJRP4xXHL6iAJBQTCepj5FbQ4pC9pcjzbsY+R
s1SBz4Q0sGl4cxcN7nS2o3LnINSd6y7Gs/3ygNd2kjYsJhnVhBaiGIUeonrEgOIjtg3U9laoDqLG
Vqe9FqY1gy+dmUQSAUUJsLRgUhhe8piB6SNW4B7aWVhS3cmpNdsLLCLUvq1yo1kGM/TodguqpiTy
I99guTg+X7iqGK8RTkT3/3IkCWMf+vj89gl32ut2OlslUvcAbzUtlOc8VPpILYruMvl2CANHlZdn
aEF5or3ExdwJLNslzbdFbafdO1ArTwHXb5UQ72f93I+0/TfRp1obZeU+qFeJlfbdQ2ah5zdpCbKe
eXubKxgyDu6f3N+skYWti2Tzl35CEI6bPRIiXoFBSu+j2vn0RVps2WxaC+RudpSmoFU32PVmocwK
znCffQxibZisQds5vZ8NCrRFWUqsnPBynD6VWFoGf7Qq72AINovfLlMPYdr9YGtdzuiXGHvXHNZg
p/cD9xABGKC8T4Aqfl978l4nFB1C1i7lg6UTqOkh22rKxN4YT2oiXfZS9YvE4dk82C1cGZ4PHELA
vYB32C9KXdqMYbPqEmtiJDd8tvQj6uI11MWcWBFSBn2vbOOd81JpBhPSoeV67/tPwDgirq6Po37F
HNrYWciDAv/163Sa0vPtWI5oN3peK9EQZGDqBnEnZK4r44ViiVFATyIJQvS994SWhGnnFfZCBeL0
tT6s0pYdp2+QTalGHY/U2mq7Tu0UzVi+wHTAopVfj9Au8DxiF9lBrJyqwkAinVQIBsWjWBop2Z5/
IUPLAXK7ER7n91ye6now6k18e/xf7xtDcZEQ47/3SA6DEL97uRdCUJtYhaQuReaXtihdNETKA6jY
ehb5oT1PAZcPzmMMXXpow27t7cB7oLwQgA9SqY6CA/ZyaV5ZG458ByQ1TomcddXO5Iv0FBaxokyB
+PWciNEFbTjShO47wjI/RIdfriY3AlvB4d2JyS3BPPrSVz08bhtVaGsQMH3hOynZHnJKz/HRUNVT
9RTDTTnBTngP6cPVuwGEuc1U8ejXPK4eR6ZlhdM9iF40dB0eGFefDvNsIJD9pKVDBeoh7YzsAVQO
bwtldd7Elq4ROPLZDJYRCFSSIdq/2tv1s024Uf1Xdb8HNWFrL/fPC8MseI9Ai/N2Lt8IAUcXEVf5
YJ7hn5zyZQDRsfB/lWzbc8dd4TB4EyycHwlUQOthBk2ig5A7Iu7r5Iy39WW/N2dITOE7Q5esq+s3
uywtjb49IPMrP8x9NhhLEIdpnLTeizDRQoAsVGMIBJm1Hm/HiMs7LfkQ1KTnvImr1+2mF05hfSAu
yK9I79BDsTPlFekC/h/YXEpSYAhSOpYAwyFOqMM1oUPZKndeTqK8eIhN8UW31vMUA0b+YdL3hWRy
VkQ+7ouruKoltIPa18fi5HVcKiZQUii9jv1bixG0ZbklfaM+Qjqbnb6K53byvM26v0ajuK/8Nu7m
YDb32LSgcH/gDUEZ/zGQjtX7S/vd3GrXdjndlqCMOLrDsqcxNf+2kG+MsUpUqeoWmlJF7bMHxWtH
PRiWmpSmabwfP6+itu5eK0+NcfwgOwwywSCCYJUz3+uADr+9QN60emNxXlgDZDiegVPHSB/5WWc3
sDnNeY09UhnW1Pa0UdMN0FACQJ7C7XO1SP1jBBHql39AiMreJJlF6VluWZgUyi952ix6ABtHYJKb
2uzz0ItMOt1V3ux0PVi38iW3sSeIbUgwzssGDJjIXrX7fiMnoiMlPFibM7K4EU5PdMzOfRyfm3ex
KzU6r96GrSMi61b/XgkkQyxERlouw3axwvcGsDRIkLV5V6DEK6Y/ipEM7A257Mxw1crgFePoLWR+
cz0aYn/z8B2bLYgYbmXutBx8PwUTS9LiqliAjw6f+fFbugEbgrKTQX4Bf+xiPVZlFIIO9EB2A8iL
YbbNluAbw3alHdiAM/Hh7i5czZDdP4U5L5YC9W1phDqne9pePxhUZeoLYDfY6V6AcLtBZCdFXzgC
0cuUvQ73r/Uf1WXmKVpoOcBP+jbpkQPpkk+ELwVOSJC0V4GsxVXfaqurLRmXrXNFRfrO9fg2BM1S
wkBRqWD/RwiBjV1ChGni75DILWeZMofUHW2Alh1QlBrU2KIka+sZtty5ux/x3x6qKWL7Jhv8zY1G
W0q3Wm0w407i569JT+oZUMWLzjLCHCkZaeywNKpLus1BoiTvcFEMUV/3+AEpbdEJmoGi7MeLGP1m
qsZ+IY5pMQKHapg2G4xFkIV/4DduGD8fu7UG50viVCYGOqqKhTpEi3bSpDhDwVQUlq3OWZauJVzL
tcjPMg1W8KP7hvXSOJ+MTE9J3cUARGjz5WSBhBMIYd/qjZfrYMQJUihv6rYopAqjvBuYgQv0oaoU
LhslIAkMmde6Wp839hqoNppMlWb9JGHClC3qqCGMLw+LD9jNixiXuIeVSoLdI++0acADQ6XwUftQ
gxKsEUjTs8A769Bu7b+gZF+j2HcH1KI9rCSYaQKzPHT4hKVpxzFDdMMHjg/pHt0dVrfSMHOIb1j1
0SW7+ipKXPG+2yWgTuKNc3sGqJ+1SKoctQTdYw+dRbHkZmKv4IrboS2ZByBU5rjJ/X1U1+xojMvU
80SNzhNWtmmf+J9Z3MmUZHqwF1E+hjGyrTrJEOib5gtJ9BCVeRY6a6dme3Tr4JmEb+mxOANadIfA
aw/yLbQaLPYNs0k3dpibLUSJP+EkMB7J0nO2zwzHE1MBiT53+r9n6OtlspKl+k6+nuupDjpux/nW
WEjc4Wpelf/Uesdd6OoLNYi6bU8bVHCQA4aFSqeE0GFwcFJPRbPlEwqA9JgDtmfZ7eorn2JFm5p7
1ZqsIV7QXTRgAXOrPA8LwDHTv7ZjSDUamytWw7sHia0DZhMFGK1h74T6ci8PV6IMTZujEhC8JUTU
VwuOEj4rU0GMvRxv24q8VdDOMvOMwdATwYgd+9bbjHQpH4dBMM5h4jax7Kjuh593R9c4j7JE8ZJb
TVkVuAZLVGk91zRFZrq9IjlBlxPeH9LSeAy78KsdyaraC27m6k7EkjIBnJXQBSspTvUZe/ClnvX3
jdF6N5TXAgCkGu2cbQ5arxIXKVoZZXt2cl40Hx5832MQ68dyt6q0rweHgZmwmzqaMKzqS9k3yTZ9
rTLy6xtUjSFDzJpXagdrpCYv12tH0hC8RVhWWlElkAoe7BmnpeyEJWlGhjxyEJAnBfwNyEuS3zbw
U2QApBE8oCQ8WIaCb7aT5C4ktgsOawxjyUgmEi68BRYQwBvvpr8A47ToOa9/ZLA72ZE52tto5CUk
R8XdwZvqnMVlj3p0kTujPFfrcRcJ/VkLjxcRy+B7gt6Pq4su5BKl+GfzYkalJiT96bF4eXEESsuE
e5BJE/YA+QHKuzt9R7V/umsLsMXFnzYofgdXmPKeIx/IWsXQsph0d7Ok38oSZCRLen/WqGn5q6zg
DqXk/GnZhXHKq/jbogwbAYBY8hN5pIbPfzr8nOsqmsyQ02Ab4FeDwTpFCbVhPnbmbWkeYYX7yHKv
ncTdfXwb6SXcj1NTsVhVxI2Rzub65L15yHGF5EW0lgmBZMa6c0GhYHm62Yj/30gkuaEHHXeJJNFh
AKZv7QHUcazqiTfoXNXiUPOP+EFF0vqciV7MPsP2Pg1mjJXDlXtDW8GXQJAErWvFFWvlsQb0o8ex
yYCyBb/fl4N/tux6vvrEMTliTVld7/dMhcnLz015d/sSpEMpNX+Xu0to8f3qY6ps0TeVwR+Wa4a3
/aDMvibo88mnZ/F7wIx5DGulg6kMDnFEMTVHuj1lE064zRkfhdgEMHUVdlVGZFZy1Z0arTkdUGUW
5M5OPWdWYXvF5mK4pvv2oKQY3i1t6Yc7J9Mk3YaDl5F1itUErMOE9udTiL5sGFx2fOBulDeeFhdt
JAVDHlAv3jaB+A+HyHIeW7/1uw4B1aZh2UUSdpTGk9rbqZB2z6F1Dieyz5FHpGQnM4o0iBMXiH2i
TuyRiAfM0yeRepFlKtWbqI8wU1ztAJQi4eDwdz1A+maccRj/77mjBOFD+GNAIoDA0BSXVJor/7nJ
MSJKXLCVd5MLmFuiEJj0rcQKwmv0XDEaYt8cOwrpTkBshmECEipHvah6xgENrVIPpy7zKo4A7LPr
JtWPABZko01SJIpokDxVEThHdnlXu5czKiOngNYs5XWUFI5Fw/DCvEd3r6+bGSROavIYmE+3WWvG
gwIcg32Ee7uH2piYlQak1GUDLJ2RO//BgQYFYBXP28pYItnyL8OIwOO3xiltEl45tlmMofFTVkQX
FI9aIrsBzvdJIxtTacfnLLVd1ounADXoedeg1RJeoGkXW4+pFgtwSzq78goQV4ceis1115qxOe2X
aapIMoQAruMz9KON8wjoZQCuh/JoqxEYS777IBPOPegyZp2IsqXuUZFAGGjDdIzV5lW+REerr0LT
cImmsbkgMWOqLFLWTym20xLT2JS5A8NenSD8sgzMoAEQ8wOTsbj2TCcswyUS7SqQYg2hkmjv+IWU
VKNWoI4S5lt3Eh1kXJlde2ndcmYcChmCLeq/gcxxfYWZKdQlioASiuiGBkB9Oi/h2onG0E853iTg
r+h/SN8vC965ICT6t6iEuRXWc4czyT/6pp2h6j/EEL0Ndi7ln2Z/EAv3UGiR7oe9tzFvqT0k+ZE0
TheIVLRyNSI7E3F3Cg8J5+uNWk42usXU4ZLHgnhxUVyvVtAmCII9ijjQr/wCdc7XLU1DJrdoI4pL
YE2IadCWUibwFnOsgxqZHNta3J1FWi6mps/DTxfqG1VeRuuCqCodrWTMdyO3RMV07kvdTQ1j2jUB
94JX2SUrpV37h8/jYLfumJUClvzdE9T4d4dAO70PvSxdMDiWMC5JW0q6XYZEXyElCmPjQiaIFWOB
LbOe6JGaiq9KZCIrH/idtxC6Wn0hL/qlZW/0p2IyL0Q2hhuyfHUB22/zqcYsBD1p9XVMDNr3nwe5
/XVsPJBiZftrbbhiX0pdyQQYG41lXhNRdfqxAjUGIy+fNki+yRdJeg0Ve/Pliw7k1iF/cZdsR/gN
UU+spJov0aXjINMHoBVtSNLFerugaqay1/BvVtbS8Nv3SfNKtHJjW6dSRT9YBI4EkpBGB3DDwrUZ
7eXCECyTBVvHGRql9Kw1B9TaL8KR5GHN10GtZvABgHXkspztiMtEdRxYK2OFDYnX+nnJn5b8maTi
6MnnlIpm9/vL8PanDY//0uAqrZjcgOct8BBJxIu1GAjQwNxOuUSMnSCCIaBWypNTWOziXWDc9lMi
ziyYiRhVrQAQEBOR1/viDBT8Vk9wzpa8FhC4+hHhgryztP9KhrYrxbl9nOZAfH60XNarOQJh77ad
VFWIVDgkkXDRJfUxy/3Y64ObICFzOmW/EFIz1HNyY2+omm/xSEuLCyYbvSn9+FbEypyztu2aW8+T
rezCmkTY2aUpgnHimiyzGbNT9ltL4UabDv5VEvSKqOT//LEZHWsnnLfmil3SM8FORlrbUgFdsNtA
/v3PxPY/YrxPFKT9Klpi2bMva+o9q9ZcMkBLCaiSBVuUE+L1MwwGZlYMxtgoB8cSZNXba63NEAOK
D3l/TWv+nanuqjzekEtbXt7nlCfhQ7R9AG39b9tcTHTDSvRklx+NSnqDiBb3MPhuERtvtSRfTl3S
/MoHXkf8x+ZsPXVTB+Y2/anZuLV1ELAgAc2AkZ8iw3P0kptIJihngRXXyNAcd1o6AxAs+taILIIX
acSmhqKT5dVeGET5609/iXeABYyBx8ccoY/DT+kyy5CDy4ObF6igaEPte9qGCvzUNYIQcdoCanp+
ghafnKkCbkoqwJPeISFZ3XXeIHG+056s3ZcuDe+72MFNCholoeGdJL2PSzDMtDf3ULUUt+r6q1OG
6mRIZVgSeY3MykPCdkb3GB3oRQN5KFQYt88dP1UlKzXvZgY/uFfbCJ4bX8ouyDZUL3rL+Rn60j8B
eDBb/99QrmrYwGG64J+pUMnWUh2cPtt11Uxd5fpjjLFTdtayu0/E+Z442Jdao8gbE+78VM7PHQkK
ag3jxiaGaUqEgLna4gHH4Iy96XYztXUjDHZ4mvE3NO/UTRBBi7AZSczEHaTea2B4DkzwMtYpVWg0
1TkeEjawub9gcMlhZDtqhIy0UJRsxSVgXkDJR1oZJqD/JgpNHZV4/PnmsRSOCTDLqZyhSfeFt9bK
pODBKFONk8WKqwfJav7Kl6fGt1tpktNxwbxHj/fWeADrjdSniA/RMuaAOHdog0nJOUI8nYj9h7O1
gNLMSpovpskw95x2KRQ3Rs0hMVlaG2+09n69rWjOBDwGivalM7tSlfJGmdp1ZZY6gcy0dixwF/P6
hR4nEXvNQr+4nNDZbF3yECIJcwE4oKWS/vY7WAl017rco5VEl28r3f3vNRlTriqumTL0v7rhi5y4
w+bDeY6ugUyiXncKfpUzOWQgzJnyVfSPF+VIqgejE3HnU3jsbOzshDAGWVhQOhy2L8pdnDjc5jpI
X0f9OH6KpfOBJcDajsSIL/YOtwr7L4zx/BHKoqf7vinOfXF+JhppfcCMvkIHHaVh/tYvsl3fgzaU
1XUVnmq8OTMJ3TN4lY//PhVOZ1b/HY+XrH3mh4HD66EphR+Uo8yQgjN6FKJ882TH6Dglw9E89V0X
RIQakw03H4oBSAWyo8C37BtKZIIymj7q9Gst7Vyl1GMmmIvY1Ocq/u3DrHMTYS6O5CjsuHj1wMgj
sSpYGIWSttJFpybz0GIkzRl16Zln5Ijs3/rNfRqTL97sdxXct4Kaj1npESK8ajJfafQGE/DaIrpR
TaTjw5mUEmdfs11ppgow/auSagb0cTWW+VsRDarXd1nyTg2t9oGUxOvIoET8oLvfpZKP5h/r3deK
s7TPa5hd11nGrU0p1RYWKEOb0AzaHE6DxUhxyKlEulLNIhGsPgpKk7OF3Vv1nHQEXAk7L3+Cm/Ob
eXZpDVUWHm82NMBTPSHU7/mTbaWNaLRtWNYl6yE1KdEwJPe74RUMaxPQVlbtao/Ly7/Cn5nUPC/P
HqfJQgqtpnNkZHNFgSAmOoxeN8TFyFhTljWg9Cl438fdmEgk02kqF0VbKYuQvEjI5uXP6zgB4KJs
vnftZU6okRnISANvvDW98RTG+34pUi6yiyzXTFKRSW/lN0paWU6Vemz6igmKT4ZeWfZnspQlnn5w
MOfLhGzQrCEiHa1trP91s/zLVipXEBZlkZRZqrqG3trLx+XTnq1rqkbWDj9Zcum33t1L+w1l+L6C
DEYvjr5iNNgh8QcXeyz1nRb2J9diWUEwdZv0thgqb0N9QA+uq4q+KJdMohdGiNL7gBIyKmIUozmH
I5KdSemNHwJORgQOnZGZnpO9NKim545ubJANZ1jgQZzqimIs1SNA+5yBIUUT3vgFBQjOPtmQ8n4n
P73ILoMjoqeRuBaRLZ1vw/fiDzSkTSfSQX5UtM2kBAYgEEFk/3gtPHHGOgPMUOINzVJsXztFDwyR
Q2uoJ81Wjb0Rdqq64NlmaH5k3/PUnHFAANxfb48gTZNN5JfFxtWUjCINuh8vTtGbS25vgIAkqfdz
dHYxz/wA8f7jCk4t2J3k8zDR6bTwfCKo8FGbmONvmOgYmkjbt6EUAWXRQsgSX6p92XXg0z2zf9ga
8BUYmGL9CE5C9VQvWmRmzZ4IYMGsiEmx9gfU8EDuiSvJSRu6g7+csMGM97mVyqZGP9RLZ7Hi5afL
/NRwR7NLKxVscJ1HFBaZB2mI7qR9/obS/2YCUiNN6Ygf/yf0EJ/Hr8kMOKWI3ZD+EcTo18Idqqnc
vOQc6tg3+ysNH+DJJGsWaqcohj5Y4TGltXtoVPisqExaqCQH1WnbuFuFt1uYFuLvM6teNGrz6v1P
As3w9K5b8SkC8qzxEdxeRlKTllMS99V1bmkF72lU4zhUv1v/H4+gFsPQAVM1yF0jfx4eZq7+DWGa
kYLLVR0+K7ANAUqDbfyjEY1WRW/vGOuPON+BUbcXyct8y/89HiTU4Ft6CaynjVa+1g0qOfPoK6gs
u3TbXW3Jh5Hpe2oRb+s9l9V0TOXDIyVy1jPJdiKszM4NyXGwFYCJI5TaDdXeJLcW73hWxiKLUE3K
iSMSeoKCJdohlSLaBaZo5mclaK8JCqiiBH9WcOeVAJTCpSHieEdz3Pz4BEc0CfGGDCoDeFq2KfXQ
psX0ESiyNsP7CRA5XX0S9tTUrJHK+xh+jG806wWoVWJ7jpq8++D31hGD7AX4Q83/ZabV/vF/z7Lv
4bSHqqJqwyj/ln9YARWLGKGgC/VOpx3eeQjs8+1aF946285fYO9LNrRCqPhXsrA0vRpSMlEJv9tF
wPwcpIB7mBZZRqgmRMyj8h3DrKfAEBqGP3LnNXpw0vfNjaSQ7cbvzZpchkibXXXhjpIkJM8Dv6kI
ah7tzTUuVUwbNbSdm2/eBLoJ421G1K6zzo2n6WUGxnCRPvMbA675fhplDfBa7nNU09Yo9kuUc/Jp
zE6UOfdSg8n3OCelJ5K2lv/C6LGS7rpDlv76M4UYixAD4zRnMR9vFr+MW/j69DNh3A5s+xnxrQSB
iQI7fqn/ka+myfJGnEJpqB4sBDzk1aX00e1U2OI+2Np0HTi4txxikL92DRZZtetB2xJFIJDCRXH4
ZwAG93WVT+x5m6nTcmM6fQSnfwqHcu823UUozlSKamSfMAbIWCIVlC7T5IsQxr7BOFB81LswBC03
eu4gehBWVcolwMnGMy+CsF7fgEZvu97lHKumSJ88VGZYDFc2xrUaZtqS6Qc53v5/hracKXWCtyUr
DwHrvdp8WyDTIPIRTep2o0CmjX9UBc9ESzv1/WPAYxBnwm2wbHE8HgQztnye6EGMe0e03NIi1Hqz
gFK1fe6X0w/H8D5czV1C3JoojG7UV75TKLP93mzwsh8bBXPZO+BF0lif/Hh7ofIzvzp6qRhgckyS
UeuFzbT4Gk+cx/1w3RZ69SHyKm77y3jmliVUttXASWpSPPPLTDUT5TtzitjokL7Ramz7fKRTNFiP
zTEBMCzdTg+5goPcy0vufhnU31nmuHuqakb2PxfjEEVdAJ23u5tk3bl2N/4S8TUXqTuSuhgfHyZK
ifuiZf511M6n4fOvVTb0QZKx+pkdvkzfXHpeKNHaweyPm2tv0RrokXkRSl5H4GBRc4OTI9aXFxrT
V/huR41jzGrB9mWiPqY4bYtemqvcTbjXGxBPkbEwMvdGPhgJaEa2CXL3GRFSN3MJfWuZqGL3dDNG
/wQI3fhJxt2A06xd0aZNHpIbjZGTtmdCky0957Nu63qvEdQyW7aX2kzBTxpVmP2M8PU7iAv+Y6t2
nkNz3+hVCwXT+CiZzDpLCkfduzVM9NpqU3tF5Twm6lr8QP8jr+sGhLXwSl3vbvqN7ht4HuDd/MDE
gvkHc7I/6SicDs92fpRFwkS0Aqdjtqnz2oWUKOOyay2Hs6tFOGG7nmNthftxoeBGHbs5qePYVZQI
cZAb/e/4LYfnPmTTyyyyv4H1pHLjK/ws/JC2yMJms1ZGn5xfAVfwsKhNbH2PVoJ5NFooEubAFQOL
nYcshurjFNMAWBfVWMsaHKPeCXNvHBcpJmaDpOEuHz/ma8nXbrUU3H0+PUiXZoyKLIOvcOLqF0eA
bIBgsHuCNnahOC8NqWUk3y3hewCt/FEKSkX6HeQIk51Vj7EtMlLV2ViNNtswoBB9Lu55NtC9zaGL
9+vwGwzWPyAGW69IK9nvolEAQmjeQ1CP6i0nv6mdbk/IHZRYQfqolTesuJIf1FMpwrZFjKcUUIQD
lAZCXFh61KMV9xsSxLHXo075m8OJOvWzveKlyXfwvhSW51GOAOdVAvCM4/kHD711UxTIVcM9+M/h
kUtezmLvpGeNOE29uX8bkqJR+tqDzculC3RHEw8sje3nrNkV0Wg8Hnnkjii2zSQ2k83xcICaYWQo
Suc+cvM0eAaIywlNiXeb8oVvznc2/wwc9pv4BrvHGr1kR1KmmWHy+I3PGvpebtz8UHhbOJH4dUd+
p8aUudoKgxZPqASxf4yfoigwaSC/VAFRGe8/+yRnM+AuMRKa+K7KyXZ0l4szsPoDqQh6T00RxfO6
pMsphftk0hVWAomoxufZt/UtgQZb4CsVYM4E/4xr+RBimDVMa9NwHpHf05/hwQ+mo+5I3eWjkcta
KCIOQexQNzp03SGfCWcpAOdsfyFK+8NFxwrjuiq29c9TH7lwG7Eq7xWo4zb8itNiWqdq1CmVKfAV
hK7yssY+2lVJmRpCxfO/u8BAU0sLcjLvV63Yp+kIVvEBgjX+pnjCRQksgicDbZOSg3D4LyDqi+c2
olVn4FaX5WAun1Gj2YjBrfuG0DJHWSLQupzcfAI1DuMQM4r+7DLD44uj6B04pRdQUNWdLvfkQfPA
TUDUJHNLJB9Vhi7cPfV7peRPo73kI15BHtgyf8IMewYW7UjXKiHOARkP3EIYkgRRPjs9MGIXqFlR
Mhijv7PNm2yGJ4mwhjF9jIURowkMKJ5oD5XDxDFrJPpHWfX2xluRAo4qjN/h6KYwAjlJm6uazzFj
oY+nocV1qc3NMCWFGkHSEyrhHp2Jq7HvddeNrPsbZp5P9JwP+Dl3dCk9TLAAZH4CAhwl+/2DhMZp
E8riFydIvrzTFCrsKhOofHMkB/J3jXceyaKSKWVIffjW7wBCniXoMRrhCPlm1QOouC1IZ2chYrAZ
FtjJfJFxp+VAeODLiEpU4HcVEO3fTng565BgjuFjo7oOMuPCRLVANxyePshPCwn51guu6pJI3XvN
s9g4pC0ACWiCUDSooQxdp47dUsuAK53L9325SMh3m7SZtIHi3NThvzRRKhA/Yr+wmjuBBNA3Yx6V
bVSuRfHWLU1yC/iTZDP3tMSgYJTH4YF9qQXZGGTE+u0BJWP66I94qG3UpNNrd+erND5Yn5EjdfIF
oc/rEbtjEGBPLD/b8uNMylaPkELUKq4hr1jv5aWB7oVangCiJZE0yjC3EZv+x+X0B+JYMatSW+ZO
3WTbvy9JJ4NOt7XmqUu2erVcpuR623gWOXY+Brf2JSpeoycZz046g+ulkzLnznycd6fh53vdjTUP
Ad7UcAPLiBAwQrx6bjlop4l5jhE4hGcJdPuaTrmD+A6ksPICN8FEmTE1PoxH/ECghluGXO54HLjp
T4eFohhtjO1TMvxOJbkpCgCD9gjzCqjzEQ/LQVtdl+5PKFdCcRc2L0CR9Ov6EBY9lvIgH7YDlXF2
HJS2G8tCY4ugxI2/gvS1tFjyiPDNIbovrLm+8f/fvU+vSPDcw9MOwfSdauRgyQlmY77dtW/58vEB
UfbYAREC/yLRVdIhJYuRVAoq4zSadimYB3Gud1nse7GIAnuWHwCKnzP0aaSeTtvHptTrJ1wPyuaM
XYrumKxdEWFgh7uTx5wabmZ86P9XtkiBgnDMUkIXOJPDe/2d/VXFW1iD7ezflbYyD9qWfS9b/3Bi
jgc1oNjBopblxvNhh5HH8fyeHyD0V988yiwqqREF0vdr1l1nygW8+9Krkei3epCMUX+k7q+KE560
ucVwC2LCAx8PFGW51aODDby0PY+SClo+D4kvSBNqDT/yLHZTqEBMcP2W52JDmu6H86mhfcTCr9vo
FR4LjH/O3E13Q0EbpvcvFcaxgwV7Di/KoGaItHYpTLZWopN4GBtFegh/HCd0x9G5m/KWTav7wfXo
flns2O5KjaLNWrAc/Ogu2aRUJPtv502O6UAtom++6hEGVycWKQXyrORiFYbiPCrBzgofV+5g9zTT
cprK4CLAq3RbvpiGxxzzMGcOXphgYSs4ERY0Lxyphyw9F4UV1v6ZeVA+QSsxvy2mYifYcgxbe3q2
Qd1IH17MDpdBoDBRW6tNR7wWIB9zWvV/EweKR/YsX8YEadmWrUPHzLaSenrFLCBUBEAWiJX/XgXd
UljkJPj5+H52AYTCvKfjfgFrvftFjFu0goahK6TCQi+/40AmMTKhWgOhcZsbf51iw/DUTam4vDz6
AYSrWtuEQgEq9BB6uFZjGxu35OWLbyNyZRQeVz34HvPi+Mo/NfK3+GPvYoKsU98A8BUuNnZ9Cnhe
kCdNd37nIpRXlsC0qebyWQXW5eTdrlNNtTdB+vJP9L8u/L/hgLho8U4L6GukaAihWEBDgeEyGF2k
j/jzodOakpdIYbqwOxIjsZiCndoR3KiR+s4ERAu4JCFFAFLy5l1milsKFGaIO6k2wvqqyPP87tSl
8sRI8hwPShp2JJda68RHN1qrTEa2uwti1I5Vqmi7/NznLbasjdeq4u4P0zQ/8gK+p1+5S9Kdk146
Rbt2MU7/vD9GjR9dKJePXa7mIuTqG3F+wwPf7WgGD8pLOp6WoWbGmYBHxpvLRHvmIYr3d3VOWR9T
aqIJ3C6CWM1kcvuhA8/wQIHFlxE56PHa/Gj9nObg6Ky9MaUaljmWqnQFQJizi/w5sI4uMdSFRIHN
V1VxMHkvQqfHs4lU1++wMW8ss5dctSS/+9NoyBKMp7iy1o4QC5ZhgJQH0nhXC2zm9wDYvlE+WH/t
gBEpLzNJx9t4XUfSbJi0bKd/wxHLinH3pgP92StYrfjvbwHcpxfrp9ATa0cR7uIvTy9aAs+0ix5U
lIguzHSsAl17ASFQ/pOJ7YIvK9dDJlmfhTLk/V/TerejOmktlmbN2A9EkKahn4KqGOzjXdDiggM6
PakRFqrAFgMbDrB1em01QOYqLj8lKtbQdEkCru363BXwcbFPDhkqPzYRpVCMsE2xy6getAttpjRv
/DgXYoYQUanzrkNeW0DTjJrW5EpgjRNdCqZaL08mSekddV8lN+sBlgfH9JQdUj22DMxIQxC8zw5i
+cU2mknGFmJ9eGHMjF5ae/tAul6g4qIHIO6/eq8CTm1SXPGNqLvOq4Uc6kEW7e4m1YKqkXL3RkJo
VuztqQ1bQKQrlIqqYBuKkJ3IpU7rILZ23TXIv1tj09wmj73qVhRdEbjj4RKbA/JKbG8jqLMS990h
585Sg/2fISWio3m0qzOPzvhEmWdJfQoMpkChE+xGsOdyryNjI4ESqpkB/HkWMzB46cm41/VmyvWx
WvRsEC6szohh9ag7gbIoVB1KEj6eKQ9rEcJFdG2k4nAbf0Nl1jHXmM55UtbQWAhOq13eoSwrbd2t
TWDXH6sd/u2anekPXBAFtoWdF61ZKRxCRtTbChr40+TYQtkYZeer+OH4+oRyndq/sj4gU7ke+MqK
aAiHbBMr0idDI6LxVweyQKgqlctw157eGw7GoiObH3zHVkEK3JzG5WMMbeui/+tn5bA4NReqlzhA
QJUvTEuLNsmdmHfbD5uhSr2EzyLPb50TLqVNJqv7YQw6Mpk/VVYRZlWerpxuAkEM9oEgsyCAJkBu
9mBGS0sTxDxFScXoEjBuGSootA/TjrYEmr5Eqz07evgWSEpWdUgPrrMqu1Z3U43QAceRFE3oqrfb
EVVEEugIA8Xc2enpNhvVO2WDiajL104DodbWZIod1X4caBsJ+4Hlngp2/J03e0D30noGi3J9GmgG
lkJ7fTpK+qNCTqLbQFpH70ja+0vNo7hDISgzb1DjFofmAsXJSop3q+BC8S1kS1Kh72LVZVs8o+HZ
AIHQjA76YJzJ6mWgU45vd8m4WTJvbogdU5q1+k9kZbZYnZ+/mJJJmCric6UfiNsivO9iEBV5H+5S
3Y29ZANo3kZm10aSKGnIledc5FgC1DFNbxEN8TERxKudilcjTobU4cgdb0qp2TjB4hUqApn7Zh/n
noaNbPpah/Usc+FhBX2GNckj/x+F6ucazOq8CXDWgJyFJQ41I9pBC+IuHlSiTofI9KG3dzTfluyY
5Pjy2/GhmKJ7JwyGDRos5HKcx8gehzzZ5aWNWzEXuA5rP/2kkGjnFMIXc/xpHGGHW7eofy1J/7WQ
+5mvHmUDNmQJkZYE2+xqkGjXwVcgn6ICpWcjoi3X0vYWLwmN6PrNPXJKnZA4wEiyeVthLqzHEZjr
dKdNBbePDmW7VgnebgYzImfP94IteeQ8LnbKe1p+W98pNRzvQZ+56LUMcK0sYhCrnb0Dm6QQ8h93
Y7+PwqfsdeVnyE8NXhqiDiYstRiyZshhlYi3cbTbxOVJ+px27a4xd6z2j+3mBkMU7BfBdhFy/8NJ
+0wEEN4cHAif+H+ENhh7Xl98WoS1uSbJjejT5dI6mBFn1Rb0Amm5shObutm7QkMIE81lY06pp35x
Obeuml1N5A/bZCYsjVXZaxjtVzdhGro8SeCrj/C+kMhj3bao0XRGnA4Jf/NkkDS3WapDejmPmlo7
FcF9uGuvBziTsz3BYfQE2lbP+teZWrYd3nbPwScEY8rB9VNf6dIibYQnZf5vAByvLd+s3eZQ1Y60
zvYEh1GDuetxVS2i9vI8v9+4n+XWODRwmjlJTy1k9AiA0MPhzt8Ya2w5t4Ar6lNegpZl2pwgVSS+
VfqM36wa9oXPGD1sJTqiVIO+6F6weR5TJpPr8ytYOXk7a95rEwHc1yFjCvMrO1iSYeuI2bH+QSWz
UdRm6ewF/2TBxndjD9d9rQ9bmFPymEFUIhH9jXNFGoy9wHlkN9M7v1W+mWF66wfCYk82dCDUah/t
78DM8/UNTlXp73J+k3psxaJUgLmQV4l6DERRzDJzzOiRS65DjQF+cv8ojCaOMq49FVDRJcFYEm3V
wLDnWlLiRrMjDl+A8okt02wOdZr/wYC+o6gb7ipgl5hZ3AiiDGuyx4ukMZU/+O3TIPwfeSa9Otpe
5PFB+tCboqCSUXfZT1KoBF7yENC5sVyJo8BU6gppvG5re9Nl/P/UnGCwRC/f7nYFQhgfdIxSRJlr
mP7djM532TPjEwc68H+WAs1/uMID2hvrJ6DF7qmdafo8vfqkdoiNPD4SxBSS+ieiOJVV+kBPww2a
t0J9DQd2+X6aMqb+3TZjWQURBwK6SjPTgO53PX5B7mycklR+bAQ7sA4dI+ntH2htWzz/xc3hIFg7
g+jWzRRxXsntr4VGqlmb76YE8q6u19kgcn7fYogLAq7TgN9nkOMJiJst4Qv/sgQqotyOHnU7BEc/
xB0/9/sho+4eMpEezvION9QmC2FH3C7ZnSU0JxvWoMnKKf8+vgZEnEddjvrobsQXyimnA5zFn+Nq
W+FfG04/aKx7PLNTnRmterQ/aZuV9fzVphzOnfZIAo0iDS0DiV3uxgkcKo1ukQLY8ZDz7aHRT180
NR99eUxhBlVT4NWqi0Ze3mPeIvTUaujQeU/xjx6s/ieFJKuW2AFM4Pp05vXLem80hjhPAmu2YRfO
s36KUssSXzyOWKrrCJER1mD6gdQvZUugtaxOBK4221iQnYP+PQYHYX6Xd+vlRZe0CgS2wafoHCNX
K+VJkvJ8HNmBCJab2inO+eWcQCxqPQmeeuplvUKEd/i4klbcqHR9ENvlaeJwRh12IrbRHlUx3y7K
L2hGHhpG50zYC7T+S46MBsg7x5YaLIO6Htc4V2+aUOfM4Dv5T4oj30spR8/Zi1ZXieJCgl9ilSS5
HMIlWa3CGqujyi6tfg8KY/RlKvQb6t5VH8lhsc8QkEWGSj4Oqfqx9CGjBh5KIbGKgIYdQceneZTt
uxdg56AK0+0sBdPp3LjsjjdDxQBeE6Bx7b+rlwM5cOwpxWu46HZ7YMMDeYLLubP1/0ZAyveCVgoP
jsni5eYf8YOQIEfdat0hUExkknR4v5Nsel42FpBHflVZyVPTPyZLJm1OM8JV1JXTzMSdqlzq1aOJ
CVxvRKQ4LHPtmu832xuJTn9vBtvizU5F1g6u5EngF6qrzIQ8h1VzjXl43Nde12R1qJvKHzyYeP22
MgPF2QTkXZtIF5sCwpmGzl6fM1NfCUtxGcagH6v2A0Og6YCOuM5/2nqxLTrF4dTA3JCngz+ag7F5
b7eJ5n9PNXxNswWmioyXfzSOhe7lR/mIMvKBaG4uGmNFq1/PzjIb3HFZVqdPPV3MxdTr6imILFdW
cgrx5iBkMlqKQIbraEXyuyEDLnQxmDKs9pxQD5VuBJvTQUhK/xUJG9Q8JgGKZbQcV7vhM1no7+6G
qyKRB88WNBb981JoCC9/lX6vB2HBpiEPhnZSMqqCulxIlZIuJLCfLJdrFJqs8+iU3gEIyFc+H7Ti
EmSKtUX1glMzzElOZaVNE3+FrODzhYUT1VW7qEnE8UvZT05KWkIxSBz6xhLg64DWv9MyaoNydsTY
qWthE5wWevDbC0irb6SDZhdOGGOGMVofidOhYY+bhT5xLuvYS/IHGNhVg1nYChkLOu+xYx5BKdKj
XlkjVtIWiQUxCWKHJzLgwF0hDqBSmaJeh4rDTPjf+iXGLfEOoJ58gVumO2Im2xMD1wesIiahodUz
FRM+/FmGDVl76vpIjmux450N+NKbTC8CNo1gH1R9tikN51fRe0p5K/UVyaAt7b+MxRgLw8xq6039
ykOpGZfA7sWLrc0o0CUABx9n95JafO59ZrueA+yIlXL/tH1CFH13SU5rT2PFNuksRk6VNSIN5ByA
L1dqdr/GbHIyfzOv4UQMCnBdyOmcaZf5TVMMrLfVO4yQ4JE5BvYYsooeeUwr9OOnvZH7BhCKU1ZD
xeGY97o8oWq7LFVvV4kG9RuXvk7ULRZTkVc5dy2laHM9imEwn6gHSFDKQl5Lb7o/LQdqAFMfbirk
CKE/CLSwMIOyzf8CJUyPOjVqeW54dg+g9HrKvG6Ec2ndfZUyNJGX8SHRT8zdboqHeXM4LX6FCLfk
b+w5smldTma6qplIvV21xhp4yskaVvq0q1GpuiC8UMpJgBGEDw2jX02pNbIUrP4sasK0knrOJGst
QenoXBJx3IuoJTQhaqx3WVQUE/TMzLmV1/lpl/kZKctZ9+vdw8gRPE3L672w7hXoRuIEn1yPYNrx
IRMEh64tosrugchlVdXTscV/ldTqzI0ShhAuouup5Q5x1h8s5Cwm70LAvr5KOBr25J1CHWvRUCE5
PipI7dHHM0jpJ8otvtchm/M0w4euPeqlOtWoqH4PQuFf4I3GRHnKwagNwKd1q4FrdixniV/VxrDJ
CV3eS+CC06TJNo3jnkghpXq+Uqh/0OGZJWG2tMkNKkz9uKvryM8X1Rxhh9OQEd6DBGZxTgCp1+bz
cRzD7n/3nWdUM0jTc+rx3wmKCWGf7QyqIb8ZzC2GRm1OCv0AFwC4b9ZKcpBjZyBCINgycfYoR/Rx
ebBwLqkVufCZR5CQOEZXvCUSF4/XMQWPv3SPJHO/uQY2GccelzTH8/zIGJ7eCsG3PNarrBcmXXaX
JPXtyiWh26IrLYWQNW4gDkJ2bJD03AdtM6OPb2gBjCS8ctIeupP7YnX4MBaDZA7P+SpsHdyqKvYe
DLSHHIzbTJju45Y9eXMfOkTWA4Vhlnkf2OhPui1Xqo6sUXWoc7dVvL3DCpruVPVMDKPsy1aGpS0V
WpfeshG63KzeAWFvrr0cT8kFQIJHwyDA7E0zxu2tdA/eCZNPegPGd4wh3nIPpI5idMzkNaU3YPUT
6U5tRiQlgnpVNAwBnbN64Cz48vKgptdQhcK/ibAimC6x/Yc7S5pfc5dXO9MJiGBtQQWhB23wnur+
/emJHJtzQDl8o0gVbj9gFN7fXFfcz36HJ9wUM978ncNUdRp/RMb6BE3jVMk6Hf5BI1H+Ucpmi+1E
Ez1SJg6tOCgiaivDTGc/NdbIB8nyMHt8VJW03P5QAX47BGnc+4yGlSzuKyTG9TIgJbmJ6o8fvU+u
U3W5U7SOmelLT2sxJL45+uqhql9wrawAQbmBfCU0GW3R/bNu92U61UNcNf/O4OZtpkBPRa4dGdfX
tq8evUdnenwn4wDp/elrjcuw7t/h9VNg3X54rgReOOUYNEq/YDn9GnFKYbYqhr4x7LWDB1W56bU4
0ebM/3Xu4u+4yPfQYE00U+ciR7dbRom3jKw/QRgjCSmGFN/CIkT7XGUemb6GhoTfweTcziYX8fb2
sj2LqrZO2Qe3CxgIYwJC20bweexxGsx88GofYbhaRCZp3J/B1uuVPBcerNVzAjzii5cOI8PEL4e5
ELwUa7GNQb3X7J8SpJL3jY/JENbl/J+BK1H/vs1l6DrIbUQQno8E+B/lcFTc6A7E95JICt4SvDcu
4iKvdeqsYgtmK3hW5YmpawmbaysgS3HIgk/Rhl6T/hJAthxSFi7wFqTxyek9vwtbspuntK8Q9jTE
4mLwJPrfyqvBdXOQJyVXcFnlPjfSp7EZbHjeuXAOZ42PEHgN9iBry8ouzLupAEcMcr0VvtF63ttX
JQxaa5kFcdWb7VzL3C4OE0gr2KFEf1BiXGb1eby3KHxR4iag7IQF5QKnKndffPS2gK4TYQKQFa5m
CQRGEJuMklLJ2b434FLX57mZs2FRejg8PuK5eF6f1m/7bgsj0ScFXwvVvY9aPZ95u56LKr2zl4w6
L8+rJqwEiCY0icTY2H01jsP5BHeH8VGe9heMd3tRlC3DsoLcsD3rNPdPbOjGf8tv5hSdvA1QKD7c
dYz1kMpwHPY7aXugMgHt56Wnlfrhyk2HpN7IWHMvsCBr865zSgvhS+CwFfcNMIriqZsIuOKnaLQL
lsvj+kQkb1l60EXDe5EhooeOYhWYOeKpQgX9kZAztfoaf4yFDAg5eZ14RGZ2DmCS+nAhzgCa//Po
q03xx8EXmOcRhkjj9LklIVYkmgqN1ml0p5QfGzhxexI5U3fBXhO0J6VQD7zik2n1lB9NVbR6jqeG
nH8Wo5Z575FIYkA5sysY7TQ/xRB8Mp4tSTWktWVmQppHhjf4OCvILHaIe6jpYtjbUAAluXswVedY
Dd7Zm5DOtWiyyPo6NN67WgrQmHPwvVp0cSRXLWu3FGjLrZ3gT5k1sfGduAli6FOEwtRJQ+nBbnvv
GuSmdgO8vGFBeirmzZPaDm8+meYuxBEnChydjH1BNZnglqRWi2ot4DqE0MOrY+dDa2XlhCN0+MM5
o8F2PdFeFK1ZFFr8NdSeRYcUlYCNXz82CaHnha7jX4G3Z9LM7/sOl80qrnpNijm+FRy7y+pSeqbU
ZtFSFXWNismVjCWZDV1G0zB5MaZD+9C/BlSWkhg8rfP0hSkK38oVbqBJoq1Mb++5m8PxwhuOHKXW
Wm2lAa6aGa+QNXmD9vH3z0F5Sn+csg/KM/X97fbU5BsQ6iHxVIBzQR7zzQf0KNdRXcgDAvHHvmLN
CbDWoJHDRaDyPOUkAQEsb4VVbBScornRpOXVklvpnBlUr0drztRzHiAjruvs1cK0d4PL/SPejFeb
fp3Rdb0T/NHDe9co2rYiRxhUm7M5pvYhamv5XvDE7kybLS3l5SuEAs4vFbH0eCPLuDEaBf7jXBLP
46ti5wg4Gwj8VtfzGxWF/ptTE9lEvuC3Ei+0xFlxQevSyZiKxbiTTM8TfYdd+Eddm61nvcM3WroM
5rbcRfCL5urj5/RKe4nNXaqjfSnqLETTosFd/jqhqoo1cchAg+0TsWfGJKNbcCS4Bs3WRbJdKxiV
RzQgKeoaskdMOE9yET9rhqRB9caj/9FfPcp5mBXrFDHdaBUVfkXamJjz0ROPQH4f00RSd88MHtg7
bwOGQgLo52nzgsxGJ4NzoyV1nK5zlhKkdtAWDWus1Vp/Awp0Oq7+E03ro4cbIhY4eFXaaZsjb+E8
tO4+IdogeB7lchIexIhAqGhmiWsAVbZEV8hHfKOtHxRBflVcRDnL4Uvc2VALn3wPfeVTN+Ov2LN6
Pd9sBhp5tCcADOXbOI1oNZtaRMRiZPKtgS5KOx69A+wj7oMigMqXGRlbvM8DOlphb2ls2Zej0gJx
A8mEh1KB8E9HjSGcDWASSmYm8LWSeTb4k1VXGN8YV+Z32C9RoRKy8UsuBWtVw3EjxIbCSI8CS2Ak
eFZF5t1qwmnnz/yZs1g1pI2LEF9z21pfOIDPmRkSNYDTwlDiunTi7RSr5MzTsZHhL8XlKjRbAOqW
G+jqwEthguldybF+2xM1alnXKxzF5Q+zWsI7kZJLrLyAKCLvmvNPo6xRh2hZIQDFtK/HBJX7J/eW
f3wqDuCrKU29ZXXggHkmDBB57pjs2TUY1DpgatDRHbIrMyyuify65OFiqX+0n/VObL79QWF45DLF
X0/f/yQpWrpBHj9NIf8ZYRS0x3teAVnmZrtcd5EsZ/KGELx+2OvZegy9u2/t9HYz0TdPFqjGusBC
gqoOP2nVem2rb8QzSYcku4PoInPpZ4PEpaQP6guDu+MFdM2GTHoDadYkMluQ+KlbxIaz9UPDdGLb
UwqgFQBwT1NTTH+dfoBeP6VdGz4W5TEb1MgILdfV19WJhF8ZGTYJen/Y9aSGUKuZ7AzxqohzdmV3
+JR/3sTec/A32w6wQryHup0o4sl0Pkrxuh+vGM9Ry2QBMn4O8fJNGJUUWx3prz6kOzXyLjh8YQZp
M9Cxq/uCXMxIZyKNZv1VQS96q+xRCVxv2t+9WozVwLGyseTPtbGUTrxy79yNn08BD3Apuu5RpIel
cCLjFAFrRaTrPxWdaMjcuk2NodrpNOMwbcGS7nAjQ8UtukG+aYQjhlVb7qvli4ps29s2eMRUvzfS
qNyESfa0Hm91d1DpbzJ95inwXewMNc9iTHPoKad9Gr7m+8zLjXN5J8Wr3/SVNwHlFVNLD6tUYxr8
rG3til7sIYez0i2QskV11QTX5oI9MiXRteq7TkvTJkOKTQQRBxL0Rid149Smq6R3qZXKLT6YbsU0
88EAjVU0xC4qwPaaSMfcDnYl0IT8GKngKaUXnY+A0Wfze/13qkCHY+MK7R8nIgTxpbbVtHzEfFFx
4fhVpzdoH7AmiUxklrpFSXuM+aVkcqyJcngoupz6m54VddkFrMwGiBKPAeEqNaDSj1XVFyp/5mHZ
4WFjeuy7D8WMdPXmtA9FP/QQ68c+pOPu5A2PVeJdoAWXwFV56997ghGKshakerwJlPlxXB2wOSFP
MLkkiZoYq44T7VZvxFI8H2uZLsRD6cHmjKtLJ/xEfSZ97VT+S9f9TN7t5/DCC+9hGLHykanWO5tn
XCyPoIx5dBYKwZLJqYtYzKGw5VmBXZeIiseE4fBbfyBWWqt2E7D29lp3KBzXDEtwlYyQloeWo2yT
V9Zxf4JiV++AkySAyhFnC3PPn0CamJsPrvOl8y+uW/YF3FvwlU6KMYd0cdQBySteXWQZomGaJJbN
/4QUPk0m8KQVgQfisAWTQi5XgX+FXEzQl32JaMNMluZpgtKp9x0ZUP4N3xyabJOTh8qNrEIHx8u7
uzqXweroubS2snMAM0sHwDhHGvlnbVNNHuR7V7MhUllrcuT6SeNxezinYqvzg+MNuH2quTyilVYB
jLgSKOV8ZJRoHPlyeIIyIpnY+taDWAXjb2XbnXLpRsQn2kppteDe0nuAZ5KGCeXBN3taJjkuaOSh
4ZDaDQtzVosLXp4kX3rLUO+ZwiJcHvERrj0J5BWJG0aQlUvEgg0Phk5kKnVgcyqJwqO34ajMpjuN
qDv8KXDg7WVTcYXebinFEaVfn/UuZZ97c8U+lWBiCzHgMLeaYY49mrKnjChMvQreUukdpJfFHR6v
h2fHFetyzkHtvZ7H7RuCGoDi1UyROc62UozNgtGuSAq10wiJgfBLGzZtgCwVkfFrC7QN8z5PT3a0
xqNp874pnj5DGS96JLLLFjOsXh0IwPF8vTPNEcfoiExURImtQLIa+selNDk4WExGePTtBVxH7B9b
8Jsv0+HpaJ4QsGiE9+xj2CECnBoIXWhLKTKI51eYVfD3cqXmPcAgTsP8jVRN9BnwkySN3cx+VXEF
z0f8vaWGY5IkqYqZc1G44YbRz2MbZD9T9e1UnUpR9vQIeYdd9NLHWdmiZPL1xWkplnM92e3ib+OA
ZGZTd3UEj9k/GJKH2lsOrqHpNakm7EPqStSu70tb7PV1m69WzUa/JGg6O9jhmUYICQXej2gBUz7j
079jhZOSVnOyjbOBWa3poarPItXpBEu1+vqAsoi+xTw/Ayp+KMvkKxQbjoQjs+j3k9HrMWzVnG8w
bAL7Uredac1y36uJjmXm3SaDON3FLpuUc4o9kG3a0T3jtf2KWYJ31dyjiVcqPRlrNkDYGUmbgCwI
6e/WECBR2RUEaHmdE4ffbM60GDq4SsDnFa20pV3McSmMofVN7UMGncBx4erkvlABIZ5cYD2L3J4H
CQJm/Mv/XXpUVgFDKhh3N3vIJhjtRarlDj0EWZOZBlnIJ7wvOWb+bBuizp43LdLl2YYzvAt8ygze
VAUKFmuuDrxFeDghpsPF+zX75PyFv6mBwh9TCe2IgiqN6NxCXvq1FL7oZCtHlxSR8sBGQKbaJn2W
pR6VoE/U7xmPhZ3O3AUgSmOX635qeEAA0dEqIhuTCI6OGQ8EWJ67QPkofgYlivNbc5KIWU1oD2Zn
EMJ2ZFgJUbKSNw0qcG7rjXJUArGG1sLjziPK560n71XGrAyqhooa+GStwEDrgdE3viWejO00korN
daAtZ7xLJccd/hZtbeRdxtv0nnLoHBL7SmQGqB9y115AVn3tQuj8i8c/SRZPRFpNGlv2NiPvvCiH
e4ddWVLF5yEhaPFZpznxHi57VY+6c6hbL/dX82NlD5f3vmYpIXGWcOjMbuGDLIhvWEj9vc84xRf7
wflEwjWXH+TtczwRWp7jxeCxDug0i8x9IUu5zGS8EvFJQKEEqY5aj79tSFkHR5kSj2BBtTuwadsc
QDuvpHCNvhV+W3ezw9y0MGIpbWSnZQ752zrixWn1W4GvVYOEbjqs98VTuTA6Z9kweDk06G6KWPml
Ntj/kAw0AN1MJmqZZuT71aixu40josyzKISaGaKiKZG28D/9dmDBn5C0lViiZ9pP0x/G3rChtvyx
RmGtEnuqmRSnycwTV/pQeA+00VEgng2MUaCQ4kPi+qxag3v2ViDFzvZXNngQdWOPiaWP7K8B+fhC
9xVtFiyk2Ci0ie5SAcRgiaf4fwkHcbHS9K/sSu86qfsfgcr/0u3F7pSgo1nP5mzHU4k1QkPHXp8D
ZA9emrPD6wtzWivuxgeeM8QMl0Y2nONW0/fsqshz3n+o9BjBParh0IfgCvkpaQbIhuYm6OPr+F3R
fP+4T/1GZ6EtwkuOAXkwbrYrloqltfsggzcRJns+eoXh7yyl+VlszaJCACnSTg66pDEUAGtGdf8n
WeBGSRaLDPqaUlI3nmD0w9RtVy111dDG9uBtIIURxtoEZ86EgB/2PhDw7pDagl93fz3oywMahOoP
vMN7JI0ghrkv1+4z4Suv78VwxvTjjpKGnglgrf0EbMNP2BsEPPYpePVi1S/wnLX4CSEjDJzojJUs
3lYN8xm7NIDonaByRYU+hPe1++4k0bvDIZcYtX+/amVwBVUrQ92Blbjrge/dK15iuyzZYMpEHmG0
KxXmOdftgYRwWyC/3e51vuoniPjmO8JaJRWbMMYYJgRbO0Q9qR7fWLBJJ722g7werCuPqDyoJ7gH
JoIgtDlNby7fy3GOoZ/9BVxILBr6hZmUZ7xBYZKQpN8P4BXY3QZSCjQ/F91nEH/As+yFofCkwBDn
I+NQy8MAJuk/9s0QoKQk1y6rFX+lk0UcMwJ+mZ+TZLwipWisy+nQmhJnUMfh28Gx6Xqvtf4fqW1U
MqyHXzz5rX6nx69cYWrCAnrRX6Glg1Tm/E/vKaAaOUQX0E0LHcbu9DRnA70/Y+yU86Zl67EA5gpB
k1akZH4i6XiRGjFCzIyKgMZygCJ81uF0hubASwAfftquFCwTBzUVXGZHd1T7+uCtQL8YTOb8vguh
WicxEEXqijlMdA0uVV5xIkvDZLHRCFSebhF05HD8TwA8RPAoCv0diCY9RygHlCzWtKrE6nJqjf7d
koN67T8LP5yochmPp5lX8YD7K5h7B/1dAc92MAcryyMWqXcmZifOybK1cHT9GDVqKnGKWg36y4lc
yuSe8f9yxC/6cxbzUga7T5zV8Q/GWI7CnFawTTwYKgWVh9BS+5ipv1/6YVID1uwubWaUEN1K2tZ6
JrLI/Cj5rkw2KdGWWG86gKoLL8fBB1ZtcYkxa52rGzboF8rdX2oPadMIbMtUzZ0X+l1TJ4YSkiUW
62CmJpMKSOf3uNK6UvH88LKSSZxx56TDejs2UPL2Tw6cWQuuhnJG9rD8ivKcoXSSMvHSxJ0/wDh6
1Cp6qCnnyjCQ5+dsHJqUEhVtyWt29FQKZZSUbfx4FmfXwn9bWf5MLDWxdrgirX5RcqmsiyA9TUaX
NbZtPeuXhliUiluiyzzh7PzY/MC9aZe9Oq7fpQf/C25MULStTJ0ZrUdYGEx0L3u6S8dMW1E/vHgT
ZMeb9nKsj7YFe+GxFyeODjT6sy9S2P5AeX0nNc/ymw7zPLRkvButomqwRK7QI8KzAV+kLYz0BshS
vqjnlhoPHb9ET0fnxkjYVAY/oFU8m/ldpvbzl3iewuUAkB3/qcdnZEoAs+7W1kmv27hC0MsvVyqm
hISzJXYOzi7C5tlME+8ITPzhwiZceN8W6eBT3aAAeYFYs5qGRKilbwakX7Z9Fy4rvN5rWU9uGUIy
sV2iWl3qRngktWsOrdtHky5Syw3tC6q2OJnKOBilBtnXJe4YpS4ebQfCMPv763DLSKeoS+0+FM+k
TuSWkArgej6V6Xf4Vq20kTBM+bfbXX68farEoFLx1or32kmJr0W7EMEd7s6K2RmZgCNd5Sew3Fb0
L0cV+qVi45wUvoS5W8SqNa0/UTG9WPrmly2ANy1n6NmhdD65U2RKC6KBu6mVGMzH2XFEtVfjfHfU
+fbIuZ3o0/CxrU4LGFzy5d3be33Eh8pkS0vBemJm/DOlDLerNdwPdq/lpUM0QYsUAFyZ6tjixvQV
TBw4I83S02c08XqJ6dYi3bTXk8vk6txfGjj3fheQZmPh+F5+hzaJKY/kJHhUpNTHQ2nF6yIHboZf
Ol+uMNvocOzl/OsLMD3eHzAjvon5R2m4sC6FgBLwjGNHHYKjSXkam6/QWKB26VL8Ry9y1bGM60HL
LCp3/d9bYt45xPcQiXBYANH2TGyj0peQ6r1ziyR1nqqkpup61cxWXMomJqNW3Qaecjqzm5nhFNSx
ZpLdiVegEJt0O6x5K45UMtq/CV6jRp6Yd+6KW8xd99Qs33sUuwq4fnFBl+vMN/XmcuuRielHoPs9
Du27LHLxwEk63wtC4R0W0pwI/JyjDvWa8vm0YDxFcFQCI8G8hxlm4mNjRyNMeC/1grYQggRj1yKU
L1AjHMuFwzHh181Z/HyMXpqKn08AUm+4eTlzrTQ47QD8fwDffbjJDeJaoJlrCSowcvmD9Rd+TBzw
1twznUGYjBYlB+RE19uA5x/chDBv7eyoi2mAg/ZwWiKBeEOr/Bp3qjU7KaDRmvb7D1zwPw2nuGni
er6clxd96JbQRi/P5DSGeAWjcNO+Te3eS/joh228RAaacoAsAp6x8dnVrNMUsYEKLyUevXCcTVfB
d/R8+bT8UlPDQm6Zu+dsC3+6Kx9OEzR7pxf1pX1udLR8Fyu0wc+gceVY7cYU9OphYUMPPzq3DxmC
hwySoKB+ATUwxEIzlHvTEcRSpITVTHBQ7EmFqTLxbTer7WRQ8t6fLAqNUouydCydBK3axZL9Vvm0
ZzSQaiIUOFPKyPb+fCj7PkFPqNnkjwYTEToozu8BGKWw+d8eu6eQ6S13t6Qv+BZaznE2rnigndrA
4tIJNQOco7wdkXtn5ucrFAZBMlYsApmDtmQsvgGm+zTTSn6tYWc3htm7coRkj3FOd2kPxPHzfyS1
rBd9p0bXsL0bpZz6Eqa46OlMIS0P10D3xs3zmtGMerCchJfK22+qZcFmRWlnVhfOoOiBQgCRyyMV
aTKhldC/1AcySQOROcMiugwTOXpsRPSsT2CFBHqB9U9kfnOb6vnHbR3l21/DHN7osJf8Q3VDlgo+
FRIcjeFaQ61nSyvwUeCMBMlOxAGK0vYRvFiWO056hBQU2fIDPvE3UbCuBmJj86zImuz/lnSE3QGb
rVWwSv5pE4Tt/7ZDWegAkS9ufVW09AJYXhBUcCuF+K8AiOQr+ewVIG/IX6AjBdRjjUyMI1ko7XLx
c/7bqNpvcN5r0cUxKF4flUFqd9KC5b+HChNwoAhhu2IqSejoummsqbG3ZDq2XDoyG74Ogv+3GMP8
892VTine/tj2JmIENM82CR1gUlvvoQblVn99T7M6EVck9hPd2fsuswH4W7nXyiUrK+d8ZXT0ZS8b
0sKb0Sy+jFrpFy0xtFULAoM0gRpOt6n2TIR87TCw74/md4d2zmscE7QUMUHk+8qTqPd+NEzgOoSX
G32a/dzOFjnIPNyx2nU2lhvK/ogC5cWmyM/aST2qby2KowgfT38/q4aCkLFi49y0X/7FkExJ0luv
u4NWcmtn4sPZd2KEydsZcYpT57tuUTIQd538CCD50ON8S9B1KjB0d6MyOf1L+BTR0oPz0Yay3+EK
NW0h+8nxJZV1Ar1jPO/SXM5c8H9RBmz3UxlAF8Batq3He+f0AJwmOGV9zIwdBseW0KWglXP074ld
zhCmdVYewRbiTxYNbN+vbvD+zEhvz6ylKP6hBNmrh+Cg17k2uoofQrxFu7Tti53ll2+iqwq0Ix7m
OCOoV8tfUismLmRHu78rSzwmRhtSQt4uApxuojSvxCU9TmvxMY6Kipa3zs/Yj71qPkt2y4+Rg44o
EHuopMOGW4zdPWLGHdC/NqUFV+JeUBO8LzzV+5vjBHIV37flh+QjjROr3nBM85lKxttCScQjcHGy
6LONreHMaSZcJy+kqK1fKQpk7BwjO++nRi5Pz9svemfSu0WjRGnQ+XsquOl80NBFrKhNEr65r3fj
Y4EDesrgr2k7XRJjqkj0nf1suJrsg+zySb4yjKUATUQTJ91rZKyKuJlFTDAOsTo4BENK5WhoC8Cw
2lFfnqi3811LM2BjVskzRyzFPoDIdeyvQqgsmcbPmHNNWxoav5l0CZKvaPqLTbNvMq1LuYiK7V8G
v8fbTgyWxqenUoO62rZYhlx0+lqKBQaz+TnFUAxdqL79/WscvClLKI0E61eSBqrY9hvn95Qo2V+t
YZK4lWcOeoEhUTyU2606xRRva28THRqUw2KcZp6V8P2dUjm6+pWnwylraG0Cb4i+z+sZNDReFLwu
8hrxoTYkbkN1/C7qgIXdT+aCdEIS3ZfY0qZRIRG0kOwykjnedcg6R0o2TBy04cD/ehDKgJCln0b4
d3eYcKSu1tmky5cRbwCA6GlzJAbo+xKiH0OpKfAfR7Hm/i7FCsjBTuM+q4vnQQkfG9uHoOQjFOO0
RBzOCRPGpQOSqYsFteMK47CDoAKXQrGDW/P0k/roYYBWq8ZNPnWZXJTaajjhA0Ac6Qgcq0G9/x8N
XZgbuhDs+ABVsyCJZdUJinbps5SGcMV3T06fOS24jRg6iUZAZx9LC5i1mzBdjNcmnOWW8sQ1Dnje
kJThBGIwe5/NaXER+WDlLz5G1/yigyraYpOKJjNYQWhEunq2nAKWqE5IqIL/7io0sQr6wlQH6R35
xV3/mTyC6oW8WdrfA+RyCMJBOvdHBmN5+ddAprqnMhC5BqDsDG7b6j99WVKn+57L21uxfcF6NKsa
VH57Qz0TpmpHnuYv+RMQTGvlemYowEhrENfLh34RUiYrm5+qebDDCiwSAtqcXy+QegMSU4JZhun3
D1DPF6gCEyFTrEWrZ2jh2JPQ+nqAkmzBw99UKSkV8f1b8hqLFEXzGZ9SANYP1cv9FGENv4Zipjhf
JUDFzXzabcSrTRDF5DzJsJcV3/JQvQq90v4ZOVqcu2KhdIyD97+fsUawl+EJRUEZSwehY+0c9QhU
o/nqu+pMua0Z0canYPBqxTRT7QyD1Gfs9gH6ykNuGcoAlI45j7ACWs+EEQeC64d3vfqlEfRVdwQ2
GlKhv0wW6O3WdUImJqmW1/3a7WXmOdGlbZ2mKFL/L28zHOeJAAV5RJDD0wquTnpK8z0v4xukpHNr
W4OAdlAzqrNq/Yo9WWYAfMazo6dBvoeHyP/CCzRKACiIGkd6asfYZu+rm/z98A77NrSmevhXaSu4
LYTpVQXDTAEjhFwNdWG+NDsa1yselaS0c5VF3N8SFd+tyEHmGx6NPPFRUKtAaWJS0NM5cLlnjhrk
g608PfZmUysixu6r0QXdkGf0J/QXaV1bx6eMdYfy6l3ITqDXsheAfv6eylkcM+uf+0wEf+qiXiBi
T/Ncn66t8xIuRK+nZjy0mfKGLSvnKARO+io9yJ6FAiVY8Q6+riv+UTryPlpkCG0OaSciHMaSNzsi
IVHFI2ipZA3jO1Lc0MZRgBW7hp6rqORYB1Zw8bDe+JsHou2G+Wnw3U0Ko0O5xcLS0zFXwr2chp9D
/8qCgVDiarL3Y4WucB9seZLpfnk/QURP+8mPd963ZGtn9FppC63rKk9K2CYHY1HMtIxnFb/LQxhS
oiqszXoMuoBvjlwoCe/5RHtxkZ7Ujsxb9Nfmk4tQRqbAmr5HoZw3COaakN1KMYBJ+1BVXC77QCsP
4qV5MXZ8v9wbAHLvxGUX/ZsDskIPyaWUaNuEHhJxHf8oKFKKdjX6vZQdY8L4etA0bTVCmvryoLw4
ukQb6+dmzAoDusW4nipLr3sad94+mjw6+zJYl0i2eNqbUkzSAHkJD+RA/9Tv+L1VsnQDQlq4OQTa
Aw2+eeSYlKHLZc6xUeIq1MvoB4d/GHF2jmeGLUHAyhkK8qTfjx9tF/NjrHVD6CuJG0VcEJfJeC7z
/sFyngXu4OerrfmNQIsoZ61YFXzPDb7WPQu75RUoyR8dtVk/HecdX4LNShjoDpggbEoI4d3MNy7Z
48uusotwFdHy+jXHb2DbwCczgwrFERvOlikQHh1zU1T7dHKIQpnhPPrBQS1jjmaIof1jLrdc5b1q
X5svRBxXyl01rVN950tHwevbo2lwEZVB2k8QgZ6wCNlzr5c1GTK2gIUGt9C+Fp3x5wc69KgFL6PZ
85BtDJkEtL8H4D/STxjjjebQy3u+Y/enHilbjY+bib2Qence+fYW48AXM0Bp5eO9NMELkobEqp/7
i7vHBVm4oJI9brRR9Zlm4XQHtjCiriPyghrTeXLVWKj1P+Gs2l1dmoC2uJmlkU8iYFRWzJwx/d7R
nxvhgLJfK2NQ5VUSarz2OuBaUCIGjRT78UCZ7X9JcVDG+6BgjL76qQ9X8+nATPz95KBkntTqUVXi
l/NJYEigGJDL1JcxpRyF7OvgUsLW75S/u6yj6SotJS0ZhN1DJztOtBcUAeNXv5RsyViRULe/xelr
4o7wUsTVCbY+ibTxLFpDEna2EVSoUguxSlDOpiqrsIilPUXrYaAkJRJDoxUwW0C7cRsOyahLoOxe
yrhKhLPPkpK7QHZWi/jkpJS48QX++8SWqUYZsh1gC2aInfLfsD4IjV32UZUmh4dQwDGwyg5keZBd
dM6yHOtwsQ8TXe2efYYRz2fKhpEZmAgpxrzRFXyIah7EWlrpibsnEA4qAA0M47lfgGr/NvymClah
xVqkevx4Pa5OBO72HTMLOaGBcgxGHePNjBcmhtkre27+MZbuUFfdWy49ls3JQ3w3JpgB03UrOiSM
uCtWplFWLQnf3vZzZ/VV9yuySa6dw2Las+GdMWAAl3x3I+Su/dCrwuayLSg1JKZoUrJHsCNiys3u
W67KxZUdYo2u5e58K2u2UgdiMf6TRkaXQHWH1XotF/KNTGqJeNFxilhHQOsBcBZEVa7kX9HZt6oP
5oxb95t1XWBEQWMYX6RVmWf71EZX9/rUb4PPLu+Lo2ckXk0I+BdaJz0TZDzTEhEVPEe8VDSyOn85
RdcsH9lMzOC3n5DbZdVqKiOZoaL8a01H8R8NdtQH6hCTuerVFWYdDV10sZ1TECRW3p/8ahm11ACo
Bos2n4QyaIVEzSBUemKjW0Tc7aB+HaHk9US2VpkvaVDeqNSKSL9DUNKAn12qbSSuvWSa58QNTs5i
LKEjp042d1P8Y7NIdLt6SKZENjt/Emzz5CAlhjL5x481vD6l7souG5wsPFkf5FtduXj5rpQLDTfe
o2mA9OMLcRvFBpZQJmlG+b5kckLxR1ayU2fLFVFjv5hhU2R8Y/VA7zY7rWGJtDGPcQTRe38MB7WQ
Ak7LWkbBiewvm8DD8rllYnJlReLDD0l+v+lvYWvfVTJKg/+ICmDQyQhttONuKg2kRnBRSPCeySUy
bjrRepLUekXLWOEv9/nAhtQCFnaNKAFxLj+F/odbrojtYClAKgs0ZQjFYDg6EBqeC6q5oH32p8TB
lHV/XSTn0wj4JUCV4yv9HLIuqE1NG3NdkYAUbkKwSCiCwctHeqHGwpbshxkkPVd12tX1aCj+CWU9
MGiFZNsG054F5/R0KF2bAZl4kdDPB3phbLsQCp6gHy01/ohY5Qosg8U6LqcIY1Z9iZRisdt2mtz5
2qaL455ERRlWLWOn/Pd8XZDIR+xfPYG+OqkZpuhwxWfXJJHQWmVldKLDOtdbdiIaclZMO3Vs5Rk+
WOJ8eT4JBC3ROlmVZM/zOHOkNitpOus1pZ8UpVaicC6echu7gCikKdF4PEKaA4d6KSDdw+qpsQDz
70J6eSNf2pnAZCFQJsTd2i8TIjxI6UbCCl2yh2CCJPy5L49GWzAmpDYz0e+vlFyAObuV8muIgn3w
5Zxz6Xa6IcFAwkybfIoDrIGahpuzfhLrea6rnk/H64XRuhvIak/zpzmPk0xF0BFPtXwkqRtJxWxe
wrlqMKCEJBgML1KisoJXk6VKU8dpf1/cjCOUc1cNOByDnWifSDQxjWIzzWuo8Ga9aCol+jwKMbF9
nFQ47DXpkZu/L1pBi8kOWb9TpiqDPUA/FvUzsj3WxK8isocbGtQKND2xFwpvvoCoY4Z0pJ+4anyp
na7zpvqT/tUatGO7uhr9H3NY9kio8yLetoOOTwnpTltwTyqyqtrFxRWSEqOhIFlpQH052HCcZ3wU
BOqv00MXG4+x4CJYAsmy47lBx6M1O2QexXuUv+mv/KPCmPGSPkAWnR+tvT1t2S/eZjF/0gMiMsqA
cMrXVBaWIBX6VuazjqUEUzcUQ2C5TNeqsekgTrT66BWqJQfwmvichhqqpWJjCrzoEeZu6Khhn+cG
517BZXcFCpfyoN5Y9LJpooDpSYCu5Ly6CRcqWPY1+4eoxjW9/Z4b6Zd1TXmkjWL07I7z7XZMELq/
GR2CCjO6wDnUUM3Uu1/4jC6wFAjXM5PO54DA0zSnNSnC7RcrHiqN70cjae0CTp4MKud0tbIgScDR
T5skDjRKBWElChxo/5Y6imgCo7eJ+0RPRFKs+w4FG4SkOAg81eDFrCwLZWSA6jYENwHHtn1ss7Il
sAIfNliyu/z/5vvc0Ipmswfqz4ZxFn8ozBmWpDu2e/z7vF+WLZqJqSuuzbZiu5TH9ZYqsp0GX15B
xHklpZ6g8RWzknAWZiM/dn5a/ZVDvPYy/sPj0iuI6AUu5P+oV52jG3XvdNelqd/Ktbpxf/kevtw1
Ugmd0tHpEf1pReGKkD0R40v/0VCUv9qznMP0eVZU2B898FLWioX5F/7WLoTSsF3zDZjlAoQeGb5u
UXbjjI25JTNtAEejzV3M8w6VHi2f5bzIkwbBRBSso+8t4Qj/2ZW9zawkhAOyDnJIwF3iaYe3ogy6
Soq0UJUhpT8TC74wojNBWzH8j3DjOnW9My1vnQ8ixOXxfrEJCPEdR85OsKV9NXngeiL1I6J+wMsS
0QWEVvHW8DOgm8oIgUDHZMqKC+l86iFjbd4QtztfMAQ5IH8trVHdzCsoaRHGh8QbBDSnuterfkWb
nxUh0RPYulrRcRWXtJKJhdj2+JU+1ccU3zehpgJVMflAr9bMjO0FCm2heFkvdxHQWQjz88CfCbMU
PzHseK02HRHHy+V5BLhpcfe5TxeqMYqR5ASCYS9dpG6vFRoK5eiy8XeI6Sb0HwJa8+PSs3mwBHMS
qzOaeK3Fm7sJUhc2bugMqMR19fINMFRMx/+wN8eaAapm70H4U8zfCtKVGK2fuV6ZMIqC/c/J4k4Q
wbFgxYbvNuVCuBA0KUBxoVS6lPQ4akDutk8Yj7+yn8d3gqzMDwSTEuwfQlIu+VrZBR2fSKT+i7h0
Ae5UuGSTqrOF+3IFdi9FCMw3PIDMbl+4xhSO6OJwRg+5UybKNaD7/00BUiOEA3cNJf/3tYTzX7Mr
gG/C+WDvNUVxge3vc8036zi91x/+ppc2rXyJS9XQDsmbemc79vqUpWzjcS1AQLTrTBgqIw33gKFB
H7fpFgtBdsRAhE/r3ilhSIOmJlczg5Jo1MrDqjj8TC8RPx/u+g9qIfibN6Yy59LLQ4X9nilM1ymD
vfKUpmKUkulHeqeZDg+CapOSPxKIuEbh9dxD8K5VV3ztZxcfKe5XXelSFSbblRidRM3/8dM2QJ9M
elK4RcZw/klSduwLlAj4y6SFHos2uQxfasG3H85ol1yeVqARhlyB3Sy5F1t4M9PCQrgI8Pet0TpH
DUYR22bJGUF2FaAjk8PIxHCm8T+zvhZN85zTzVDbh8lyGthMedIGL7yxf7D3F6PkO43bHJX/page
VEM9TtA4Pvud8eR7V5L0hIXphJnFIzPXGLa9q1U8jk/XfRrjesC2ihaBCyljkxsCCJWPRp40KEwm
uIIxYuvYcdZ9327lvYBiNkM4RU2ErTriKF53i6Q7gANNiCjeRx5Y33SqgKlpQtFss8YzxiLFECk+
9VgKV9K4IGLuUIAMe5dWgKRGIxlIsf/EClFEw3mQ48Crng1vACZSRkEGSDdfxtcfVYgveOA1Wvjs
lRwpokfjo1XQ87l9g+s9FfFirCXDOG0IeeYoWTZSmkdXX5hSyvEkpASnJlQgZFZFpKyLlThA1kJA
lQM3jJ6OKZrGw/6BATjPP39juIlPmJIe3xLgxyEGJ3oZFy+AYVGL0hfll2wZ8ieei9M9cygn7XK6
XfIWxhdHhrflP2aI+POqe6NLk/QL9MVZE+H1L4GnYfxhFBQAxYRU+P8Htj6VmrToSS9c3uMTj06b
7mTiJkoqGPjbM+doRUYqMlhpQglq3YlM9ZWDskpAbLMEp3eeEv3O/zvxI6zKpELvZF+dsxnQHfNH
8TVfJJNZMUqxjA44yAffcJI4hUhlATy4HucWRodmkLuUJt/Rtjfjh7nO7TT325ehjEvXMHkf+zYg
MnDsfhbKWMJ0SWm9VmDLBQ+6D0zo4/1l+HdrbTKdd8lxIbYljhYYzYeYOj/jcLWQJ6xduv0JUDPy
+vFZYbuGfp/v9NQ+Pj65yC25hs8+f5QIFtuoWlDBN1UeS+9CT+WYEgyfliwp9SQ92OqMQSFFW02X
bgPM0SEnhwyvTykpFODg7SWRO7Xow7qFZvkDOeyxAPpk9kDlAIf1PAYYX4qQfgoOhspOAs0nZptw
LKFr9XVILHchrivttaMWFYT56FlQhvq6po99o09FL3zAlEvb8MZ447rJu7jElBTc6x3kri+ktDZ8
zEcdFQDqubw1SaiBRUaEZd3B8Tyox7elJo3xDvfVQiOJWV+pDNzNV/toMogmOYH6p0MYtuwWvIe9
50m6sL1Bh7TV2gigkL7NWzuRhRmO/BK6bdzB3wfR7DshhRkWER80cQhobFajXkTMenETBsI0VnFK
HUgjNkdkt039Rc7gCArdMRBP6eZeDDNKuk0NgeTqda4bgTkd64ZT9JuzznELkmuu0ZLarTFMRInv
LG8HXBiU/1R6H8cqQRN9cvzs2sB7sIfvMm8FMVrFYmFqHVaWeMrG53wKfbC7nO/FrsPaGpdGDf9K
JiIITEn8i3FRak3bz0ci3sVh8JMLetFbMXdNtnbf+y/3MCGzbNyNFEs2dBvEKNUtFX4YFJsp32kY
/dG4sIehkzfntCYuaDEdOnSCuY6qNbizz7pIJGOXBifDITa1vi+0n7nCjw3+gSbhNSn7HUG2Ah9Y
QIl+bhpC+1G0FrRZyCgaVsOh7UegMqtGx1CcGZd7/9KFonk5g2ytFX4039Wp5rTYd54RcgUUwz8h
gM/mWm4h+6EV8O3iVH6EuGxLrXHV+JbnHiWtKO1q8F7bemfGZwWQJkcT1rtZsIhu0mb+J0KtJJ/u
yGyTOqTm4kg1j+m5Avr2y2+OD8/iJ35JYd5eIkwM87xSG/IIMiAWkU7/qmWVQU+zr3nNKnekXOTf
89XEqK677xQnlH/OAnSY1/h1USiQmVJByA1fU9mKfWU0WwTqVvouQg1nk9vgQd5KjMMqDM6RIDAZ
la+Fm0ZydphLuvR9/cuV57Qsan/9H5SKOgy1tf83u4DLMCdD9HSUweqR3bCIOWOjrg81RP8s/7XR
Zedid+zNGmEK9P/+y2TBPZ6xaLiykaWRkSNfjvdKDITVpCHbc2xFQGs7Y9PiT9pDlndPY/KEowS6
R5IbDwjv5yqSNu7OlakssXKDnooEeDwHeuOay9FL5kkSOn5BlVi127gKaF6freWDnnOZeAXquL5n
aXD3B87Tbp6uXWJjJNkfdGqrR6e66gkQ3AHmrO/8S5rPSZ2v7+QoTrOHkJ0s2MFd7Cl2sjID2fgv
r8VTEoP/noyuJSCwuS79beUmNW6znzyKkuwv5YDtwb50byPi7hL6RNVf/mCVjvrETzFl7JZeOyEV
NtON/TmEbnT7WoMqCTfxosx8lZRtIIp4yJKtLEox65L8jglvTnsglH+oYlU//ZkfXxU+kRnLr3MW
RW+zTDvhCd/Ne+wad2ug8pr8EtU87V7cim4WHeaAFQScLFi1eRK2k6UO5BXP0zPwKAirX00AJUoC
jknS6lkp1vT2SmN6a2W97LT7Maq9vJjhyJr1vlfzcT9Z7UzzZl/6VQFlNIRDWuRQiAYrXRzdYyf4
Iz6bywXNdLUQbr55HNZFkhoJMmSq4AuezWro6LFNk0iXAwp7ymkMwtFZS++yuiZVa9ut/EQCrfMX
J5PiSWI/ESk0XM+Qx+V3yLsdwJo4CWbkxBoceYkOjxu8QNvn/LQR63uQlkk+9u0RO/9KCGe89KUd
yY9oHUF47erPIEt6FfLluc+mEkIBCxD0EYp7VBAcRTLFvFgaZzYgCMH5vFgAWpiNvf+T6XTjTbw6
kUdTgOHM4X7XslNxp7/xxSkYMNNPKAasmBNfmucKGixnHwyW1AsI0zRbznO2qyrqEXF+/HLXuhfa
13oNibslfOH1F+EVF8KTj+tmigSpC5onvQqxNzueQ1dmK/S/IdUqo409pMQU0fdKGQ0EmrJkwBoZ
C9dKx4OztO59+5wyvvBfrK6QtRzDB8N5uJfv8EPjs17syOchfHBZFzh6ofgjBmL7khvxTyr9wjCm
yenOV0dVmwTq3YKuh0FYeKDzzGuAK4JgKQ34FmkZTJBnJqA+lC+uEa6TBwYociZ8SLkutZ7/y5S7
Jh+rRROc9zSDKbEIM+EZ8uE5GYUaY4Qr059zUq7gOkKqtumf5vxvBqbTVLK9qNt6L2oeuDVvQcFi
5KFZc1OdLW/sFdckw8czAMwNisGinetjlKj/lmriNSTyWyOzmBf14iH2Uhn2Od3sEXUsVUzb7ju3
fgdrtN7JTmPavr7wubxqcGioDwifa5SuHfXX2Rzk7hyjcOMyDNbun39PKAzZOAUCZxMnqL50c4yh
Pja43mvQ6Elh/F1oy6CsoPxCiCTSA4o2mdLWSQQqTvNPe5ckUQU1TguBEy+Lxxa7roswYttePD49
F/0jgw4Loc5YholLti0n7jLy4nc2ADBvLXU+AekoTSybu5GKIivrM9hzrlmc08ffUtA24Bzxyzze
ufUX3YX9kL5CkTfPS86XSu3bGX50/qUJWj8CqNn+4SsMDlJwhqtkdVcHhYWAtdD8So4TjwXBTuBZ
AkUC0kdZ8VqmSIhZCsO61KW+iRxwgLB8PD4qB5rBmBvhmGJuk8XzdXvNT81Uxulxpj9+hUXdiAND
h1qTFWiFFFsLfGw5E3KhNZ8DuY8JECZWwK7g8FjKxzE22pmDrIBT1blqh/mTDgUeDMbuJ4JVZ8pz
RLzd6YxVz5rX8jhmU7gK4VCsbvn26vNFZfACL0F35PEsowWBEMgjIBsr01qc26O31eiU8limo5xi
rCPwgkKj+uuKYu835URt3S73cs5rgtDs+c2iWKpEhd9Ne95bu1otWDal3HBDLOyfHraBahdSSTxr
L7vjcuT2sFDPh7by/N1SLtw1LVDjwTBRDUSD83xYJf8PX4nB37OTQma/DtA0/3akMzFbki2yisSE
lHg/8vQgz9QX0h6pbo8WMaT/3qghGDPOnZWzYqdIGHjwEI8NOv/h1Gez1GEexkK+XZkXofAd9V4Y
rhHmK8bAjGlvJY8JhSBeuYeX7ryIkxtNKlqZ5deg3MgFDeKJ3TOlTG0n3O24cdEAhWDOj8LCEFPV
gfF8uK1ZdUtwZidhv8BHwGL+34DZDXwUtiDawGg0ROCEuA9nbs6N2O5i0j/OY6/OMEST+hUpd74z
L5WQHnW7YMJBI5a24qC+bFxkbjMLj77EVU4sX/oC2BxctbpXrNgFzZBgiYkGcMTYf2C0Jr8nNiIo
wlMyJs9Llr4dszIcqtnDh5irgRA7XbHxlEob7DWGmgB6slBNeM3yAlRKcfsSRveSgeuz4+dzBomU
wvPX1OBeb/ftSG1Mcuj9xVsenwcRrcK7Crjvw3A16Uujq0sCBZMGHmfmK6tYQYAhwyIcoWf/glNd
cVUNNL6xk6uGks/YYWhCoDlBxfXRocTTjQMne04HyExqJpUmg4+5w21MTPlaj11Saga3EhOz2UF9
v47hGORvaz4qw/QOcatxIE1JvX+5Bh2LzEXMIh+ZqOVaccEG4p/RfkDRD1B8EQDrBox1MTCYN8AW
0XhO3hs8CIWthqlEduhjvC94bIa/Q9e/ddyKZalOs8uXx2gM+1WRv/akkglw/+AeCQZHAVCgoxlX
Rvpz9eqWch4hMYCtw9op6Zt7ZB2gKTPR3i0CSKS3PCx7+SFw0bejfTGLxKT7FloO13IFLc9yyC9P
J1Me7Gq9RECDwaj1FOQlZW0RfCU9XKr8VeaMJPG5lepHjeppOK9O5/Jc6toM3aIBrjLY9ysJKt1A
GETNcR/C39u9CKSU9RnFx30WMbAD1jV163ZvNng1GkjM6PxAROtOcKLedJcc71bI+fWnADFTzTBw
wXr6PFk80dWtoHjZMrWwHSY0as7B02M3yINef1ElGn+jbXsa6QT+aDma1BFOJs91FqZ+bOibTuHf
KDaHF9n0r+Lcup00JX26T1zDkH+vlTdcW9Wh3NQEIX+B+5ml38Ta++aqJbILrm0NXTWV2WIyszfg
mRyvZoNX/7xVVvNQKYZ1S3ZW1cxQeCbVf7UYtfpQYpQVbDj09t6dyqYGh3PtegMaczo3d2ddRhfS
ENuS99Z/3koq0A8EjZloV+An+IeGk9fYKgOjVt+5PDQ86BW/1jC6QhZzmzo9fRci2oaLbxprPEBv
+ZmGnA56SBcFsJhJiMaWPB62ckm5fOm4FL6TAkvqu/EdRrv7WVrqincij7guAOqdivQu4LFnGJr5
8jUKq9LjFbGdNlqrsJCV3SObwd6W2aBeIKVkbg6a6blEmJ8dTB00RHcoX+kfunZYTVnU23lhatrt
U6GjWctzJjC4cDogVbrtaoTJu4R6c5Dft73F15tx+j5wd9p3bCR8c08E7tqP/fuMg9oBRGXiNyks
a/3Sa5tLEbYlhtkyzmQ2ilDi1IoH8t61hLpoXL994ZZ33eTVzjg6DEg5v43/FNHzELwFuJp3vZ3r
Z4rVwF9cjB9mQNw/faqXmEjPD+aEFVQFcX1YxeccOcIsDVmwpTwC2H8aST0C1nXUXIMGbOd375rm
jBhR+ucdmbk1RQVsEDVGEJPEki3rEVq5RxyOryfjf3rY4hEX5TqltxcXveUqerq9DK4kIEu3tifd
lb+aGrTDd+QeaCILbgxh4yamVAmJTeE74zl5OBY37hHpVzG9sfRf0ztZOPcLEXgBFovs3bzOC1no
Tg8zVN9vXDlr7XHGFM0cWWcDKJtJvYeinjY6JowLUDgWgdipAfRQXSARy5CL1xKrvxJ+oOXT8R43
99xz3AZNIwbFfD/5QDTtqf5G1uEZkUaSsCep1GWYPu9qD0PXXaA+b4A598GgQp+9gVlpDmplHZrp
FANay4Uvn0xx+4R8Hh+CqlxTW1xjGmoYw06tFVmPaNdFkrtvQqp/rBKd/1WbE4TySH24lrURRgKr
/Ww3JakJ6RwSLqR5tAKTK/ztzM6iftAWMB/2WAfdYSFqe4Y18Ps/7n4nIqKwvS6coelH8ulNW8Aj
AT3yktnOz2VMHWa9KP3eRmg9698YDMvcKwIQtFqLOZsTo8tTxv9QqozcZOh9Xq97U74vU6gCnIm6
IbymRmh605D4VqR2p08S41PIPs64aKW790/5Llu3UBp/BUjnorBgWdhZBo4T6zylWTppXozq91z4
++H8rfW+0SkMxff42NfHUsL4O1+VCH0ri53tRUwbhE/mUR7QMDGCZgQ0sBUEqAZ0rU9EFWkFd4w1
GtpM+yoqqFlPLX963+Y7uLkCcUcgXn5s3NgE2+/qZW5t6pHMZ9gOPKA4TPHsNje7UDD2q29LD8HP
IlD3QEInnPk8UJiAahdyTtVW9+Mr+b2mcLxfREY2Da7AvgQQY3lBOsGONQFsAyPmICTXWahInlaA
u4IRXyWkQcalpklqVGW1pH0U3EXVwI1v/3wHQ7TspGu9tQgbj43v4JhHyJFRBDplLI3XX+p3Xq9I
gF9EQfFCiXtQhq+74Xl3UuwuFeqm29AFF4tDr7UaxKmSx98RwEVcpMfTuWdvoxY/YAcTRLxu/NZF
jI4hXzW5kGwvvC5wulX98Q9qxrsD+V+G3EJjRghLGuT/jWDfq6V/HptxKCDSe8eqkpKGXmIDZu28
X3vCG8LRgOxOAo4Y9jNgk3CO8d+N8CzMJYM/GqYG3VNZZ3IS0RKN5zbiFKysY4LUXNk+8TDJRRy1
gXYgJnHus05dkub23Brm2Jn3y5ZvweXwRteyO0YOIAtOExQAvFYwA+EKm00v/2N+tjamfMumynMN
1Ee+62hqbzQdtOkKAnaJLf9QYXi2nfvCh9nG6F1JdZL1jKzvCEvX5YgXiGgHXy7dmZlVcgK3krQY
UnK4+sf2bR/25bibdZBDibQStUS1UEo04HyytyDFCQPsqisEWY3D7UpSL8jh84geIGfAOWd3gyvD
LMhqp7wY1cqYd8/b6mvYoVk90eLwbIVyDeQZjoU3B/86np3JSyPyrsYCXXN8A2CFZtuYWwvuQkeN
jioMyh/kFqG/9Rmb9fL5hswOMKw5XGOHSH4xy+aCd+KemFSBuUCH+5OLIYYl7ttzGzWfh8H40uvJ
aAZMFcqsQi4AmDWP8D3bJ1Du2Xe1ICTHIKLn3VJXp18JEyXYTowFKwN/2zK0R0cHbkc/Wb0NjDTD
mJXNPpXX+20ZG1oC2LfjsSVc9Mv4olYLm68KYH2L388ClMm9NA1f03FEo6YnzdmswNeGZNq3Zb8v
VfOKaV+YvRv2u5dqUn7EN5LGF0CQuBUyp30KMvWSO5Fy4sp3tYklIKnNX5pEzRbi8dMfxcfJo7xd
5Yhzej+lh4OLkNh97s5VY3S8++0XcrjmjjD2Q4OaW+EuMUTjG0RzbgbNYAw9Cf29kL8csTnV/JOs
PWU/DqT+hkVqyY9owhmii+SnpO5rh3Eqa1hlNjnpsCzOEqrdm2ztiv2QUSs+UXTxoFoSo0TtKoAV
ODXctk2qiU7z/nYVf09LJJl2+e/0clb05T3Lg8NPGZXMZF6Y4Wilj4QG4u5dfmp9BOk3496Ncldp
HrufpvIZcBpMvWE9E/eF+bXXwMz7w6zdpfOnyMzTKEHt5jQjht/5auxck+eYwKfpmrQMMr0rn9NE
ix2ROlngA4ri40Y6uZRB4898hdV92kRZJtYD/O3/y0DiG8+nOAlM6XW3wjMlixbC1GQwYi0JgU16
2+yHdzzmqusbVp2jn/NAcWdmjPBcTZDl6Q3v0d1cjiYFUrLPij9oHKBzRhZ3FxOfvgoaJzP1XrzM
EinMKGgXho7vsyMyxgLEcK+AWCP0MbUs17DVOPtBnxUa29I+ri8bNx5whfnnQJzZXwZkaxYVQ3hF
yRRxQNr/XsT1FGd7808X5i/1CMnnPDcooA9B7xtzJQRsgV8btJpK3rT/0CWBAIaYelZMeZZZ9eoW
sxcZEF477SgySBDuXBjcFlL+emwtqdant1AMUoUVIWANlNAzyF14UXgr3Z/k66w8sgwkzMIZUqc0
RjXCwV3+e3FXm5AGkOImkTF4Nzpszn4eau65m4VTrGeeHd6RjXLH4qkiFEMojP1NiNP8wPNuKdKz
a5vqCyx98NTT0RZbQ6CY1ayTHjaWc8ezyh9sbb7k6YPoj50pXOWhaET4phKfnHFgMJo8kRkp4p9f
mCUGR3jx6muRp8DkndFAsMWVpYiS8t68WYW9SUsLertbEWNdt0cEnciYwRkmYmihABMXOSrfFmf/
D4Be5WXlQ2xKcdIZ1/7IqI4pr0NwQqNFzsAE0t5rLSh4eQOpAYVMnlwCBixtJ3CKBfe/w1i6SJfm
mfUauQacbK7vh8pn8UFB3/PRP8VVaOR1s3Dvsvo0SVct2DTz6H9WGq2SotqWhPjXsDwik2UW0uBd
XT1Nm5Rc9W3rkt/PExRCH/0NLQKWugU0/howKozAl0ixCo2ErFeTMbF4DgdXIU49lqB2abU5Pz08
MnEJUGxlPNXLprY3tvi+3DUXXylIai2XplvAsWvzddkEB+2YATlX+0AL2JdLsP2MYMGko7+dXDeG
6ed5EnAnfbQQjk2hc9y5YTo0AYW3GYePIaCIcGSzP63Jil4RNfkmdLvptwOHUaBJ5EGSCxd7b6T3
3My0F1/JCnldpPmsD10eELByuQ1fKBURUH7EJqkRowUnpkfZmdnjGoYSHqCqoiFTolflGkr6znsc
d2g2hMc3pt7JrD3214fKL8l8tltkwGDPhLaEC4Tk/KIYXxnvN6Yho5t5LyMi4JCOWa4kc+vCVwVq
hghzAmFZQYCLRux4cSImVNDXVdZ87x/XeXhYHCcgSdmQw/+CKDudF7sjQQ/fXuUW4fOAKqFEozl4
k8LzVcR0JK1t1DABwYS9JYKtwW+pPrQTQpMKIysiXgMn6TVljPYaPGHPP4NmMjR0cpHs1NXq4wxl
E0LEC2xxLXG+A5QjbCS4LyXQHn0VJ6Di5nl00PVXeDvYHGYXx0Rpu1nKqGU5lUP/3iPRgHR4EqUT
nJfHQGBMxoqxYPNz/77QFP/U/IozvE1WPTcnqkj1i1cujjRLmQorxruxZB6WkxY/oklRetV8oo9u
o6eIYbZz+0NF+uV1PMNqARfYyMu6vvOIqVeq0ksUvxTgGwyzT/HNV0H2mbLnrvs0fFV7Wj1khLRB
j+3mKhurCNBGW5SYOTmHSnWwU1g/MBQGf0FPinNPIpW3mXfVhopMUTCl+Fkp1q4YuYLqSPEF1cpu
Z4tnxnE5gMvgcF681yK0C7yaTraGRGuOrSvBT5cgotFRWC864w4fz2XLabfyAJVEYtgOY5fiYGW6
g2xi0A8n61aRPARliwSOwvkv4fUBg1BVP5EUYGgffpDJZ4OOTIqAi2YKmu9GZh7luNKJvfsDZ47o
tumWDHGrAyBU93zu3LgnnddYuiyEdCC2xXNPc4QJzQJDtGJUsvZUAciP7SLUZ2pwZpZtFaJBj3B9
F7TWBdYgOALb1LuRUWbUtPEGqy6J1jJJnDpRGjwQNipX9ipQ0+bLJ/ZYY2Fsf5CGErlEbo67v+az
XuFsdOR8wivwo3RyOtT3cMOJacVLP3Y3v0ZT6lnT/I79SOpkwCipAU+p8fzwPSlvx3PWFT4bN8bj
jv+Qmy2D2etaoSIqQ+SiOSezpT7/jEPM52WGgHkJal+bJJXxIST/sZPPgf+u9a2AQRqOylLce9+/
y0+1FgrzM7ht+qFEJr2jMdCYZCBKnkqmBydPlog9ldq/kgikqFBisdOxgjtDtFxQpo1Si0B9nkmJ
vdBbO2uaUOG3b9ZEWl6so2/u3PIgLCCBPqejfP3AU7ofObbZxz0+NaTo0cRgQopjUEUaFOx3z3tO
BlrPraeIMwyW3/3PeBMRidBa4ASNccY1j576NxYY8reFEJomhUv9G1JX+ftO0H0zlSLe7nqfT3pe
4YBjOIItAYHet0bp1x+3yGHIs7vif7xDsmyiLyiEN2tt+waIJ4jyjG66baYdbm7t1UIG7d+APS3p
xKXV8WntzHtFxrwGXlKPgqsyDGBJOuc1CP/ko/4BobaQNRLwMuA6rraOkn17McoP39L2uEfxQcXc
Oco3P70CIixEFsurhiiKEhEkP2+bqkUrp3QzRU2CCxc8sShlZgGyQC+cZkWewMFuZGp0Lc1eKsey
kYS+pAcEJnop19Z3OFu2AStHPYmh4dMAVBJcxZ0jfoOb6rf1YhsFcE4KZ6BOcbYQlKkoMGymuO/q
76phXrSBN5gN3w9BnoeM2c15qcFl/XebGyxy8k1k4LSSeDOQiliDAFQ8uTUa4a7bzA3Drm69e/bO
MbXO6NxMNA08ljQhkS4Yg1aHw8VNfRSYS1u5o0QAXkp4lBsI1phsPANqDyo8cWCUu2UEnScF12Hk
UGygiI0nc1iBOTGb/F8ZCnzBaDlM2GAmECqGMTzF5FU/UkZyUgYWOkDowhSsdN/ayCiH0wnl8ER1
eopdcgXlwZ0BvHmcGXCbamUOswbmGy102FQvwmQ9nEUM2gua0KXwtA3c70HqB2EOALDNQHSnUdNj
x7dl/MucINdPqbBptAJb9tDkE9BAu7NlT7d+bfNAIpCQVvdcnmdHp/Guv0xbluIqWftzjFW5udy+
F8Orh9vG92b1UaVmZnWdQCz3D4xPyL2IB2ssJInLcmUo2hnB5grwGINAyVTfkeNpL14Hpz3hUkoW
kTSyDcRELw1Ycz3ndFEhCd4HvFEn+wzJkdIYnENwSZtT8fVEgFWmNUMpKWCCYGF39Bwwas4hMZzZ
zNcJzF2Nvpw7sJ0VS6yBgPeKBaOGBWzbrJzCIua210SujncrjD5MvubdxpsZuOmz/s8Ovj7dijif
QRrC7YOAWcx8Y5850Mm2WWWwjDDxvvXpyKv66A11V7j++145e0lGde4GGDEpg3hckiUcOmxHMTAb
TN4kteh4x5W48G6rCqP1sCzg8RQ9f4lHMFc1WZ+94w13BZqsHSOm75CbetliEyPuKZCDQfutXR8/
+d2mXncXUDq5C0BoWggyF2wP7wBZn9FUtxbpjT/9Km7p3+Zc7FvzGcVfaNVzKkkUyQSpsgJmu1dy
TaoIOWOPJgjc5moLZiErap2snkXfh1GoTrKx2Ni7zpItcjQ6drt26g4oL8fSZcKplDkuS9DDnEMM
hD/k1H1nSDEA6fPIGOn6uFL4MQzcKuVVB/l5wAIeF4spWaR4i89Pvnu509PPVZXUpJoYwo1m9QeP
KA2cpB88HvEfPPhlkVmzgftg1Jd+14XjseVirnNDsdcsgjnbU4QOgOmJVtnkJjsDqNy+X6T2rAky
5qfrzLWDoxQaYqq+zfLoAyJhW2Gn2NuRXbRxdpzqnZ9JrpsrQPyTKl0SioDfVr9I9Z3oFg2jLo6H
tkIUSOz3zfnIY23YKPvInEMFZEGOEvgMFPORpDx3JVF/HWZOr0aLqkSTRxzsLxgprsjdiReorkUG
WUa6/1rsxanDjt8acLKlpu5qP+n22/GLaa6da1hW6pgTeVDnSvRnXYcLYGUa155aZ8i8LCbXVwTJ
EZ4KudylR76I8InqnWxvatDTBK/SBhPfm7pqw3JuIHGJxvYlEA4tLtOR+fN3yP0vnm/nT2WNIZkK
5chNaWd2tmGmWDP/MgdEPZexyY3f0vM9xmyS9bCkQqk6vLaCvk5zYxaNjcOzoMV1PsWzNJpXjuYJ
gU7f49fNWNFrElWduhsIzlf44pqipzEVW3e2S3zIsSfMAy9yfI6BJCaqiSOpdj0eRh2G/B/+4Jo7
s3SJxpVPl9errOChiWK/CGNyNdkNvh/stKjn+5/YNR0nGvA9rknwukXs3b//ikbt6wf00mJKBhZ8
VCsII4QzIYy7lAib4paM4uxKzSkn0SNLRQ8K+I3YOnk4iirrl6apyuQEEz8MLX6Mba0vqGDEoS/R
cjptnUK4g1Zyrwnu32wumDUqK+Yyo6xnXuTsA0VcadMN4a9PNCUSVZyqqbdFgps7bqDbJaJ8TG8p
T8XugbJg7ZDDOnj4yqKxNUopepd1SMd6zoxviD1aPmQOeex+mCbUBPId0z2qc+G8ZyEX0hzaHQ39
Z/uA1igKCBk40KYBmlvjq2fkgxoxrSlyEkn9Ls3hoZgmBnG7W4AOGWqcBLm67YGseaVmPrIMWr9W
ZVqDW5pABNY6ij+Sofrb3v1zEqxOY9l759e1aUjsrEqilZ5CYvbIRk2YEyQai5V7f0cMqJGoqbUY
fWo2Zj6B2djNdf0kwCBeo7Aqwmnk2sK2d2yXbCv0aZd9ZCHb/OxjyBLm/3LwjOnk4mTtPdZFIXls
jo8L2Q7ESw16CQBapMMaHX7PRfWvEM7dCP6YYmZFAPS5H/iTmnOBAHkYpnW5oJ7ttYaK2XUMSb02
1NycSKW7PwD2zVkCHn5FXrQGClJj4hz7WbGFy+XHWjWlMf4nlbiqHdwUkFxAnlTKzMf8+QRi+tG4
1L8i9kbiVYh4JGx36FukeUa26/aLzBD0wiGVwxQ1dbdWgumC8xtfhlQrriBuvSQtcysU+2yiIoy4
jmJ4mHJ2XMJ7MYwtLekmDq1jZTqxs9YYBU1VaXOCqvOv7PhaDxCehQlnhXwzh8vl6Cqbm74Rnvm8
EZFeJWiKm0sL3mrW6bT6cMnrhm/+Fh35inrRTLCDaPfcxPcF2SjFv6VvnrdvM2bnnefKxWjmx4Nk
RXuE1CkKB3RWpta8/EFcX4X2rTed4nfKgb4/9HgOV9pQz9unWUsM7vrlO5QmMwpQfj9J5g6qpUBm
a37lcxvmxjJzBCHbm1xI7Z/5PKHp/ZLx3aRsYv2V04QnAnHlR/3Rt1eKSVtEFQwtzmRQE1bLexM5
CnWTNiHTzA0xCUmx2SuTSMwVr7y9EkcZcEU884uaWz6s/IGv4054r5Afcpq00XGH2trXpXHd/pjV
zOSbl4NvSUnuK4O4Fx5o85v13utmLN36SQO3m9AF+hwlDC+cRhXVRn8XAYwpGWfKyqIsewGi5XOP
nc0zsBl7eOmEZNQJ6ZXn8CgbZNZyMjt1wojJXdsjmAF1sKhMdMlLn9ehNUh1ED95Wpc0qIjhCKKl
alvBo+9ZBKA6Ce1MPvxWAUQXQ1+JTc31mtJY0MoNwhymBlNYOTv9RNpuF4JP8Rsj3kIa7gSFegKt
mI7l/GtONGksqWb7UElvgKnfTygDj6cFo/nSQ3+xSWkD1ajsUDi8ibPMzsyXTKeS803N2fcbJCtA
siXehwVdWch5G8ZvI/mTTT1RTYiZE8kyCzvUDrZGVEeHXmYOrqwSAxQtMg5yi594M/3Pd8jMQ1I5
sqt8Gw5kwQ7YIVc2jtWcRyXv77UgMi/g+OvhC8UnrCWiKbAs82HcWLI29DlCeDJJCmUcQu91Mqcu
QxBF2cjoqF6PP5Pp+z6nYB30TbNN4mqFeSd/55yJbE+TMKthGS2ka/RQrEbDqBG+8NsXdUDspTvp
J/clwGJaTpuxOQBWy3bzb/XUhX/fprSwvyEL+RfQDGR5J1eCYFixhxYkhtO8bFmBHBNPHlX9Udl0
ObN7LU7S0rQWo3KO8C1ojhDukpI4o89C7u7PRToHtANlwCTdAmV24N8P7i8hRE+7h2ErB29igZPS
N7HlcircwfCKZmUGbyAVhCvUUH/RBTUW5xlKC4eAlx6jYmAPkKgBRWX8VLijNTYSFNczUJV0nARU
vVtQjU1ssliqOJTclFEtDRIJX/+rwyenR2Xbbr9xzB0RhH1TR4GG5NITnFVSAV+oVPtGaiG+4N8u
UdngMIKMXWVtc/ZxxCh40ZFngSkTISbsHzAkIJM+fKUpj3SgT3o0LAM6oaT+NrzEx7owzEniAzk9
jgf7DTOYsg7flrIpJHZcPLvJu/KEgmnIdyK/LojbecQSAEFeiKRRmVAde0+k/iOOJi7XxEglwa+z
ey4o4d2l9zVwplC5U8mwbS0KJKajVG7No8Sh/gV2IeGYUle4Tq0y0mhkowxIc2GR2IBA8OBCwqRO
pZlSTRlBrbneQDRYEBqJojdjvk4jZbJ/HIZMKkhCFe1WMQgv/ZQHVzXFyHDYnbjFOUMmqlP1/7Es
Cjg6r+4yUvbIB1qNaCoJQDVXym/0Fmz1wiL6SMjoOSxWf1rAde/CkkAiKBukuUFo+sAidCJB/+N6
748b4bWNtbbX+7MLnVDmNH9RhWwAYPc4hU6UsRlmR5qmsAH9GZbcRSN4vwmY/fJa/14N/hbemW6k
Ia7YvQ2xB11BGZaBBNq0yrd08sgmaRfwBMPju6ETRnT3XSZvHEPLg3mmlQM/J8LUX9oyqzvNcdQe
7rDkT2re7AIXJMsnsoAD7W1DzvhiLwFBUWtaiMl++0xAmL79e/1/FPMIXsuQDGAzIVXApksE3K/o
+jkrCtUBTvy3dD2q0A02PX572YIC4PGkXjy/BY342Z9uDK7iEjn1RvefPwyUpmIlS4L0+4V95BIz
HwFmaNT/NPm9SNpEWQUfSKBU4n5SVfHIoeHKMyOzyKGGcgpIZEMCdgzkEqll2yS6gT7lj+oKzayF
upsKgSsr8m+u3nhtd1cZKmc/LATKpJfLDA8T6Cis5b9hap8mdaHHFf4qZ90WrG79Yhd6qM6kOAmF
nJqSpb12JnofefwH3nOAFoPdHe0YRMot4+NKiVXTh8NOeRMrr8/2gMETAdhi2468EdPrh0JQ/o95
pARoCbLARExvLfQsg5fFfshwpvUoI3ahP4o8HO0/K4qGSP+ojozdn/XLa6ChS6fIvLmyMkwuCQRR
y35K0zr6j67G9XIth9kASstKewFMTzMlIppchiuapzPjzHyXgo9leVh530koSYN4Vn5T1/c91HKM
VzxpboI5gxqN3ArWPdSgfWsLlO1QqSiWCRO1SGRYTbtIJexy988kog03Ki6kuMcwV+uwa5dQgiKw
Y+LuSj2of3qnBAQLfhCBrpvKrQATKKKpraRc2t81+kdv2O/pj+tpOeS5ZwkBHJsBNbexkfDxrz5u
Pilj4AkdXMSvR2kTZ28Ba8LOGHsJeocQFCIZjlDQBfklJykdDb0whkPPUJV8pmQMrncJWcyPulE9
S6r9YobIvdH7DspV91PVkmhsIx85W2qYkgJ9avXer5HaYPtFYCvDDUVhdgLeP8A1P3B8+MI8HO2N
ri/ZLW4XIkfO9VvLtEaY8PuEkMZSN8p1V3An1BjpVlc/zsmSoyGiRaJH3FTpcCAg+MA8gm0J9BwB
M2BzLfIxu2tSx7ogwZITfevxOXZjZ2GRA99FYwM/hQQ5mtrf5SArPfI8w0v1yiyqfoWtJNss+YyW
FxrY1D6OQmeMM8yMZm0ciZXJf9SQuFir22wNQ5e8DJsw5AQtcum4E/1ekHiQ161kopdiFMMejCTl
mlG/GlTk4xWQg7o1wHUvs85jotRsFJ01nsbaHXaDc83wYp3H+LmIUzfPIjNyBXeF8zfo4PtGSMAo
fyyZIxCuZgIi9D/SLVRtBphnK95BBeXy86tuovBZ/2GlL94vz/8HHe3T8WlnrGd6VjibPoDjyNXD
c91f3U+umlh1Y5UjBAesOlq2T9SgNeqajTHKEfYFnz7aZdqVVSCaQzn1ojHXrIldNfVAO93trbNi
HFsNJj5s8wAcPAeJnhw+LqE5tlm+cIF1TCWfyVl7waRN5aNNlkMsxgxC89GLKJs3RZgJu2dqVkob
ijaiPrgHjHXvJ7RpdGy4CMXL1p8EQkzP97tUv9BDS3j0SF07DeD3pgRSk4XDUM76OHNVcTqL9AY0
3Iyf47p1iQNvjUdC2PsILsEFMOlgr/eYCCQx2scjf3c1b7daXhNmwSu12WKmE3uZbkangG7oeqCM
+0W8E0mB6n7Jkh15qhvD9FqSaQCplF1paMuLcXZ2/26sNFy5vf0DPQcXLF8t6D4n1+KuS4A9HHKm
7vI4rg0KKYNBuzG8P4cE6U44y9lD5eYDJjag0YAxI95xZA8W2jIMl+sixZBxLBeKtTkWshjLQWr0
7FTWOfKel4QqjcpArvUKV/UEp0Vi4dIWI0LldZ4Xv3AfhK+0TR2jIeWoIU3K70geNLyc7FNObVpy
1HTnX+gitstRWiqkHWC02n+VOZ9CTBBRyJauZjhdFGD4EUsIO9ccBcyLpms49js7Gq2HIw9JG8/z
2rmzn+kDU9khPUQL2ItHkXiDsBW6WkOdZU4QIEKnxK1oiKuUpbBq9QnyAYcI6e6meeskqapMJGUV
ADLDFlDEYwzQS82RxQYBNXSTs1QKn01yxQC+IEfpYNaI6jejAEriQdl1BE91IT64IA3MS9p6fyPq
cOKLVlR49M3N+dDZ/BVBCiSkbClWpqNt1lnrh35IpeCrogVolPV/h8e/3HutYwgCoO7HpgL3rfdG
Bd+rUfBW0tSRUr8SR6IFX5U0LWchrItCclUsGmntviDLYK0HwxvfA5TjIPfXBZy3imw4AVf+OGeU
sN9eQ0TTriuJxQ03RNdMlIWO+2oiq4DibmToJJQKLAHaG0MRFcao1OkhHm/eC84OTBouFvQaR79y
4cxXEz+l6lfMYhABGXNUCmbLKlbjYEFbpXWwGyiXblv2MaD6aNNtcj9WVzRLtBjKju4VbIQz65Kz
bpeKyRDIPVxO+r2Co+BCWgen3s4tzcFOIx+OTMPOrpoL+atiZyrPmIkILD6cKS6K+Mon9DpHxcFb
VzFvVG+8Inho+xl3vOwNeI3mQ+aAEgZBXh72zRzRalu2FPd08/cjCVxI1nZ/6Z4dds3zDj6Zy3jZ
UK3MKgIIvER0+saPi8un6ocBy/TYWypQ+khcwKda0FOKGkSfvSfRA+8+kqG23AzUn83TP4tVAg4S
PEsYkQnOW9CzwQbGk7eWENfKDobiPykHSERfrOSQdL0647GqhdtkHStWJTMMI+niHz6qYuNYJC+2
rIfVJJDp+Crow6mAGjgwnTDoeetl3KigCqqNAn2Cfx/zHrWE83eyjYHVWVD5W9ynPKMGqsP+jG3o
OBgHI1TDxlD1icKn1Gt4wGdbL6nCkEmDYGr+RNKvFb2ixJvJepON59cZO+KzmMgybHVf735AFkz4
TT9emSLi1Eg0JamJKzn8vxgz1+Y+GP0YlHX4MbAOwZNpoyWlUrMSf8VytHWOSt1sEGS6rlKPgPvP
15pEd06gLJF0IPHBGj3YQcsm9oGSaHAyVNSCaGLh8obZH8BNILWTjanN1BEcpqnGT+rsGJ+dwMIt
SmXbxkYYDN5dEgwwMLBFDrXLTFch7ptXWzPgQ93HNhiiIvycPoDHzHbDYODGG8KMrR2t2Lb9ZD34
DXkI7FNgprn2cFNfSCspOgjHKco6eRyoQNG8UQ0HNrUr239HtWfxVRKowHk44+cAp18A+4qYLUbc
mZGH2QzNPOd2zpVQmn86cvCuGyM16+RKa4WUEpADqcHYsakjzYbJbocjfkJ/iqGpRCgRp+yl3PRu
cholzF/P2FE7LltljGs7NxDcw6S/HvcN5nR4m4l4jOMJ2SQBXJqSETK624YbPb2WTyRPPMnffiEr
rbStYR5GmTcu+hm+UIuOX8Z6p72aO3Sypklfcj7wEFzjFyOa13wrdOTgfahfoLRzebs/lQjIjToV
XiRlNp50WCYwuNOIHZKL3Us14TEVL8XBYSeLkqiWctRTvWRvzkLZW/q3x521zAuI3QuagMeI2uK5
jZhmXWeYNndyfUxjeQNWuZ12v+Aqe0+zMVj/jBQ6EON8XS/YYyXzLEAKEsCdgfd2Uc2XxQAxuivA
ntWqG2As9Qb1lV9OjjQNOkJ8cPgcgu5s6gbbcyC6aY+MshI/2VvBnslX5zg7rEBY9kPEDO6epxxN
Tq8fDnboqK9BzkdnEIPln6670MgNVH4nk5HssIukUo88FZt2/wx+x9bloH3HMnv4bnwDXK1vqwsv
cikcPg6jzjiFzqWiPSxCAWsABRRPM9AQYR42ZWmcjfgQKbVMVP6UC78vgbow767Z/Dr9aWRYL3xv
w7VctNRg7LUVTe3lZTEzU4l123Z/tbVItV8u8W30Uk3Y5TXgLR77vxAKEVdZTYKEZ9jjF9Qx5Jpq
rWMkMaovGPpTe7BfCZTu1gOt1VpsiCWF/wot3Z2M3tfDEwKvHYEVyL/74FDEoS3z5eTB2C4hvxco
OPEMXJyfAudYZoSHRMMm0ytmvPBm00zjZoZsxMq14spmKf8lAJUiSJ1exRj4ES149XE63mW6lCXJ
KjQ0axx3tsuZiMC0MPL32kpEJCB+07Eer6WTVG4tdAkxXfsqtiBsKIAe8BrWLnMPHwEun7gwW5jc
AxcEWSndfWQbP5Ts4j8lqxPcwOjBoGi0ZyjlNS5M5Pjz4LqoMZ7xG3F6EwunRzeTwlnrnmKNwmHD
K9EWAsr9ev6qE+EocPhCjcJbc1G8AOyCwsogCWbJiP77r+gVN8VnJWihE6H97CX0Nl6vrEj3/GhT
uv60Dg4V18ppSZbFQiN2YiUe5PDPW66Wg0XZ7nQn4rlXoLvda52mWAMESNPDI8Qbp2MTWrXaWdNR
PLBUkB3k1z1Gnp6KvLWUTchLzzY9D0AGcz99ZTpWyBZyIMHnOPXoXFzQ9vy1r2Ha1YapB5+OsvHV
9L9wHQssatBJorgSo3mvbY5CLUx7LtkTDte38tLHKZsmpg7VSGNh9LtNpEwNqe9WKNogDLDhApRt
rlfSz3TfUTQFxsqgIxIqrMI64tIQ1r5KxZRFlAtDOEdeapvHBjhtoclo5FluhfwuJnaQ6UW16+xh
DFP048ygqt7KxBN2UEFfMRu7xp7z2e5hanpQMw/Mzx2uUlnmEeRJ8DVba2mVPcJV7Jg5k9r+rZpC
8vCRt0R3lNnGihwQgC32USHzFksuoq3td6uUVKnFtTVjJnrJeLGjm8DQYX6uxbCa1cL6ZGcCE4Yg
BDo/jeIjcYQTuULnq6zaMq0JjkFIQ7303I8PP37gEfRzHuavTLbgbZJSFw/HJs880ewFFn81uM0e
RQAjFTpjgrqOtD32dfD8qIgkJbKKfmYEmsUZN3a/0VS0WwofCboOT3v1ZX9WvME2qGA5nRioyjiA
VbJqdIY6VfsLGZKm+t51h3VvBlRoyvR+UMWimPYbLZR5KW4TzpEwIu7Tgtw0+X/b8h8v49ufUIEA
QA4t0fR2mqhkAUMDJ7jy8ffqobS/bAWsPzJgim11/HbpIiCrPVg18ceDNmjeeaXZfG4WpLoclSoE
lbvRfNZkdOD3WXmBpErA7imaEUAjHz0Mgvrq/E6YTN6Evs/ft+KFFMADomT6Q18xH0sfBv1XGKKo
UtF4EIrFpSn8aaVoMgHkGKYSIoQoF27+Au10KdKLDkK5NusS5SQO2oxloYAvbaCucQY041dnhSpM
t2b4QuapdzZz28++jJMnpBmDPeC+WCK1EdpAqzpOC9jLMQ106D4Kb1l1tncf188EJs2QOK9URLRg
woJ0AOPM/0xqS869A/sXLE3GBNign4zTu17YGWCrfb3iVSsSTD1WPJKo0mzmbVKe7Se1CjbSKCOE
Nnv1isdytiNI9S/v1HZzr7Vmpr7d7SLl2cSIfY5c3yGR7S6bddOKhLYcRVksL5z4daXXKx4SnjqJ
61zAO8adeY3tcPDM4U9/3yhzM95c6Jn5WzCh9LV94ZjAN4YrHwhoRXqiUzecEpo4KyXd9SJtMjgn
xlnQwP4o8Kt7YXfN92Elv7vEoAM07hQsnRU3Io2kGAfFEzKMIv7qlq/wMhxEkgWbWVZVv+3PxTX1
LYfpK5O2fwgv17xUO5L8fMbXe2iUhcCTAN/kxUxiUH4vZ53g6m91edpmWDabrUeQ1YI2ADzt0moC
zbdgrHl9m6MMUs2KBdQ+hk6CGURnBiCrTFjOx2RSBurhd2GE0Rx2EEOzLZcGOWy33g/P7c+tqnH5
Yj1GwlhsCvPMPi4eGfsG4NYTA71N2jZkep6DLB+AfIf4rjPpiAx1m0LJyNJ0vlEwCTzjY5L2rOst
Ei2S3uApkt59hKL8w5dYZ6IVb7otUAbl23qx+2AXQ6Sri0NjKf8eSE4ExIBHGPRX4/pSqhT4/325
LTNiwwz/Y34IFZPWAZAj40piBXfiBCoXPkiv4X4wkKmSt86yGBTC2r+yWEbahcBUJP3v1CNbVBMt
Il8E+A0CeTDoKf1qPYTj6W9T9WTS/SwO/NGfoFhqIWa/sLWd5rHbKaN3LShSHh/5abdR7H2xAFro
D7yLEsPYhPIgkbft7xs/mUnPSiwWoNlb/pV6wNEFuM6bvGexMfX+PHtTg/hpn7ue85OgebNiQY+A
ZMA5QhvTWFjF59lCKa6p1g0kaiyFhh0e7QknpJPDVBfdU2X1NWsJjVdEB0eN+iT3DRDtcUOCpikH
eXIkkxZB7QYXPYvpJ/7eVRiCi4zRshMyafZuUoj2cz5Ok3RAx/qaPWJPA475/3yCtUj3dg78X60v
rDnzbBeKF7+gCi3gDsmbq4g8WGIh+YM8cWfPtSgU4MdjJsriMe4bsxVLMt7G60ThWZb/Ra6/l+AH
O6DH/EkLs+SdR0FYiPxUbYoIMSxHfASFyJs/TqA4D7RpH0SRshb9Qpua+tuIefTNkmJ/dhS95pxb
VuzOH8z5Ft/61QqDZVLHog4Zx64V/9JpThylaSYB8gvYGjOXJBtBxq1wgmN2saai1i9usttOS7j9
L2/FHgC+r+ibQA/pRUNabP3c1h8rQvHvRUH+nVuZxTGEV1nroqHt/0cHHOAvHRe+iAqDuUSj+YQO
nL9cPpCdAw5gTpyZaF4D7sh0U/3dil6O0cRGl18CMz9YE2bn9i3+bt+nJlpq4RKsC3tVzp3jB0qw
MnM9UaKnVl51k2fedwTN/G0d0ON8M+JK7cHFGEW/FsHto98+yW+8hYk6PA3yf5fGEFdUDHDRUPJa
8dJeNNY8z59lm4NBX2dcbHkgVE6xmIKjWwDOIcBCMSsMlYMbExvPb6KoRzxhvaD1Vdt03IhNSmZu
ifUNQyTtQIY/48na9EPcmjPROVw7YMICZKV390HYDXajkuJR5Rh2z4+CVoY2s77bbOfaAsZl5TsO
wevlrtEw3jdd/AwNGcWQLEY6Y02A1RidRfnBWUW1nQvbSX1cJ0kN9i3g1m9ut94zJRD0Xi0ey3/k
W6EpdZMMxqXciScRiA6Q9JGYIx/B8QIkmB+n5KlP4CEtbH/+aD9jFTex6SgZlbDZ5BCmLFA9yqWE
zFyc2d3teYO5+YVbWxWQzj5YDc+C1pnsUHVhA3L9VR+Eqad4WAEG3/h1xP874NNNuGMYQJoVOv0/
GOR6paFpamZA/Bw5PyH+pynga6zLJ8ABMG3x+4dyxm8AKq8vkQr0hiIvtkM0mnclk6WqZRanHAlu
e+MsKW64R+f05HzD4Fg3I5FMrAupNfxhPH3FeMri0tmFGschmh7WsfmpNYpHjEnWkj3ilQs6KE3O
/u1dfLnb9N8qA0oQs9g5tG76Sag4OBDVH7Lqyl4wu1CKxHUFSKMaksAVoO0c43yDS0VapJSotfIO
bb9DpHJVp8/+6K1FN1oi7w1Jw+T7Tng616XX6zQbTiEzhG7c46/SZVjsRTn794RxzAg87xMQz+2V
pT+8fQqqoFfITC5lbxyyxFHffeWyful+NGFdegRlnoYEW8QJAaQ0YftVaWbYbn6DWItmovSeuOqz
CAMAqbzZzZ9ucIXayT0trkylxGFRfAn9I8Ll01PNdfgIMQmr4lqKVW2+368E8yZfuAlbVHwjwa/x
68i+5qKvhxvrwmNIuRMTtQkM6LgRwq6pl167d+xqCBBBTwOfRoaddxUr6gXnnI/9b6AhefnpvFi/
cQFLUQghtDpZmWMi3nkbEoUdnVgcz+TdEM+iLC3YUv3iWqEISnAlRmnAVleZByK7ZIi3VfzM1ZLP
1WRI191eDgFqrRmzdcfz3pruZdVwrujBgwsP/f0Gt9WmMDeBsJe020DRWzW6koXhDIEpq7JR4w8j
aC7U+5/JjxLBYzGTOvK1ZzUbVnfCgC578Cop2ts1g8aav2B7qs9+z5mYHQTr0SsmzNDgxvqDTuCN
gtnEW5s+n+CUIqPaVdBnIWBToHGbSfBzGjBuXvGiaNjLNvU6D1j3YiYyi/+XEtWQd+fzkA3bdePF
t07ss+yr/s4H78cREYKDn7NLR4HrYNNxZCxOT2/AyP4geCRvivSmFPyqp6EL70GLD7vWWzFI/OXY
aKrPhwVZJzeFIds9dZci8dGqmwCBoXhGUHxLwKQaZvOPo8+ADZEAmnJQrleMPwVsgG+PRxN+Z+m4
D0eb9XLI9vB/Yf9Z4gNK6/IdXDcxfltF/NghlfVJZ8VHara1pbW4WsKYbF9y+Xa1dbirlmqpq5pl
SJUrqJva/67UCeRg85dNnbIFnFfJK0chYrtnOz0c3CrKoVnJ4jxZkbUFMRqIqMUuOne2D2m91Tbk
uo8jnYj+rH55d+Y2SQmH3we1YBQW2IEy3KbD0PVnLDaTjPDglnJ3HGWjxpkRjEwqOLpDxB9gJ0HM
MxpD9lat6nDvjRl/wRMaMuZUjBs1EEJrFkH5Y1Zdk2RYtMLi6zxffCceJkje65B0+mT9qMTbmvn0
FxU+S74m8SuD0E8rRCqw3cDjPHi2/NbxlI4tkU9lGPLT1ROTEhnS4qnUkuGPzXzliEVleJiV1EAV
tS0upxqfDmgCtJx6ihe1mn1atFGLWuzUBmq8ZL2aj5Gd/6F2v9lm7Dkxa4BfAxUiwCas+Gy5OTDg
8P9Q2Q9YIf7Bz7LjfXOxaJrJdKgGDb0nHIWPD93HXemLUkjtViGqf2WrMITXe+EV0byjyAbVTSNT
XQpUnhBZeji4drpNS/+4ZOKVPYuIZz2dsiPowjoMBVpWbtbwEjlbUV09uA28GsLakXRuZFA/bJpD
rCLbrOI6aHF9ja8k/yiRgVwDodGN9LoyFavQQ44Lh8fLzTRWhrAc693TPlMcr75uYwkxh2AcVGaY
+JlGavQOL/osYa7mOMLmoiPb+66f5N/29ZsESloSStKZ3ndab2OCP4sWMjzqWRH4WGtj4/DrgKgy
x0yQlhsalZ00mWpsiiXKgV8QDaQKOMCK3Q8UNx4W3ggspYoYwmCxkUADQvNbMI1EwKMbxHgkcOsr
y8baYMAED/U65NVoPMTmLgPGQbAdYYhj6C/TyvSe1Z9oa6Gbl9/CQIg0J9BlC91SqA/akk2O9wia
ZnAYOIq2aduLaJ37D0qOUdR5yXEBGxCgQQlxwAfXqRhY4LQTHC9XCrO/xZmsf2fyClQb+gM3/WTn
72ihePRpcurt/rZx2vDF+npdOT/5hxZoSYrL0EmCJvBTEvKL48yaFjGjYpJ+8dSbdgE7nLr/NgCP
/fkpI1nhNPKiKPUWPHaMlCxAPIC4/ZA5Lc2wzDne41lXHY/HZqOAHlhy5oMsB19gRZc5Ad9Btrpe
BmI0SeEPGgeSjHKzX16wnvgvRrzQfhXeGUC+81r4M2LiMdPKyG7/ORxwylRHR8m4YH71WlPJ69v1
UQfWq4M6r4FOPcUjXPIZsIxC6pcBpofA/WzKhh9D1O3qEsXwtZylT3r6Ln1GeEKEZCmsc1MicIyx
nJHJY5h1Dk5G26s8MhdsM9VxAetiFA2WhAEUixbanlzIH7QG3z+1QDAhC6HbUeo7vZ0YwgQcxk0m
8XAc+EwyNyUjPhDcqfYnx94IWs95lLUKDEid5L6UKIxI50dwVy1CVv6nu2XUpfYfZAd3pDMoRmEs
WUNs1vK8VsFp6y9dMYGK8lu3VT3V3eaOAhcSoMbps196bTCYxiILTdbE4Wz8DLFF1/vUiOgcvDGn
ohKDeLYR8aqNMU1BHWTbEyVKiWv1t+R6OE8bSqqmADBlRaN2M2RoQrEERnIMFB2Wj1hQ0u13hLJq
2DGh0XnA9LX0lHLVlra2fM3hxzN3F38mpuF5LSWtiY0XbUU7VO/Wbli4efUK2q2BvXVIsnjd7hPN
/6cMrRxWpXSQ5tdJbIHr15C2rGO/Jy7w37heS1AYzOCw2FCuZ+oUfv7AJ5+4FrD6tsTMllGCLZwa
/jY0oY9eda0xNtQ+U8k9UGk+yH+rBFD7a86VMD8rRfeEWNRFTcVhBcPRbCeM+NywvU8ShYWCwudP
5uOceF2YEWTYts6gJ2XPpC8UKqVVFsLMOHiY6U4Pq2kIjyIuBELmgd4D+ojVv4yNyuc0I25YWAmn
EDZ3PKUwn7ricI1SKiAMWkf+mCvZB0ikh36dl9T0Lu20/ZW5GsocIf/REzwkth5kWJ8g3tz5jydD
dkfMhNLCdJn2LlWlM4WMwc1rk99qHcumZYEdS1KfYBNVhwhct5ulokd7rHqJG5gY+OvsBWOQH7Zq
YBTvfxKRXLhkIU7uXWYOIr4YPoaWpPtVe4F7diuu2DCwz2DQAUbdXlMHCBy+gVKnUhasPp/GMq1c
Xiwgr8tIdESisB25t6/g+gCMChOw2tRAwjRuy4FRzyMrvmHLGcaJ7hdNU+U4jzqqAeP/FLfjIzvn
J99F5v20L1ZJU7iiaI2+9VFcPn/3ZV+ZO8P+xftZTw1pOyMv540zLeKE5S2XgDEHpOIfElL5G04U
lXuOTARuzmqYMwmXJere6yN5jswQHIAzeJXL/wY8XiyFXlQmiaUsD9r9lWQS2aTgSstWB969BDgv
MWguj6059R/OYkY0N/exmuApdWvgrXMjmXHIduEgXkWkwp8iCIjoc6+gxdmD56lGUxhK4JuChteZ
Q8+gi3sG3tOXp1Dz79N+gesXUvoWXLjE7hcUgYENZLIbMjSeukpSzmShNvpnCqJvgTUXQN7ymj32
j+FREpgMh7+zZJNcRa4woZNYKn970I/2GmuLMVb5mYXoV0awQUVY4fyn/NMkAxVqBtorJMc7/Eb7
g/tNccW8bBQCGRBV5D344jcj7BNRQIeUCjeIn3fVsLmuUIZinPIPlADJIsCM9uMFH2Og8PGMsFjV
eFnLelE6FD2+CMcYshq7hs+6m69kkmtO7Fb5CBa5zs3K3mE3oOgbUdkCCmULohYAm/MpYo9g0794
9bRnulArx4mNCw288gfsqqoxD+fizIOhPtd4OgA2oXA0hJa5JEAGCCEGB1smjohiNJfco76mMqQR
GsP6btudCShU3y5r+QMmV9f1S1pzgnJQiTozwn78f5SsSM3eKznBHtg1CjqlIafJl1YsqHK+dr3o
u3q+mPbxiOnviU4ZObmntikr+ZXessLqE7osSFLI+BhR+NThCawl5GI+5oP6kDPEO24UlBGhr+c8
crXPhvSCbq9h+RsZnrt0UguPnSLO8ncrIMbwYQWS5pcjYjECruPE0ZDw0SGsJ14WlVeXrWWHuRUw
cmgNpokm013Jh+2ZsYqZfyiPWm5Xol10BuVSc4CEwH8GLeQaYk0w8JbltDSycTKacjYQ4qMrsU4z
zTeKOVrSalOzrPfyDzvW6sMX7eBzeB2x9zUC10QiXM/gfKTfpdor2IlK5P5OqegSsfIBcUOfkfle
j/Xg15M1PSjz/Ej7i3GtcsbzMwT9/5/nhjnVuqY1fuIKCFQSGtvPM3+Wuz3LDfzd5kNHsOxo/gqH
9xyluXbYGyrM8wPTpskEGEHXAyVTA73mnMHlqYkd9Nd7iwu8cErrqLDz0xXlhsl9Zfc9u5ph0950
Ei3+ABVP+TZRaaZ9YShA1I8PbqA3DFrWd8z6kmVoKWWiIf3BM3TgzPIK+050g9vHICflJvPJ4tOK
5NtIDu0JnSSPniQCyskJuKog+bPWq1LZu2XPX/EQptdB7NJ1TVVUaxHD4/FmICAgXUuHCnbyJoZQ
rBYzQZ47Ug5wqtsiXEyUnxV5pjio2lFzuZVF6nVZwBlIuqXff6KAap3yF6aSm4SummXHuFo+FF6P
prJPIDEcRGdnjck9MlwC8RX4o5BhF7+L7Fh0eFUZCBuprHnZ2YDC1PTpGJKtwGKJP1tOLNGWpKyZ
pCE2jwmbqg5JnCjp/Mq+sAJ55qAp/sVE2zZz+n8Z9ufxI5UOQFdObyNngSF0mChlX3VdGkt5Rcvh
mHWOso2tDPvlboLR7BqexHtuRLIjTws4yXVAdSan+rrBWnPQxD9fgPZOBqcn9Uxd9uXRhT7B40zr
TWQQDEc7XoK/nEUe7y/TwqKg9mUJybdul4DERCeCmfpZBvZpQw3UQob8oQn0dzJ5h1TG0KuMpbWw
mhRiXcCFWVphuArIWhAJvE8xlflQI/cLDiBAFOyMJaGMKSdbyvoitL/W+zdFMQb65AZxJd1JFTDQ
jN3XuHMtOCQEwY27ht/j3JfZ/02CenPToZpC9uFf5aqmhz7y3SRl8b4/jPGWl6qOBVYIpI53bBd6
Hcr9I/u3tNlpcBJvcyfjxXKP5mCFte1AsfKkdC8Gw4NqkJmzhr0q8T8QF6zI4FiC7HZvSmvztvUX
I/eidRN7pMVo03qoqYOjB9hJHz6oGJRa3+SMeSCacEX3EiQIIYVokVFX/ksaxsdmKKqQ2h9YNPog
MmWi5hkyKE/DOMP2BhhPmmWGPiaBXXWFhoGeGuqPB6WfJ1iOeqHt+20ZkQnwoTM7tFmoeJ7AY9o1
d4e7xajuZCAhPUAejoxGvCnDQjAG0JBKt3QMl94y1w67nff67fJgLid0om47XXCbADkSFz1yDl0Y
CfYbZJ3W+98WdtMaK0mpuYprKInc3s/JrFhw1cy0hv8yJ6vZ36NsFITWlcnm1dNt/F12ShIxmhlI
eQSF2jTKxRAH9sv1SyAeGQi+gV4TcoJIsEF6LlcHp7G03+GdgFKpfHMz37ysQuXWaMVE+hO/mEbM
ABFXGbR3FRO9FpFKiKjPxzT/1ILm+WlurXYnhfnyiYn1pkA07CNgW9AbPGX4ZdZb+TEB+TJzcn+o
TxnR6fIJRapMfGMQnJ1lyT3QJA9OH1CTIzLF8qufRVXbg8lPoe3brNxUPeJh6B0CJWtgEB5zSXFW
s7ZTBtvjQ9U9ai1+RwfY2OKvhKoQPH3rpS2ynSY5q01RkCZzSV6ZM63biPynLOgM9nbbBahctVKM
gailfsXDde9Qt0Vpb5oxyEwwmwvT8uayQORns0ArH7SUbijJ8KdvhlEy9EITMVCScQ1I5XMtN2tx
cFBjj7ImIQQKn9zJHAMXbgwBLersNMqn436Gekd6PRtA/GBN5lpqtC5XHBenbngDtZUFBiSib2Ie
x2Prmjgh5ed7wVB8QJ6+wcI13rA2ufGF2LsUCFwcr/o6nRa/+/PKlks2u7r65RvmNWLXhR4txbJ5
x4rYJmffXALd6lGT/W7rOQTfTkOmVFV96QieVwUiQ77iqizzGRTxFIGQu9JtHi3f3IO4TKISXMfz
CSLqBUN94ohabJiHvCWgMAA3YFWHN/TjMre7DIeLyJo3khOfdYOrX8HA5XLjee3eqiV/IuF4Z38W
0puHwjwk87938LA0CAJHttCu7ELaOFqqheRb2djK09olNaO0mLC75a+4YoOMjHBth8EI/IQOtoLC
BYSjutE9egJjPjmKBdjN2ifaqiHucle9dTjd0sDAYLbNcf6E9N+XpZmi/9JC4ZVOX1GPQ1Dmd+Nw
eRmh2qk0ns5npZTm0L4DabQwdsSUhmCXxzPnth9xDLYJJyEwRS4IdUVfPx08BhYVCEM6FGlYxlHn
+ShWUUs1yLp8evdxTCly33+uiAaQ4pJwMSzHq3ZUoYQAYXnpzoE4Slxz5rpaz6ZNrIx0BDF6fcZB
t/DOaoSP37Kg1fy2gIdmOw37oI5NEc9othzI6zHq/ZfBPCMaOVmGN2aLP6Zj2GMWMJmvrIxw22fI
0vTQVMErCdsN8tn/SuI/X7+DKjOVyl6naNVVn3dGeYXvx4aYhmXciHpouEGPVQXqOKtjG/J5PLK6
qO4tf1qCwB36VVUOfQgZ4jQUwjOC7EQlHFMwoqehmPfjZbMRmLnZQTomhsEXI34z7mV+N0Ll4EgK
MgQXAMtfw8PsJtk0YfL9M6itagZ+4sz61EieHyHRlhcJdlAWw8wZ4mTlEChJJGYZ6FG9d23xF5pk
qR3Fv8rzTvejjEaPFfq/xnEdFzwtWv4gmBHaOhgL29+ydg/VZySDYhwmcHN0YKw+eg37EOyX9Lb3
RGtFGN0n+tLVbUvTqFqMrSl6B2uVvjNVKdqp5T5CzKiVVM9oR/Mn/4EIt7sy7kjRDT3OHI2T09Au
vzFJnRFJ8YOOFWU4cczyLQiBg9N113PDb6P++L193ePsynjT2KwqmfH99kMWvlC3/uu6YoCKy2Fl
KZ+99oLU370OmkwqJV8HdQQ5GzxEEeqTmN2v66ZlpTaxBjhLByLczda49t7gBajMTZjEpP86J6fO
nDG0imyp539hGJNrTEBNf6oW1dcSqHxZXmeJORew4GGiKBW3mn3woylAhX6ZiNUWfuSpWiVI62v8
zOStKOfjKw1bHCYBpAt9QZ73j8Wu3u3H/AXfmNPLYPMtdRnNLR8VETPZ1bpp58/gZeeYQMyJKEZs
lm1Db06uXcqC0H0w9Xdt+Xo9crZaPw3FfMGw411JsGBB5Dr3iIXCTVSdRm+Iw8pzRowNs4OvimE9
20SsjQGPiDoqudgtm7k1r8BwzCky5axeQJ6an5FuuxEWZS41puTx6dwRwtepMSXsoB3k0S7q+HNj
+GJXs/23WWUCTwjyKONtHRP9iDv+f6nkCg3A0BB2qNaklsCjzjrTWB0gLY58nEj5kI/VDBO7C4QH
FS1Xcx6uht6kjdrQz1WtU4Ti/p+ZmBTAKvB8Cul7ZynFma+X1UYVBSYJZOgljxP1rAjcwdTTFTgG
2Adm6FPU28xOY9V3pR3vj/9tu+4fj1dFgdGFucL5cJLn5R9nW+60qL6n/lfeSrw9eBChRXwU9Ffh
Yf4FmOwzxL/wv+QooZgzaq20ZHrLCQuZdEuq61E1I19L62kX20ccM7/JK38I45SPya/BgWN8cQfx
v6BopNyP0RIiiTzY6zrQ4i7lXWORFdPXT5mWi4Vc6o+WUSsnWiMqXk9FGqDBBFT9mcb0cDeIpND4
ytR9GGkMBGhXENeGEawpT91srRDU6SGOpUYQILv3ehxfBfMicIiA+6QqNsT1I8pTOZdKz3vHEzVS
UMxA2npRy1NepdlsV3kNilPLFqzi+3B/VBfhDuk5TivGeU4ORjoEksCbN8rkjQIYJ1/TmVEIwNOm
2Zr+2Ke8oK/q+OQtO4FuUk0FUc47HAUbxjJTEsZFHUXHI3pmmM6c6ar7h12kmGvE4XMUhEqT9bFi
XrpdQR8vVJdba4k+DQzb48ODSaPzj97gLbT/eDCp2m5MEQuTIsI/RLy4JGQM5b0ZDlbue55iQZ8Y
rmqjKAavDdXdUIcFMuxUI4P27WGo+mwoo9pDCwcV0FIu9goJ4Iuk0G+ZQOuUaZKvg1t6elLmsLBa
xbswJoqeQfU0xd14k6zOfvUtOtyVZvRXfOQdoGVx7GbB9S9xG3vauqMgiYncEnVrOAIphBJeSpWD
oUQ06GfLud88GGCEQ/Um0zNoCpwt0SgWkdCb3Ei3UqYxjFc6fVlwQ0McDWl2sHCaxu1SfwTEac5m
16gssxlb9hihLnKc7y2YNvkGlrcRHVcR3Zv7MeYsAFOYkyjYhqPyWE/+eoIVEJ3EcEf8aBLwxgV1
er1gjZkPsSJxCvCEaj9MQKa9I9O1Wv5uUtFW4BT6U83UHBgHaTV2BlRDPtffZWhipp7Kqcw9a8Lt
zIbtNtsGNm0zu7NEqQvzywicVpNyMHKHHLOi0VJO1YH8XJhTEIkHHNqwm7fupKfOb4FWhpXNbpO0
Hcy/9U3JDcaRwJJMq1dJtli9EaCeQfk9cavIUAv+54sPLAONqFAkDtX5+zE0I6akOAUWfMcKKS/j
VjnZ3mToqVICOi4gO+SPoYvpiAUkoT0mCPsM1B/ZQqVYh1ZNlscVyO3jjPk5h/8RJ780d5mLdUtM
unQy8uRsEyU3zB4mCl+lZjTZSpTuxMU8v2hbwOkw2yogz3DN+urfrXHVNdp3dFMy/poBE09g4r0J
zLbE1kG+wte0xY9R0x4CX5rEMGFmf1pBVJPoB5k0O8q4qBRGoNnUknJtcM9EQ5+baNxHSslVN+kp
WY2o0pBwMsdKmMXQFyXLkxu9g0qrhlJiY4HByLaCfABV/WjGS8HrUwzcrfMgtcwjhe797kFy1vxe
YkZzfDcvSHfxleC4xCMPesWgNyuVCc5EHfzk5khsCuCpNx2+HAf9Ir1+c6YauQv73WBdQBD19Tbw
XhpJXBEdMgdWaxJTQf3n7594c9T0Wa+/71lo23rg/vxzToZVbOjc4VMrW7eI3MUBxaU5eST0W0FN
B+/Z6XjWmdcaDRI+TTYKNHmzi/JJJDXorT105KfP9MSzJcb+14IMiprqddlCaKtp73uaZhQR1ATm
ZufiZCaJ2BzBFIgAuNzHmguskY68Efty0mo5P/7cMgpf/25bn/toj0CgUzIF8+b5XRjatzkv4bv6
1RNuCkzXeh2SMxSISWoNR9PNYKiXectGjUYGVA0teuA3zyUr935Z0C3Chau6i3XKibn2syJcM0Im
W1L24AxMvUXBPJ0qwcxBYG8/xep5GOFlBsb7FFBWOT4zNCtzkJynKHaR6gZZ3YbWqjmfxVzTl6S/
dIYf+EUNyWtRSNHxaZp0uS3k5E7SJObeaUqpK7yoLsnJflIX3WcF83Ix/FBNEYudWKFEiEspAg+1
ta56YeffWs2MIwA+X3qIZpmE1lSQd0+4zaTpbxOx1C2Ojyc2kCG/hUtriI/gw2jhR6jMcGtu7zj3
1aQtClvLw0dqfVdlnBg52WUpxVzGuSCMXlnfT+dP+ELG1x2wupOt2MC2FLWaoKUW/T3ttFVCCOW4
o+v1zK+GjCMJuYmNEBy+gVcfykJ3Ge3PNLcmVtTfOiXO2wCFv8tW3VfNpmVKkBtYXAJ+4heOBqti
UTAk0KJbIdHjG9nhmOUv+PJfHFIwF9U/W7W/SiWNZ9TSHmacZnIMDmX4MRlzYFJiPgaJUZNHS2AX
9k19LuB4vKXbQLcpjAzSSbxeMn8NHRoNoyLYfJaYlteAH52Y1ma4gx1bwvp3RSmzUQCm2mGQ6ai+
hJ6JzExeEhVUsU+Z9xLTecG+jdy23Izg1xn61Sd/v1YAtJYJFDFp9H9OSSlx/TtciP8wqAJlIKZR
QRoz3SiH7zgVIdMM6Fo1thPFV2FvYwpB5WGdVh1qlSFigoaoJZ3xTYIwXReCj+wwzMOVcsnG6l7W
ocBqUAKoXiKYN1V4LhU/+6d+R6cq2u5FE2NjYh9onoI/4oLq6P9FanLk1ibLGoalJi65PbXIs3iF
knCKu1/e47Jp1RpwvOvA27iSW7rT/Xm3nIFWCc/fmffu42SDZOUIbLJK8WESHLg7a6QSWYbTdPbA
DSHkBWH5OthbGVyHmi+QBgac8BbRyKGYJGG2gA09LrXUdpWkw51zEz2Z2JLV2XC69S0pSRwK6cWb
MsjUH/Gdx0yQfQq4SH0JLLxPah2m3BPUjzM3q2oSDWrfFZTgBLUVIdtiR/fi4MJPyVcdWPInmRhD
Fg3g3ecX5XzscAwd2qdvoceOxMOVvBZWqmPryKOlzRCQHRvXK6UhtCS1dzLDUdocOSR4r9vhh1nn
1EElfAqmon3bnB8dlSUHGQL7Jt+PdAopW1oQQBAv94IZ9Q2rPcn9UGictj7NGH2X24409E/ZLXBo
iVD6VzanHn/68SqXizPWnqZCkskxpuUeUFXkoFrm5PSm8Xh5p5/Ap0COKOKeN4BsdtdkpWCslAyM
As9ORY8SOtN5kuoZIW40OD6EfBiUKbitdpVKBJPtqf1Ep7I4ISOC1+OsrjfPBwu2q0KWpZ2LkQo9
WHhWwbPvAF5Bk6YYvAK1d9Walxp+IhcnSb6YG3GbY2syV3FBtQdG0mTVNouj91Ksb0ZIW9gXQhYy
9TOgDf5mESgi3O/K2BGvLetZEyUSg9lThRmolaSmI6zBGXdN5aVU4GnTnyK+U6chZGMEwbngblkR
aL548H7oRPd9itdGsLil5geVGPksz92rHSlOzU7VnRZFJervOOASnlBzKoBOdnFZ45n61X3S8sZ8
0w/zy49oZDgyFuj6Tt4G+yqexsXejFvTH/93gRv8UBXijpob/QyaCBTvf2YM6KWAaXnlsxLUUPnJ
2ocKRZPiKU3/pLLKRxGSBq5rbVW60QkdpZNoqbQjbaxEu3LNEQEcCa3X3gYDuPXfXA2H2fuomgwI
cIm9O+6y+/GtF1T++I1u43BXlIZKuoOXkgCQ9f3PuKJcqLC5X8qq2H0X/yKP7vDh+51xj95h82n6
b+ZovnJNfyC+J/AnhlzfugKPKbQSWeZxXEX0sUbW0qOd9V/bz+ztJs171nAL+zYVekN/t44eTvlv
6pZOGLm5Ow5TsQgQU6EvBvBYBhVvSrmIh/PdSKXmSeslwFAxwaWiQldH11Bm63mVBZHGKoN6oBGs
3MhztSNu3l5fmhUJtUvI55TdkcaaOYndwSsNSLAZkm2Y9epAmSNvE8ZuDjAoaF6Qjn3qjsPUQGVe
U8648juUa97iKIm4/kF7jXHcNvoovleImOTpQ+1ICgoD4SPkx9OL1G5XIDPtJF8BHBB8ksIVbHCc
0aSS5D6LUIT0cQqUW5abplZwseHsiDaBHHErZr83GlDttoXYYPgrIiaqOqeuZiGlmJRjv6g3dQgV
9rLY7fQZ/+qblDr0x3WDgyXelMp5kpRN5vRiGKex8ctaSwSzISyvKRD2QdaovN/+VN1nOUwTEFHA
m52mW0HtTigRndHtLfnTh/XNRudaJ1CafGPHMwiw7tUEr5dt7Ac5Z/MKDSSgH8Lxdvaul1g6HtLN
g0Xl7JMs+JfLcvC8nAeptKCVNTvLG/sa/1Xpzt0ob7177aV3z6fvirkvTGuCMe856UI1EnzJ3t6K
VAIjz1Ta9GVB4rz3PHhTIxSw5UyvXUSEkVtehVms42iozVnfu5nzNkTKHD4QwwVSFK4xe48os0Uj
Gp12N33fbfgUHkD7mY5Sf1wzU0n4MpnQhKVp3Zu/EfPaHEjYqEz5DDqG8+HMI1dxXt+0iq4SNTFS
XmkTTYpP8INCDZsuPtsxMqQjgnB/8o1pvnbu7wvhp5mvTQjJ5KjobUaUegBxhTUCV9TQXZmkTIg4
S6nMHEEpXR863L2ejXv7hjrr4G6/16crW1SkgSRLNlJC7m8/iv3/uBxAflGwN3BcIVug//4oaMPw
/ECPGM7cbJUmWcF6flKSWUrlKLMfizZ9o6lUMBGOgLFWnV2v5gxw5xVtG8BuyvZLSDNpF/MQmaEy
ShzfStke0SbGofzqEJ86U/Er3f0cTnPED/xy0cDMzg677BGdM+oMRo9xXyKeRUlfbYuX8V5yPqw7
9TRChnO6X7L7wZ2+ZLYCeiGwm2EOvbvtBX7fCnsnBMdc7mt9BgOdhzc8FIwuSvDT1C3wwaj074I3
fYadMnkwdacnzgBpQP6zbi/5CgYsp10Lgfn1TeqNQMPHaq4AbFIEo63y3pOJWGcKi1MmYUd27w1G
VD/EJ7eu5GR2wxKOmS0pGHaVYM/DhsNKMVMnQd/hn4y0AnkNeGr6Jz5kZqZt4d3mXiyGAWMrViiX
kNA/wQvAnNlL1Q4Jx4Q7jQV46h0CgDx7nK/Eh5jmzoN+MLKYZQt1RnkINg0M+9x1QNkiPk1Lym/k
YwZo4xLYyEvnaRkVXgYOV7w59n4sggW2Bgu8j5zKkkXeskMm36toACV/pZWqiCQtqrgB+GL+TeMc
Px8tN6RHALbFwhG9XdAUy/s+2cMC7W4LEK3iuNrsziiBX+foLZyg3KXWAMdzfSq9GSoOjKzMLFJK
yeXfaC7oD9JLEZmoraU8Fkb0BzqDsJqaHXKqHAQ/ptLg72qVyj7zWuJddZhLum1koRtcV3QVQ+Nd
V7k4IRJeH4ut/KkJ7eChPjvyrbbE8cEGbapJTsoLrjE+RILmIm2xQc/ljE81H4kPLlv+SN8OEdH7
ybLcTKak1V08hoSbncdTv6eGf6zHaz02yY+xVJQRaqmg3Jz0xq5swMwE+aEuRAHrebCWFSft3c67
2YYl/fe6Nt/cRIR+htGFl9bK6enTOvZq1Kazq/hFiB7CnwQ3CEDP03STn1esu89In0J9TGvwltu0
hVX2HDp5q6oGaKH94crySyPlaYqZUoYtWVo9EBJTx+EwsZtG74GS4WcUglb/8agox4NcF1AgCpE9
4uJPOKmtJ0k8HZYk1GNxOUqlR4jNP3sulg64ho6yae/8j7TSR9UbHBYnzvITow9uzwrKXQIz/7ob
Z7I1XqQkzuonrX+WfsaE1Ed0i2XjvVGgmopp4TcL+3X26/Zk9J6H0ijVoCbQ5/tVWSSAJ9in4nju
YdYsK/uo/uIW8merfmkl1ooJmB10VKIlkRJeBMCiWBs7C+UomxjZqfiEApvGf3pAvcM/as1/v3gP
FqzrC6ZElDHR/Ba9afEaYe6Zb/RGOkDDQC4BcUf3T+NcVRsEmn2/IBs3zWw+ptEVbOqGxtZwsEvF
YbyFuAuv2NxWUUgIOcij576SwWsQQ9hIKCGMxDH6dXupKCgWoVipVAU9eCHxGCCFS+moz05tE+kc
Sb3UhISVM/lCahAjoIcer6XQrUOFBr/EO6qMxNJ5rqf4DEiMrmVHcllT63y0okNsxZygzK0q93IX
XdfVd5/9KXWHHL3++7bjzze64I7nXlx2bPjQKoxF5ZqlX1gH1gbmbnZLoCauEG+Vbm2E7oanGy9A
WjwD1uC82tTiT8wPbzRW6qLNUoUADcoI856L7KQPrfUF+DWEWqTmhL/6kimrUqrwdEzmnIQvUpv9
fFpgEIFjJU7YuRVLUUW17rl8sppRjw4fHn1jihOLPHM8h7tW1UVpQ2RJ0yUWno0VYFviLiVT0lWE
Qle+mBpmI6qnwbj6cNWABju54FQEr1U9Y/f4TkwcO7kBmDvrIZccfcPhPyYXL1BY/EwWx6p8iVfr
xIx9eBQ6NzL7aIGX3mlWbOSCeCgnptMPQfhbb2MdqWV1SQc01fMcr+MB/Uqx23igBxlZaa1Sb8mD
zRnS/L2AtxqYlkUtB2VQB3L8H8+Q3lDN8ijtsbNllPqiCNNEse7xLbmVnjoNK1Y8TPlp+y+JMVX9
TbJdVFunHHJhedcRFS8t6iTwyzFMf1GSgkE4Rm/Mk+OncMC1QS/KNwX11lnOur648NFEWKcqT6XS
cYFeMD4h7PS5CN0IBxkqE4ZxddDgwsQcY7wFrim+EDPrsujroogYyKw3qzXQ/eKg5QmNcjeL10IN
BblF4rrTCgTBXpRnQ4BG9OiVJqyncMzAUHqGEsms4iZpxZtw2D6kdz4VB8oDuaphV6MamauN5mkz
v4Ltx0Tz5VcJjSKHcUJ3vb/Lkm56jI6NlJR98lHM0MqRbMnuh7vvsniSjwuayVnR2IT0ASSfe+ea
9sIpyMXMcrjtIOvs3SURK1KcPU+GULsuyyYiSuhKMkUxbn1AxROubNcm6VQ/pDrKZPA5GnfsJW7C
DgcEUvxsLm+T+DslOnK6ifmPrlLJUCD4MrWWC7a/qtKy6fbc/53TBuchZ9GSaSFlGKLZDjXJPAdi
ifJdPizaVQvqacJvkatmuFv+5XKrrQGetBUFuPnvW+FFJg+EkVbPng7V9qV3ZeNPDDcsQxgswXOr
DwqTIWxngXvWqrILF7jtsgP7N/32wYcg1sMvKGZOipPpIIQ+g8SRwdSaUJLQSrHUdehAYjqchBJp
9daciGaQxtRM0wXPBkozdP1VxKOi0igST9cMnfxVDpfkYNGn45bglqLMommm0N+DyW7TSDnYLOMN
hMKXQowT/RlaZyPc9lwKzx3b/Vl415JJ1/vloq00x9bA9BhZ0dquaGfwYAHjvcpY3FG00k7DhYJZ
5J/0FILsfQH8NfRSN8zcurUKgnBGK0oAQo0jDsKmOPosLwwvFqCKNpesHrsRgUOCGETEi6D1CfON
eQ/Fc9910VZ3AKvg0hiF1vka4S83QIGAbX3ciHkiM4cvZIreG2U+9xqKbD2MRH8xC193jzg2ZiFU
qKdlUWELox2RCOeSl/G5+74DZwxNG0sx+Qiyky5IzUEUm7+Saa4mjNY+1mbv7jvVIOVl2crGwQ4G
ljVnB3WvppKnEMTp6g5p6O5+LALsoS9iiLQdmD4sI/XfjTgz5JjNfmmN1DnTsEf4YpvphS9RMi0Y
tcQT55IpR/6AEcRHS5hsg1idb5UGhJWR6bDc4gVCKOPxhVQRWOswra4JVYkCYKDkRI1n71KgQteZ
stbBNS9+DV5Hpt8Cp7qkL+aM2B441khIcBudTIcdkSzg19g4un11yRlIS5GafaGp4QsJjd950P7N
iSGp8P27oJYmIB+BCBxHf2YSOtoWyskqQpSiqX4LAzPel6HJl1ZTzGlp3Cumv5uXtn4pkhW7y+tq
IZOWIb/UwSM/wgfnSGxzEi/Jg9JnnTlr0M5Ly3e//8EsdZZIfllS5OTfotkrtsn0iZAgV5k6bein
lFct3ylQ8qTSjdvOgqXqSWwif8Cq+SWOsQsmFa3B0sSEjOWAiXlqU1DmhvlecEsH2IpxHS02xdax
027uBAYj6n51WSt8lVk4ybWaofDptv7+nsxXU2d5pTlF+R2vTa0iSoyZ9/LrH5zHBgmD43S0q0oR
OJVM3OI+gvjZcq+MAYDJRCmlpRFq1ZzzE1EGZLUl9rSu3Xcja5SG5qeqNGCs9VOjdMDlVwMbte9n
IMXWhMvIfoEoQCdhYfAYjDCZBKu65PAeqr/6K0l5rB2dTKFukHGzeWDdfzL8WPJ4vtNwDe7pDjDV
GiJptu/KxB6BRUG/qUwfhcm8ZhAm1gW6Aw+jJ+oFYTao/eTkZC/5/lHwsX7vs3sxmyANEeT/cIm4
i9+bCWGlsyCP6HhWZy/51Q60yE4Y/JahLjAADa74/lCpqeXDeePecoJlwnsbMrSftnm7xpRz47Fc
ae9CxXX2zH37sSlRFIPLLdM8dON4Z1XyAYr65RXyjuDCKPRQeNwcq0i26Mm8t6hu5/b5UwCz1X8t
+o1X/dEJQBYTgrWUUfUZXFs8EaTOWvgAD2fRKo9M8V6OY4HxySkBYGpo2o0EYYzXXWTvdGp+K/65
piaVNSw0rsNexag7UP/k94RsD8b2muQ74gZBRhp/NNl81oWaKWxanS3VqdsuWenRrXd1bIkNA8yX
V+K8Tal50HeAhU0SjTY8RiFzlhcvG+XCpH6EbxnFUN+sZoN4bURy01UwTiOAfWnMq0gzgXBqUbm/
4m2LgLIiCdTk0Yju+A1nIrx/m7EKQHiEWF1ZMQ2qKnIugLh20johdV+tuB23SDuARSwW9Rl+ZS06
KC1dyIV8qvdDqpRdS974gCgHfloG+OXvcJLvaGM55fGageRIV5hFIcwIOKjt2AcG3C09S8Tmneon
XnwKrDdZo/A5iGVI+3RjTicaBJd47gHm1OHKYos+yAerOTjD791eLL8FT4o0TjlKQKVMxe0d3nVL
eNLv6YnWy/5VLQWzuxPVf7wr9wKbfo5z7qeW2hr+nIrFhR/aiVac3pClobAN5y5YfcvJepAYdIsZ
wPSkn2NsBHWn9SPj0Lf6ByIQSk+CC22BIFkGOMhDE0+nGvepbp0xDl9wiEy8BRWO02af4o6M2PmN
DPdeDhbHYFcjcnDsTL/i9g5Y0UsDp8Gi2hpCVK0BmCQjv7x+6IfjN5FrYdcy34npq2DK4fZ3y/5D
cRj/xfxcQeqvPM1Z0UVQ346W/+49V1cA6Dneo/qb1QLvB1Ow922nnK+/aYdafsd+SWQxRDBYDyQF
L7tdfWrnJUC0Pt67K8Sjh8JpYccozylWhrQqo0IRv8GQU4S+CpytWbyTwmwBHgWgzYrl/vEjp/wU
pbT9ytgRROsKnAo0K7R6wJfIj0KiLqs6T9DNU/XJ31F6vdcfePTEwELMVOpo7FU8+yF4K4IhywZ6
/EMT34w0V9Xpx12aiWQdJg40oP42uxixVf8nfpQ2yZy56ElxXN8VtPSRyw5mv3qr5Fnzv2ZzAnPX
c3ZYOHL3o6JFWRk9wBeGyQXoyoeVFGfRJvjV1nbaAQwv3uJ+gp26MYh+frbk/Qs3SYUdGD82o/th
7j9Pi+piSjTbNVlSKsQxKDOooouNaZsjPLeR914dpCuu5eWUb0RseH3cpcF+5Wsws70WtwiHSOz4
t/iVMmg6iw0Hf0AUZnIF3Zpcn2StFIECJH5Ft8IMl2pJGNahX1EOm3SDENOwaE8+WWVMdCIE6YWx
QCfA5dIoLucYWYA/2kqxnIcoQDTOu2+QQapamrjpsM9PAzeGD4Nv+B1gh+GhNoUzcvE0YeaZhQ9U
KDnEFvRAw9GSZQnb0u3eBwIMXgpt6YbC7MfUJJNkJXRkj16VvqtGta4sCFWn5tFxYf40l/orVTF/
/QofmLtD0lGhpDlIlUblDQ7zaY1CVgE8WQpg2lClbZxp9qgtkTYJxu1KQnd9pDfikoZOIc8NGZwn
BArT5KesuqClWkjT4aJDZkEgj769yMWKu1rBVRxn4zQwOLH0DDEqkLAxtUBdQQDrjXh27keU8PiT
pIoCouKPIRj2KV9o3aN5RM2Qcd2YL4KH/yjphEhLhZFJWBWy9D3ts1BA8YiHGxWZOlnk9XmpbhmX
cO15M6tVbU1tm6qwcnKMDG13w2IoyBMYItB9ZzLJOFMNYeGBl1leJSRRjOpJuWtN2XqGwzVbzGAD
5buw7Tc26a2hwTJgMrK4s7WGmz03RNjXth6zlGzU54PsW5c07T0pXKDnh+ENpcjOADa6KUATX2U/
Sq1SeIthDTUS7V5MUfbrhYjmox3bY/G7NQlzGs3rDAdQQcxesuRMpNEBGSJWnTJFjXhXgmlvuM9X
20y+seIpzDsCHZ1CwlXsgYHJcP+L360XJ/KFaKvhr10a7SI8ur7opfbnkMFUWlGNOErET4gYcXcf
4z7nnLLL3Rx0Evo1zNA6vJ/R0qZifdvtrECImBol1RDu87fSTb9kZ5G0YN2PmJFjiRdWgB0AHfAd
pqqQZOGtXNVKJ8//69pFkdlY45aA+Yt+ga+2Ca3fPe3oEgufTXHNPaLBC9xo9pM6WNbBk3dbS76z
DfO400y69YxfbLkhl8ukBdeJoV0HTQKrSpNNhfFNfLpAQkBs2ajXteryfI6JNuylcxYqwOxztJlx
+ZfiK4QqfJw9oTLpjA4cT60VbbRMnRX9lYr+0bJ4iUclNPJ0pi36GYojYvFKzg1d7dMtsG/wdF0T
MkMC91xkgnntmZrF9+tFhcjEnDnuor4O8b6qisXfp9gznCu//fuY6aikgV1wWBv89AzCOrJhX27z
S3EFGsqZJunVQiUHK02ppYI2Oet/eferf1/QWtrTVDEEoxJA5kVDAJ9uty34LWydG6nPkOnBjUCy
RcAT9ilEY5KBHdjAAzqrxjESgwiIJWfAL8SqyhKlsmLqNIlSQbNwXuD6UBgitpIsTXJLNhmfsPOR
KeMWYkczlcDs5kHFoa7VAkFxsOEmAZIcTade9hTztTg4xRi9XFcAxDpw7TqUN87Ozh/Y9gEOcO2d
N5T32UMD/8K321vSUIXrqJopQ+CsYuRk0xa5rHzhwY2f+wPexysg2CwDRjGJCynRbvIlH9l/7kwe
Ps4ml3X1HEHyP83EEviVMSg2OZ7IF/a/988xllXd3xE2yuu+Oko+Ic9u+IlR82RWJK4iXJtt3dUf
pqsb69MAbhJjNmCVdpX8O8uD8ADRzHPxCsQuTE+LnGDQf/5/+RrWI+8QBnn/BPBT0LYDWmbC+4d/
WMrY4FehauoPv1/4uF5hIDCtHPZItuxLcI1yikDmv+SfqAOCL2IjoxdtoHdpUGycKkPtvEFYgRi6
Hmv1FExvXtjYp2zff6q+6pjQJ1znYGhIGLm6Z+Ah7PH+ZMyPW1q2HpR34BCZ9cZ0JtGJUMmocpMo
KTTmQSRCoWRGvCTaCOBpTvRxIgPixg5Y+twhxZx0f7ZsCVJrnG+mZW5BWwfld7mgQAEuxcXf8Hul
rfwr4iqrf1qaAj5q3vxsjUt31oYspb3RCdYAwtsh2MgDPLTOfDy1t6xeTMlCYG0dV5Fm6nIGJIBY
KAPoH7Hh8UyZJHiP4qQ3DnQ1nFgM/ssHY/NGPI8avZb3MEhAwDJz6zO6fkYkSIMZH8rg9jaao8as
pbQ8beRK3WTnBQVxvYiQCp1ey82SQ5GS1JG4eS497RWMq0IyMC6WDoARSW6X9e4sZjSOpYVvHaYD
QcOpgLhcVeHMotfVoLldaUkl75v4Z89MTeSIofsC1qyD5cS0tbtJRV8rwu6nGeTyBByGqmHHy4dk
rV1M6MAp4W2GttnvIsX9z+0BOdXcoTOjWAjYbiUqXgOBfGykcrmHyKl9wyCbw5UPJosvjhstZgAw
fiAOSo1L7XVHsENxDXOToNBnjpQeNLVW283p9FnEbYnFfmsZyyKpoghfpBOIi34RQvEZopBCJNs+
/5FFcAXCRY9RAZcD0zIgPIggeXIj64hwAjzHCR6bo3V42z2Oh5lhTuUPxhvcZfnX3kOqTMdNhr2C
Rxzg0lVGfoAufwqsWJ8fuVVMMN0k9qh6TQfoVvQ54pVx/bQBi1Ws8APGg624mW1juO6v+yxM246B
awlJCeLjvrsv2vzTWbOuYdomOrsagTtJv8RvxLuV5L+tskNS4Klmw082GzxwYF/gaR0StpumTB7X
+Sssur9c24gQKyCs6EiCe1lgHPSML+SYgYPkTkREMLmQTjLbBn7MzqVp2WcbQdMOTX/ZEZgpVoSF
/U3zA2uSzTq7+NutJ+6TEMCFMNAuoFMHlXMoqu8X85C/5S2KGX4468+0sB2ct/tDhkN3I9ClKlD4
aA86Z5eDUfU01X/91kyw455WCsnmisHIw3gfNd+vLS4QlFW30995Xf2Ii95R7AQz1NDeUL+Jb66c
OSDBszvGiSYn2sA/WhAWDZdI7q3HdOUJgK4X9W0dCplzThaW69ax3dp/Paxbn4R/HyHucDS8cTLt
+++ijk3yCKOxe847roY515wBIOOIEzhE7lasFS1WmuZGMuTTpq1reJBm+r3Nz7ATtnjxCCis6BzB
PhTF/WmjoUORK5F4I/4twL8uNDtG+bwi/zGFO/CZDLQN5ls8zwvZM2HbFtftMMZR+FoghYbYxxJw
cSSySnIoFYv2z+jOu4Drx5MZDRwBFkULPYShTHSxrD53NyM3tzAaJvO4QS0szuTpGhg65C4oZXT0
Aa0CMr1KJqMFctjPmnaP9fKz+acBXjC6+hIFTeVXghRyBYuPLwC5aWHD5mp52FmRyfWCIqiC1QK+
LlpENMT8DwXcJsi60JNwkLZPQGdJQ3g96Xy+seXWtalnrTnWsisrdMZ7+R90L3JLrn7VuGngDBrE
/sfz/28X9G8B5M2D7Ynsgljjx1jGMMZEt65tQ+kx/Veyins039P58NowZI16gJpNs20k54EwP1BA
hgWIn62cyQhYehKWf3yNoAy+Hc4WwUc/7+VzExiPgs+KbR5cQsxBoot0vQCeifro07DP57kZE9UB
qSWZXoma8S7HoZpiNhU7PTOLQtp0fMINt1ewGmbMDxe0/t7dAqxiwD08zG++m1Kq81RcVeDY2Jzs
f9nnJgDctVXZhW0iFh9BKONogwRzp32NM1wlvaeMsMiQnGOp29AgHIJwb8Oa2dX6H64qoYJOAR3/
Olls0X4WGyWOmgPUof5FnhBqXs7fw2fIOGEJgdl7b1yaB/f0992fZ6i5aVY54imQKEhPPDRRLEPV
EC8TFOc7bgu5c4gasdaQEbWWzvpKQhSBberStaX5F+SDI6Op82CujYnh25Yur1Z6EUgk0Dnm0q25
1Sxb/j7HpFo1QG/5Fh68x42sNVz5VQ2vjMucygNkrc9eLZlJkRDKU3JLgQlln+V8ga49YspX3PYR
dSDASnDwj/KB2GwO4FnGzwNiF2hWSe5pC2GuUmYNbf7j2jOebYYDHtqCsYMsTip1bnQEBWORrNRn
We2s0COKisljNXFZ4LLOgPI3swn+5reD0xVy+gW456HOFIIS3x8ZYhGZ/GJxcXLVYF5UwvqoIN9i
R850VgUJBD+eofm86qKqcsIleLCynig1cYKb/xv+YBhUNUSRID5yBDU5RbDc+11szeQJXN3ab3ip
7z5AM7zs7Ogn0ZjGJ/iSNQF2GCbEIrp/3v6w8gI5O3kXa9ocMnHpiwgfSzUjrx04SdFQGTTjoidy
ERfFF2sC3X/o8FxpdtMSF6x4PrTopjvnlBlFuhG78qOiu1VUR0xIW83CbMxaqnEuvpZJ8m0T4yXq
I+Wa5mzF7hhWwUlbLPRj6Az1k+9ZPhDVOpd1BiKuywH2+BhzPDSq7aSmC9TPY54KKNclASJT3OSx
EU23J3PlZr+Hcj+0pnsWnIZybd/ddO0KvtpPUzJYpHWbxcC7FNZMJThzpM40YZjvetELUMRB0/gD
xclxfOJrsXwMRtao6Dq4NfCBjPcqqWJ1Lbv8DIOji1VkmCPiLU7iI9DcPsoat/7gAMHHhuhYSQk3
JTB27xo9lFLzsO7bJZBS0CkJeKMTqukCf551uciFDDazVmBhOnZZgEVSUbSLwaoc5ePDS2Vl3m0N
uTPIKYfP5eqf9cc/xO5wAdAITN6JLbUw8mPM3cT9PAT8LHhYoeZ9ZAs40n90WIEiVTKagmFrphmy
BV95ykd8INSg0wBJxaokehNiE1MJv4fQsSbCqETzRrBFuTLhZF9OjPwFXTyBQ8SkkyNJtJVqNowP
4FAb5QKULAEk4J/VfxULI/G0LGyhny9iI3WtFsCsrRapdtxvJBFyyyMDv/a2Ns3GMjC6xtucWVy9
jMXevx3Kb8LEBKRsGWAHBUqq/JV4kTauRUGVXiVWQfL3fGrojdDRDTkLhQ0WNp77K/nQBjoKb3bw
4RZzV3zSJThfloiqwEoZkjxoOMHs/1LAA8XHSDwo0I0sr0cDWVF/eTpVOAy5wohi7WmIh81vxlPo
IDrBFiC5poFFHEzHkJOZ/nT3g6d4plep8gVEH/PR4/SpxFlaqYlF9E8IDkW9OhzQcVA/FP4PAJVO
1fd9LPsI5vwFxYaFFawCgzJ21zGrzjMe40cpYlUt6nYaObBkcIVrjghTobzFEodj3sgjEhGQCmO1
nHtmLLz1m9MtQ65JaEMUAYoQPiyNG69WBHtKWBhIGpCZHrGW4/Nz5WTQsPt3RtM+Rcm+coAhcnad
pUUiTuL4S7Fao+yiiEt+L7VRBQN/XN2GEGTMKeAcsP2b/Lxp4/QBPSX3wrab+Zk4CQbcnKVp5m4W
7p9Np+a1Mvca3Gd+AicJ+ghGI0NIA8AX2r9KuA/3sd0Vf4xCuVBov2MsIh/6Pk//XuleW2taO3HM
59Zc1T7nHZ7pAPsI9UwBt6VSviUnIisAnLbMcK3EFtrQdftYnQ+q7Y8BleVCrj3+b1u8BGVJIQn6
+ZrfQn74iKXODM13MvzoFjpuejXsbhJ4LUDBmxJZEW7qpuasioG1XBUExDXvna1/YpuOPOJuz7b4
lXYctD2LHPEm+SM2T+QjUsBVE642w2k6oNrMxPRfpdH8ddT/aQFNNTnw6nv2755XedEgob32/kE1
r05ClnBKgw6lCRteWFhg6V4qnqglmJe1DpLndeoEgWyAUhIoenZmHSB40SELhFT8DQWCdmopdHCM
jwWVroTk2wH+JabeBgNJMpFFfg8DSdUo7pH0YyL2PDYnj6dOoi6zK2JcokdlnNExrlJclOXq+dHB
s8ilejWJPcHp/hZdpS4KTtVNO9JuxXziYkoZVrvJJyq/re73uB8IPz/MdHE2Vs1QeynjIYsEFA4a
NHsLvI1o36qJp/PrOwv8b4GT+3mpIMBhH722cZXKGwODFk0zH/RwaupkcLoQnVCyu92AFLMYv6GB
1VO4AYkIfzFJyKz5f5qt5YMq6CNk2Gh86/ndbQUMGFPQabuluEgUvpre3zj7wtc3I85zQeZaaCih
AFTX8X4lzBL8ZK6JxyGszz/ptDqQzlhHqAibtMqUoK8WeC7JQgOIR9hhjtPvRbHMfXCNnc08yJqa
8KTqaZCJv7AEpCloZOHXONZpciP8qEu4U9TJpYHiXpWT0MGHwVf3lndWBQ60ClotHCGzyckylw0l
TaFLpKOXccRRsjO4h2hW7gtyMr9sphDYs+7xO3+wBQ4byKqqkHJY4mwTPqeI5BrOdGIeRUD2F55P
wTCI1OoptQUUeuWTuealWvuRtMffGXkhIpVso1+ygYkVXMsXrNx3xTeblIoL2Bz7ekV2ivQ90c2M
Hqex5jwpz00RkEr9Yppw2d1hHN/YIW6Y6hlm1oGjVTBlr+sfgxQgvseNRftzf347BR/SkcsfCsIf
M4nhAEvGM7I9A1r1+6jdk9dAvBtOx06BmVCTg9txTAyjTStF3V5aqgCFQucmJg6G21wv3sBHWBTo
RpLbByTzYj2gshRmXSVWyLNgutFzmD7X1l23fQPPYPHuhtJuzVjbuc9Qf6REeChl2bK+W6nHbIEk
EuVN0EVcBcZH8CicXo/dtNk5uqNS9u0jh89BdPH2fGMDjcLIU0nQmTn3cPqmjISVJPGEFvkzd8xc
uIRCV44eOSqTzDrCvI4IJvVJNWhsqxLk3PMnRyjGyfn0weyM/3/K35+7SLSLIsrgggGh1OuN2t3A
c3WNYjxrcO4bvzcs+o+mtOKgxVdFTDekFbgRxnERL+msL4pG6r79N2WNAnWU7zvTjImULaPN2QlS
Nh+r5Im8m1J5p1nyu5GIm17SpUXrR0euU0GZ5lN5oHcQ+FrfQd69W2a0ABDwtSo4cG2Yu3lTCr4W
YxQ3n5g4eXVjC7qwGi+3u5PyhiWERhV417Uz10Y+Qzi+9ufkvvu3lrC3qcZN7NjFzXBFKOBb9UWi
vpXFNbnkhnkZSBlS3amrQhIppEEjPApemyhfLhLhnbVBncV8Vv1qy6COKLcMG2gQA6SC/wr+3sbJ
/Zfv3dpyuwCax2glY99Z0qf5FDpD0GlcfEjMMc+mWIwBW42ebL86ltI1d0ZlmlLp0XjNjkxgh4SC
Q4V/93bAsq7yk5U+B46eZRDB5k17YDIa0ItI5SzHI7pGkf8lnNG6Nem8/ISFCWEnSHgQKJdfPnXA
GayezQ45vanhbO9baKEPnO0LR+wEf23oo7LgPAerXy0qAQET5+fE7/BvqAcEHDP94do23ypEe1Uc
UMO58Gjbx0jK12OZ15Ooxld+Qoo/gSTKIXBwo/ioKQR78pKktxnel/YZzwlp79VcdCBpoWz9u4Gq
A4R/DHavsOheBjTFZrVJUeuQRufTDk2rgfJSCHt+ofaBUuNEhskqgNdQEx1/uElRjFADDQpD39RQ
66/Y0ggwXIn9tjCE9jTctZew2nrVYPtGX3xm8vrskhp1cXQuPEAz8mJqr7TUh1YOEGZOX5J8WVfV
abP9doB9IRs9b0JQLnWbfq8vlqNFxBAoYkmoWH/OJnoKVceRq/WPWmn/ZS5fYpqLx/qwQk9BF7mK
SNc81pfJEWcO2tiJr3YsTh5PIQTtTxkUsvIDUfz/GjLZmvzdeUY/BJg57fckqYp6H1qzO2xVzMF9
4f4zJGCaEkau5iv7QvUGUBpBmklXCQoHXF749/36KfupUMKVEGmA/ZxgHNYdV1CTyZXuZgOKkwoQ
gQcXLEUVQXXjbSVajtmx8uc2rmKLFrOMOFCgNWmM8Rhy5ZYy3Gqkj5y5xVeMUwZE4lND53yqhOsj
b6hciWFdHUubmvqrqfHE9CBBhBDYTBH7fBB1F5FOnZTZK1Ay4iTOGWmtQ9z4y+tWASXzG4O90uOf
jj+ALzLsof4uAyWaPnN0FYgQiGzX5woDsftw6NkGrEPROhpNhXOSftjxuFPg6DBeQrUqeD8YHtja
2tUsVL7LVoDkPdBCJ2CsHzrFWyAaJoMeAIHIAVY5dP8Ngw/+11td2aeoWWVWYV7lWBmpH4rgPYVI
U5aVzKZao3s/KoMb8pNf2kLpg9uaCE4KvAzDrtutwXchSZk7BOYcN3gxgUSmDgg/8SX4Hl08Wju8
sXE0qeUOmVFr8AazVRf7E5kgHVO+6hf3ci85NMJgfMmiqSZM6z8nN4HHS1KcV0LmzXWdHIsypeVZ
LjXSPCRrE5Ls+H+Vqxf5JvvMec3XdDNapd7+VW/1GKCVuDDoS2aLkyhiv2lc9jnsFwoB4jHEUtkd
7PXRIxe091aVTucz2pYxS2SG4tZMD8V8zFqGCnfhLi8YorEpRhvW3Ne5S61S9g7+PF7691f/Cwzb
yVjWhZV4p3Or84GOIVZtc4h6+RXD2ZE0mTVNJTEkPLCg6n+z+GHnqwO95z0NRnConiS/53+KN7oc
GJF3XJ1U/vvWgYdapFXIFxCNeaNfNv4loDSMJ6mBI5Cxi3kFcQHyFYbCREAWhUsRNkIZw5JLELX1
1q0cVDSD0mjI2jn4qZeGa6cOSS+m0m4wwCH7QRr16tZB2jNBJv8oR3NMAcoi6FW3SxVz1XLIo3f4
T7DFuLXIT8DbpVMP7L4IK5MLq4G2FxWbVo+/wO/L36uQQqiWB746PCThOtC1E1+9o6AjPX/FdrDb
wj1JqeaX7LfaRJ0Z4z3A8IPpNT93w08T5KbdtyUUGQDZmO1qLss2/nOTZMJGv8pGqGURcYhG9ZYr
K62k8vASvfUvEVW2bfD6dJ+/LnNj+j/U/rNUTugn59+2hO25H6PDkaYJqdXHfZBFxZcZYn7jyTGz
sAK/HwwbfBMRksnYa1OLthTpL+l2T1kjWEGpO7wX3IsWL18LcW7Do6aO1kMNGbZyKe/lJ1OtAzbD
H1rgLppe28jj1gi6cq2kHR7zH3taVxxkS5CbpUqTK10Wq6zbE3w7ACv5i0p51NylGg5/TDeOdM90
Ps+kqxcvr168QSgUg1febuhyxtF30zo2Iz04ItyUY5XzkrMlAS2k0fq1XzXtKXgGpoX/josmhq1p
EREdH6Glfc1juwp1oMF0Pz5Q7gS2QdJWLOs9VQw7scJDJ9ZP9PAHwWc3zoPW5OP4ueqbfc5Eaakf
5Yo5TqfGPvnnz9kcTPPg9tb1NBPlauGvu5Uqf54Qk5Yyt0YQ/zTjiazMcA+W0mXf0dXXoxljLJUS
Ht/6BBGWm86xdnluhNYY82rCS/Z/eEG7mbGl9qIISI07QezqF229Fk90kHFAjXdaTYt2HRgDEcN0
OYiRLjyk8LuN9Zq1cS5P1D/LOkSEm84RcqKXakFxHYoMJZsUwwO1q6KnNEv0M8A0f0nnl0osnV0a
d0ZvXGXmfW3gqvr39ZT2TECJfopmmqYSFQTsFqkcaiJyvvoAO6Zgg27tRNeIg6e1dvngAwua+7Oz
R6iBbRgBnTn3vCQwkMGQjXAWnWsZcepHOrqLEcP2TzTEWLfXgeQk+qe/yBI+Ah9U7wpn7dvRWGUE
c/WGsViHV9GYDE/xrB7GWi83VyHHfUfidnyodnyLeaT6jupGfNJWbN6QEGpQfJIVi9DrhtPsCimK
qjzCj5+toLoMsYO6QKHqkPVLj/PRRofxjG+oQ2HrqfvUAiRsJknZWdcsJo14m7ZJ5NSy40mayzIt
aE+noPpn6dt+j9xiQLLlRBXobNEt5zvbn4OZSFFK41y4wvyDC/JJxwnqdxsqj0qtfSdhq/3u3/s+
5NmDbJQ3LNWca7cYrHhftIIa0PHHR6MgedrHXE7aiMiBHPuSG5lYNK4L+R0rkuHbP+/xX1HVBEZe
e4/L4keNdy3F15zQpY+KfvvlhTYse8FPf1TmKLvVmDuXL1O9ZqwN+PT/BDGCdMr1+re1t1gvU7Ox
UsRb65D3Rpja3+6OqSb2HMqefepW1aDngiEuy89kFiLQnKaB4Z/cUke9jdiXZt6bDfGojROiT9gI
W3fHfSUgZqRrfQPYXqw8EIXnKqtH/eqhYFArzuMtdolRder090rnpf7J2XGRUK2DEaUFu8soSBoy
w0rVL6OMJnjgm8x/sGuiD+2saJE3QsxjTy1LDTYEl/DPbnxZo8cGlBERfKBU7Prc9B+ubf2wwNVc
O7vhW1ZPdp8KJwphO3V3jlWUkIio1UkkTwpjaYzL3VEtlH2C3AB4Zjh/fMSNVeOa9UWKGisNo0Yi
Er5y86Bhq2nr1Jp3+QBjxbZ4BK38BF6vwIgdJ/+ChcBXcaB+5/MLk2rNsENkhfUfcU0OcLVLU03T
HcBsdi+ibTIo7xLlrO0lgzjCu4M09Ia5b7ETYhdN5vTb1+Yw4fZV6fHxCDj53EmeysY6bA4XW+6w
heIwFvOykl6lToE741MIPD2mBEMaKu8HTPOPo7BxZFxOvDiQRhl/9TXTwPK1klECTq98caaMgLBw
rU3gO/AacOPa0sRixA9AmuhgZvHhbb6D/eXMzT6ShZFQUkJow35Xs5f1IZFNcWTS6lhZ51biBUb7
QQ5LP1iCn3tR6PAb7X1eEGVN2R8RPFxXGvf5gaY2GrkLKLdEW0iUoHcyZn5jYo6LSLHZDD0mG00E
k6p1Ja4UI4wbCYJbd9fqt1XQgCxarTgYZVz/wRrUTMMkGr0WalF8y+0sQDG+PYFROp+mkl0HQ1tU
aXhVm5+lmk/Gqt5VNmGSdBnNuzfegUbxzJdIF1b0IVtnkZACQiUCvGzxSEMl1jM5Zfnz5KwWcEvo
57kwl0qam8I72wJlQtlx7iqKD430AynpwXGQRVyPYSbSadEMAP8nUIZFm9D7v0qdWweiVmRkS1XP
PjeQ/1a8bpOsCmN3XYcZoPWPWOvFkt7fPmvGJ+T/eV3dVdvwxAvv7ZJmvdaf16auB7l8K+joCeVf
Uukptxi6MjA+0l0YFJALePqKbaeu4W6WG2S3DD9C8yzVfYWmuaW6x3TlZ3AWBYxlHhj6D8LVPa1J
oRmsFGPm7uu1ff+87b1Wce240FJgwnjBJCKo1HJpXzDJesnld35TFmNIsneqTo7BFsnVA3AW0tgs
+BNa/GnQykImyoDk/fiKl9FqJFGZojAKf5DRdQ8L8NK5/tS9U/PdVREPT45lO97T/zRhJbFuNHv0
NC9tisIqOQrYgmhMSNjcvbyb3iMzsiIjZoTtzlWslDKanjCSFGXBRyBQ0Ys+T2sXIgIerbkDjPI4
H+fCEjYgfBJ7j8RZhSnp89ozd+7JlfM8dmKc+NTktIumnwdPaUtLFDlWWdVyBOv+EYPHxE5iiOjd
prn43oZ/7QtYq4rBecw5Ugxj6HSORR4dn45Gb1IiZLkXkK3VCcJ4oujn8dtgSn3jeQW9BJ23ZTtc
X56p8towx6LdNW9DmFH8zXevz9Lor1eWGBL5OQQUW6umxJO8IrM5VbZHJ0kekOpYcA0u6HPsnoC5
9YoDtuZaWgklFQCZlq87tAfbITd9KRAC8zFY+3VEDDURErp4fwWv5NVuHQLgmq2Ri0HBzwqFNwie
gQw0dheCzlBO0EzXMTA6hGOMh34z+Rt9fOWHgrDjzcCO6ga6J2P7r7cHPJTyFqf1Xss87FJhZzTJ
HiZd1UR9BGy2ASQDfelCQwpVlBlCdiFKdjCu7lVIKX3lHhzdV1JssOma/a244HH0MQsoviP+CLWP
wFgdqzhuZV5Kj2RhGmxEVUasViozZDthmIaIi8hu5sDY9y41SPv3VVUN1M9ufSBIRtdPrXDB85no
aXREKa1EzkfpRKjqSVzbenaojb6l2+3S4VyhoEnhp3l9COjm8bKTj4p+uVMS4o/+RtgNIWqC1dVX
d2JjD7M6oy7zBvs5J9YFEcvBZ1m+wLd4zKZ+6qQffqATUoLUs6dwlwvlZ5LKiKrs/iRBKvti9+PB
fxidwe34VbhuSocnKVwbG/tbwSvhMtlY+sKGRSSUABEBCVjKWOmKHwzIETmqb5Swl5emvzcAIJtI
nUPwElCbDWRptghY6XmFUmzO3wyVF/igm8/AK2HDVZN9xwpMRJxa3xc4Rgu+LPTF2QJblhaOxeLY
AlBrZfF8i3IFr8pHxev8Cfj0FKVNnJb/w9DExfwSjZcAmWuc2Ez5mVLms3XyZHCWCWfYM326ODHj
+Yi5KGzEhi+rjtVs9P65W9SE1HQa/NWcz28RAOKgkrfIintuHzj6ZmTFm486mAlKgIWttE7BLpBY
MXZh7wF9D+I4r5rLsId2XhaTgFJtV+rGzY8ayNDhtzAhsM2JHbSIoynS3MFVzEHe3x5TjQrxMUSE
Yne5leaMPZa4bYr1a3vg0bdWtnMEWHpMQ8ba3UlA9cgEd3RiEUJisLMGTNBYkzmdzG7XDNuJ7onE
QiEgbNhvbxJi6mg7t377kXSiDnE2J598MnHkb9pIkK2SWMYmOe5JoswyJsP7uKYA0+8o8SXOfutW
onN07pcrkmJEO91saCIrmY7ZCUO3zKmKY4SPAIYlq/jMOH/Cls48iu0o2w84uqSszTx6AZhFEGqM
8yybKs33hk0oxqaLFWgl1a53E8bNx7TfSOqpeFpFhq+gDM7hHl4HbY14f0lYvjcILy7n4ycJVU6w
oMRhOwqi/UlBg2XwAxSQJfsbjrGyklMSSdqT7FMUOIE0cOs+pAAQuWAROXt/23cA01S1eZZf2gZn
5UXF3FyaSZeX5/nlC6MlEtW1309JcQMpYugtBnwHHabYitLg+0Ea5bJiapLqJXkysF37wTLpIqqZ
qsVpbAiQkbrNLHQhvVqlbh0lxhxlGyJq/sk/DhZReTbmdO0BjXjZ4lsVgcJXuqpi1xJsvs1SOu2J
JGUr3UlTAsV5UhDLj15xr910BmPv/O2TN0r/j6ovTQ3v48flgext+ZgzYDF9mWpTl6FD5rClKKH/
xs0gxiwqwfozLFSKBEFIttc6Xcr0xy/UJDH97IvTE7cmBUwizWVJA80fcXRbYDyLwC1F05s+FDz7
iiNxa7fGBMr7laXqONcm+ig73jigpd22qMee0sLSLD/GHRgbgvk2TvbC4m236+5qSp3xtUWHfFVe
H0NoqwODilu3s/S7yhZdeKSe8xq0+P+8VOqBUIWPYenJUoOgdxFkeryxrDiVSuE5ll2iYMi2xl2f
BIXmoNoAlzsq/LfaBtnDrQ431+gEkM9GGtjm4iRSE4GWlrKWZDzcNanEJ6iZ6nP1xihsj+k2ZtvM
nuH55Icfpq4M+vIZEKCuoQ391YVt9GngREoj9gigOLN06t6HdUoYBkrdz9vIqqp7+3Oy4aKGyuDH
1NWHtZsZeehoIpm7/xG0kPIdMo2XOXPUri81LMB0WEaSlhYEU2BW5RtvQQ+8foqBXVSDCJkzSS4X
9F3EC+faDgOBlX+MldK+L1QF1intRpAwcKV0ydkGHjR6fYWa/FwgkyiBBbPCOFpdTJjjXpBju4K0
Wj2EAproyiv2HFHbTkGDU7736WUTnwcHF39VzG7r1+BG32LaU7ZguclJi1y1syYmx6FjpkJ93ZW3
e9iGfLpnImN7qVjKAZRvfeR+hSR/zaYrPUIQxb9X7kcLL2CikzAjJD5eAI+ZMcHGOhx4rpsx2I/w
cVWlrIMyTxhjEJDrN2DxK4b8v4qQ9BEJ4AxPclorMKoeZ4tNh8ETJL96eMAsqwNW6dwD0hPu+r57
soc19kRoAWMIHLJg38hjbGiovBO8Uc7V9pgjv4CckmE9b60r/BP6SMD6Rfkw2WuR39pYg6SRcZUf
6mYMr4w8vt3cyf0lunmWFUDP4jUB2K1p2MY6XutN93HP3f396Do8VBtxDX+nSTv9VUCZb9wz+s3G
srWOhHaVL0Qh9OhNt6RjysOPM1z/vkQBr9hBRcu+SXXFBL7KlfL2ijfF4G87ZA3yZgSn18uyo+pl
Jj3sLCK7Ktyi7xf4OZ+8hm5lGparx5D2FxpcP837BYDwHJRP2ql9ECRIBapVFedHr40x41sFihb0
1qWes9eV+GaI7wV/qTvW//+DstjkZWNf02NBKhEFjVSFpeRISSwbOCNjtfHZT5gH9Nbk024g9/to
109RjROiRhyyX4oLaAxD146R+gyoYxAtcZIyoIRMzdx/eQXX4Eag+0ksFdZ7mJzSf132NMCWU/uo
xZMp9HVFGyDIituUhvldvxrL1MX9Z/wjpIga4GaCPcqb6NajamWsyl4eQDzOKOuxI1uihFSlDxpE
TSo7Pu7oGtabJAAzStbZLerb9jotyo+O+FrPCTQpDqh3N8m+3i+F2GNNIA45XZ4qcg91yq/TOajM
HB6e7S95ghIERh4Ed89r+IS2M/KbU5C179QbBiTLJDcmUxNyWA1rEyUzhLjtSWxdccehfBAYWr34
k5zyNpYEhd0K7ojxayKMFzXKVOX8PeBjO7cCEmvOw0VRLXQEg3aFHp36YAFWkinH+HS08nM89Snm
gmr2YFpBMJi+JyABRa9Iwxg8fWKcGMWsXY2zACKybw+BCgX3APxp5ZbVzJvC4djYSUNL0SXpMsoK
mDk+hHc+asaGfhAm/6YLc2uJR9PRfynrQVslgRXI4T3uAYVT/GeM2krBbFxsfq8BScUaPOkVk0Ug
744uwOjQXqRTvbWlnpq0IRxonJ7DmSGjnfDHqG7dYZky4NVhPVh23BD4GFTW28RywTxqrhP0Opf2
8rvAXIofInNrB02QKE87rs+cZITD4PNSq9KepIWyjmP8ycvEAVnsKs56oDIECjHt6WPWEoNRREGO
fgV9dHYx5zH7580qd95/D1crSD0yBVtZJkruYVcqxReETVXireXyqpHHoKcfIUyVmPrhdQlpX8jD
074AmtcfjQ/Dl6Td5mnvItWpkumlAWFf7m+4+vMguicEcKfNUJopJhK64hkTPqTMARNpbaIJxkk+
rVsPWlYAuQTbBib0X0aVskrKb2K3Fb+lZB9mViduoJmlgB5KzgAhe0AlOIeyh0xTmz/jsggPVgxb
jrkGZctHrj1fkNQr/dLO5hL6d8L+PonLwbQMf1HeCM0K01yr4tXhVzF5eV47cDPQ9s/TrviE75Uk
qPQb2YrXPP60kqTRznbAc0LF40jMV6EcEFItbMaGaPFMLLQ/3PiNcjYac/FW5Dl5QsFnXiniXTgW
5jYwzDXcFTzabETjZ4yqg82XSVXrw4A7P1u0eKEpO9qV9PlOQQpKaba1lfYB6vy1tvv2Ktn51glz
poz80yZJhlx2M+zxQNy2/0OLkJ7IZiOYHxzWONf81KbVj6HYLs+kbpC0evmgklXqPogLidxxNyhW
7mRY26rqt0j1HThQ7U7VVJCQzO+WjHqbDCldPfPAASOBkno51Q8qda4uS8UFcSlNq6TdSfRjlUAC
Q682rVzKYnLoI7pxu02d0tuuoxfjYyb0/YSe4g63BVFrIvgUiKAPVa/1dhgrzWoWrpWapYl+a0nL
2peQAImLtE1rLJyaJMrKXVLKCHEsmcL95jF/glPN+NFuPDmrtvgok/YutLKjiAAyYyOUwh9jbKM3
xSdgLA2uVjUbN1OgblbxvFoYAr5v66ggiAGnrafraJPaq+/h5qij47mv5X7RNGVb96zjK0VI7jJ9
4Qu8zD8LEVmzluD7jFV1fBdcr5INqGNzfs6+fonPJ5b1Ly9/fj0Vx0KhruiNfjwdBcmUdJJzngPC
0ARlEzYUm3XTlcSNc1XpJLYX6RYX1NaiCZ9fDmgdGDPE52RwZhXrx3OoaQ+p7KP0DHl1GSX3iZgK
BclzwzW8ENawgx02c7AmDcJWHy6wHVeYnZ7lm5uumyMfDvSkTN9FFdSYYnB6w658JMSeRun30rCX
5TZOBkkvRVN+bPSQ1hp/ig4im2V2BMf2Ifz5fm7DYSzwJROwYJFeaqpz4Q/fbIx8IK3oifNMS9Cv
2SogjRfdbYbPFe0y8AUboLrBZSbAppAKLQbHAHavAVVYXebkn6y6h9cUR9W8MiqhbuaQfMoPagCK
qg4wmDMLwSeqAQbzuAEjIEScMpILAwCy6PHE5VPK/FdyV6iZ+iglGOEQakGCtDTuWnA2ioadT6HH
yIp8bhhw8JXahdhSbmU8/s6hvzbkyLfcLBQno97lczgrgrfD2IP+AMi7aBB+LDpDfcIrsSnQIBZ0
Xjlrao7tw73kuK48TPoDNRBuunOE+39Pe+Eg04u2Fd+srnui4QvKhLQCdOTGjXXH0LsPvkytjeaD
a4Hdyb1TAmB57RQpoz7gMdL3dZpF1Cocl5KnyFpmuwNX7ZM3wnTyoF7bradLWxXa+u50yyImavIX
18S8QxwG6O4IklljSjJqlxJg1zWk0erHdf5THt1Sq5aJC3j5nKQWL1aUTYeHhchArRQlTJAe2rTH
TFSgk1Eg1h2ExBHimbJDald8v5Vzq3JWK3ADEPUJW8opt+3t4uMZfyBcPsAlBUOFs9cei5eQgeji
PRKg0hYPmoL4D02+QI/HYZevTAYoKQ+sDygDlIh0WlnzU5EQXFfFNKmE7DHTIuOoeGxlW7cPVwV8
2y9WpS6niReF0/44xzALl8u+tjcfe2XQrmIywq51GfzDFMy7SshbDkDgQUPi8vfNs8ChxOnoJUuK
p1PA6TSNB4ooL+S5jGaSDqj8ynU1mgyQvZDPi6eTEz0wPB4ls+wOG1kbKnONkjihcceCFbJJ7h7S
lY1sNSs6Pzx/8ZPrUShT9TBJp9u08PD4H9RwM7yLq+N9hzrv0CYtjddZW8HpRWvaeJXznXGTa22t
PEsOhXplU1pO0pwFOaokCsMXGZ98mh6fqWOA0t47pmHB/7DY0dGGbMevrMmqD74mR58dh7/e1rdU
onsQlqfOHsP0DXXRVjyHTxFG3FC8Md30bJlAOGmiHDl7TEeUnAzIoNaH3b2w9KC7drQVnAjnaKcw
CTqBTAjtDh7Fbnz9ft/fDWKCXpJXj8Yn6701CA8hoaxyyNFcu14NeG+JA1+Ca+KcHagdsjb18TSH
1VPthx+2fsETCNQ4rPg4Y8yt3QB86Itonwul7fKqAC84fSVFde1AZh1nCjolNlsdfBH+30r4ijfK
WY61OSiNstN/d+6ViOau4KUkcGAaQpFjW6y0KlK1NhgabHZHdoSbYNpDDgruZIxfbljJ4z/A0Zsk
sPXu+9kMzdY96osaAc5AUcr6uslJSHCBbsuTOUcHscfcAca0V//QnlF0P2fEDawfJLO4yqllP0D4
1jT6mhnAkdXwPRHpNPhyQfR1cT7824TUScxB5M0vPVgKMg+wFB0sS7fisKJb+jJXpqBYyGcsLETT
TYPIPDAWyODDpIsSurS69AFhmd7GcXbZBqtvlBM8rnqfmIu9xO1hwoARmCgAD577mcikhSL4y4W3
UvtqV9alvsTxtGHfepr7FKaOv9h9Wa6chqOL8J+cZJgn1sPnrqaNrQwYP+lPHWLRK/luKr/Rj8hj
ujMqtjySd6iXGdJ8nFqL22EqmyFaBTFFCG00zQwHKzv2CMo1sHUVdysptNmbU00ZsQk5zgpkbMeS
Q/LzcrBlGlXA+2TJRNhzqWSYG6n8staBfNzHwhQP+qeesikXpeved0ccoi8WhKpg2bxSqtLtL5eh
uWLuxmTb7jSALeECyka9m8tVelhMlY1Yje3JnzjJ1X1pryUIgtQUGJcxHGT1u8ZHMj4BC8t9IPcc
Xlv+2D9SsEVMiEVgO2OZFjVrefULh2daQE3y846jNyzzIK+j+2Sw8rgF0nMRVbK0I3vO7ySpioZi
9IMXbXN5RbAx8wU2vCFnYH6+kllCp/RqdRIQq+hD8wogwi1Dp4fJDbP5PH1GLhmxDb6SSpa7ytsX
wSAUx9zrwE73naW2qpD8ZWTIdD4IwyxqEebPMqSl95MnVvXfYomIBWIQ60o6AYkESgFkP5qj0XAn
w2AmjbCT4zIF9D+kzlj6OEhBBaq6UFkOQX97u+fOCdpu9i+OfeoAXqjoIuko5U4+8FkfZH8hbqWW
E6ALrWmXkoPO0gmsb7NPrObT/FkrSngzBqNnT3AYhdO0Jwqldtj89M4WkqEYa2lHENlG9+HmLKzF
bTvlHVBxmGq2fOaZCrcIodN4uOrV8gcWIKMe0qiW16bhabq5VUfP9OzY0B+YHSe1KvNanMrKtewW
SAto9jJQjOUHnGRDZqcBSF4wGh2lo7/bVymf78jCEmgCvdN1RQaQvZNVE7zl8XsHI9PNd0bBLWSP
mMPkNgV92ZjThnaXCK0TnOn0zJ1KAmb0CWcSGQsBhz/WbMOsfpodFV+mEsR6odW/MLSwhed7GH68
aK3zKYAimnshbMplkPrk3F2L9Rmt5UIzfiyj89BS3vJ8w+oF6niWLFSxnAtvg2Py2imav9Qfle/D
kJqz9XpQ8e4O3rTT4Ojwl6wGa9tQurqNFdaNbmC2ZtHlJ6Z02rWXYFTJ+ng2Ns5ggxoAD+nXkn02
SMv7WrycTlBem9oY8eCYRbkgFv7dxiwYciOSNjtbJcbWCr/FSTIIEAWjYbYeEJDwJtmpY7fJRW1A
rUkKoqXtAbExdlfyjn39T5IiwtG/jR339yzgTkJtnMMTOGNXTHkCOkExo41Z9GGkmgYo1hJ9mVr3
U5menVA4yOlTsw9SyGESRHWclA1hx4Es1FUMdUSmbkhGTOgiYnFwEm2MByUYkoUcZb5SPTZq5l9f
Us/AGnpIvLL8gF+aXUwuyTFDfNvCGhHYiquVt8stuELa9K4Zo+llRm4YWKWo1NPx3OgK1pcDYkkx
/zkndzeVzPh6BIo075DteowMqUv2getGQTlOfzaucDoIEbYaiX4uvdne1mpojxDWSEYRpWzooAzr
XGtlw8O35sl5MLRNoRG+rup7CjjgxNY/UBx7j4Jc421OZqb03aQC89wWy8VBcbrcMI44Mnjt/aGd
WFhGf1dYQHZkd6UfcclhyJWIJ752TIBW01yygNS4lHTo3nvxelcH7nJKFqy34Me8SZtRlTTgKNTT
iv0Kvvp0rl/bCKoBVT1viSNJkBroR7r+CNY9Euq3MB9r/oFcSGsvCH1YLfL1y9ENZp2h5yfIHct6
FlmlpxYcMrmec4SqBOJP9qZKrY3IOxOjSFI6v+Zs8/T8pQoqwJK/+67AEagC5xh9MIT/JNRecGSq
CvBi/us2Xezw5pB787Q7MFsHt3FIcZ4cdqaebzF+DcijtDhsUE/IN7Ky9wlDzdoror37eGG33F0X
hGyYAtgOemArlwZuj2QVpbXw9kf1ep1G+cnPO5CEsw+v/MFkQckcR1XjFbNVWIp6VpUHp/xEtIjV
Ajxt7gnWBsDa1i4zoUKQhvnsATtNRueDtILexC+dyxYWtG/GG+k69HXuLZIGe+QsGs0XFxMawVuj
+vqGH5M7kz5Y0ZzZEiZeXlCkQUKs88hb/YGuebZiKyi23dtZWNA9aMIB07lUF8qFOvINGGrh0TQK
mwYa2TU/QSWN2ONAvr5kUIqeXSB15FysWxzUt31xzP6BuEeJjA8eQqN0c9VDNKh65o/1vXM+eb0l
GKi8lbX/4xx0ws2QPIB5ddnlUgmV+2vEP6Nd8K0KmB3sJXjYBqne4geLkQoOod3AfcCWhb3ED8N0
3kpKdnVH4kzRR12f2sGIzdX2quj9kr5C8fLki1RZBVFOlIGcfoQ3XwAPYknIr9naX72xkRl6u9Oy
JKaMgeFXsCEFx+OV+hlI/05gDkvoXRG9fUwlkZooFEmCfB6U/LNFRRqmvS5TgYcUvjXNPWkpv8Zf
mzJSfXWXVchqPAZxdIk7mbImM3IQ1Sq6CjTpsRL8vwlUFIWw0A5CS73aM/nzvudFhTFv2O2bM5Ig
odQlv2a0IlEHUKpmLSSuAm5aE6S9qdkDwyAI3v4LHEtupgHzHmQrn6wbtKkAodK3zh8wgSbAPAq1
XkDjDzGW0gj5Ckl7y2G0NPjBWQeRto5gJ2PjB9H5MaefJHiwJdh7g+1E7yS0ZaXDYV+Xa3wsUk1G
RBhavp5oYyoRoy+uXFXqsEVQ+txNj3A7EqOolOtfSVuEqQBs3MVIKSI86oGD7+d/o/N8HQLEVy/+
sA4sA1GyfYeMeGiTFcZjCXrPVBpeZPb/d4UEZ0Xfzw8JlqaQUPGkYqYZSLclXGBmODWLLYudV3r3
fBQQ6r/AwM01PhUfSel6W715vffB8Zhqqytkrjb2yCdZnUzDrgbysMtWI/k2DIe4hJmL1XVFp7Ou
ZUqOw91q+HqWPq8fqT8rEZCqicuYuHDtPRcLLhR1LJjD3pdOW9iSs5vK887UcsbIpu8+FVtJLJ9g
jz8hw5y5zZuJwJWaCkq/mRJMiEeM1bcRP+4CVukmJNo8N7IcpY4v4KeWb6ODZAz0Cfrh/pYx9Bzt
2T8bTyM2xf4X42EQP6cGm+7JmTtDk84D3IkAfJmdNmJKROWHl+WPlWSMdEZHLd8xmN7tbRns1/IF
T9oJvLAw9ZlJw2kqCDKxtjRhfo7nWWE0ALNti6xy5E5goEY0qj44EYY3ga9jI1M1orr6creo62I/
WWxXti5ivIim1W1/L7Q7VZF4M2qDP4kdERS+dIe550oE8gkxsmaZVp9voQspqO+Psdk7DXWdoRyx
WHoqgEoEDqBuvYU2m0py9J6jRo4YEdlvKkohRaK7EHLEaPdWkiSA5Fs/2XhExmMFf5cbUJxe/a+Z
L1F2/2XcKsOUE1WS7NIlyaUJnTdBr/8BUrcDJ75TO38Rpkc8Ng1TPJ+7dDeEJZeNIfC2n/EIso+E
//eqemglpqr0pYBg9VZPCSgZ254cRFFTJfVR/C/xeM1G3FloaRs2Z6BQBDfPGIgQess9mv1P5g8f
mShCRWQDgHoXeI+mrvvEoykk0IVfc64rxr2lf5g+elMLeSaPYwKBG/yVz7kL/QpRbniyqoSccugx
BJJZQxdMuqGh4uBLMCc5Mmh5uf3wZnFrrN0c6BTzYSGxXSwb03rMjecat+7CX6rwdVvQOjYkOGrU
SouS9EtRDaT3fbTD2Yz+AI9QUjfGPYUtt7MgjW+zyPTU4rHWRYyqTGViNg5IPvpbOgQGQC1m2MLj
1irhZiv9xHPal1whobRzPbyEKkIvSdKiSYH5NGr5llm2VY0C22AOHyIp4XGTsQe+rOEe/QUH9gxS
eZ9fxmTY0cFGmVa2lfff4S4T/ExYFsk0jFpMEGklHHMSmZjH3Dsocp0ifUw16DF9n3fOuWSQmgsn
4FdDcK/J1k4Kay2gf+iv4ncikzyj2ZJsQLz6laqyyD41iiW5vDJvc4eCXgvNjxvfvvLn+zbLP8kR
RaYtDluzM5WaUwzOHLPDEf/USooCgbRTcGu72ls+ZTeObD3Ifb10C4kDLi1Je8o0/jpDHT97UAbM
MkOD+dzHXogp7DA/LhC8ZKNCc9SeVGGkMPVuR61evu8Fu0MC5NK1CX98wkHv5B0GTjf7oHT24+8Q
NMhvuHxKKJjfa54mX3VQQPslew2Ixd7Ijrh5aEyqkBEW3eMBkFLBk9oNxBeIjcZNVNA5QuwUraii
X+YRW58jH1Z+ZN21x/ARz5La0ytM5kB3bWEGl4l+eFlAwAuascdxv+HJMv0He7KALF9b0n9mDDAQ
PqiBuhU8IvHKKQjgScRBnZbAPr7SrvtvyA4psP0cdMm377FwoXTCSPi4BvS+mYFdyWpv7LMaaqu8
wo+/+YlEudmScOtvtyoL08NqqdMyDABFZxHAXzGbJB3z8/Re3h+9uraFY94W0UtKCOB9+vj/qnA0
SXOYMvjDeV89ueVs0LS776lY4uitrro8xKw2AHU2caMrFsew1k4gZ4em/TiKgJj1Dc/4HQ66oHpb
tYT8XKf/Sz54fJoNCOsImsAqkkwg8qxA8P/JroOVgb4eqxy+ZSiwvU38BE2ydibhrJyj0oMk1Zwc
24iJCJS557fBEGhHZL0Whklu4WyXI++2JgORpBM3GZssaS6WY81JAzbd2YKs+lpXf8vYpSddfsG0
hrIKc3GQWORjUbCtjeROFagnTySzN2HPMwAgQa4N6lZMYlwrK/LcG0Biat4EqXxh/jLpBrEyS7oV
2UwvGKyyo3/e3d8KUSo2gea84sLwBGrRu5ykUR/lPIQ73rMsYIItbW+a/5BFJY7mKezF0y/phruN
bOesMWhwjMw/PqvfgM8GAm5k530zxmMsW5D9vgd81Pkv+YLZ016QE4HUgieamgp52OCXqd3N6iEB
NMpHxQH3K8F0dRwJicrtCHwqB1gBjV9Zl20U02AsIcCWZ8YJAV4XoAddhjcigVLrWT0tIpFRQJtb
uq8iWD6n0RwbAYOsoeMtydodODWSDAQPAb8knLxWlb2qs/ebM1EQrkKTc1FwlZngQL2GhZyjH3VX
klHtQXbgc6EJcCBeNm8LutAH8O2TWT+/wrXQIjlR0IqRLw8T3bvEtJg1z+jGC7WH699I8tyD8dFT
tSf5fEAJIwYh33AIeCRvt2Oo1M/IJYJd32QGAWuM0N/Vz9t47WXBkFKYOGeA+D2PWR9AQmz15TJ1
PBrSEzsfoDh7hRStZvQKEEqTldo88LRB0+sldmAqnX7hCV+x4jyDXAlvu1ljb4UAOWmfF3luWa5u
Bb6whSelmlEYLk/nKCA/XloKxpWW0IBOiTf8lug/TG8JzmLi1skHPZYsO1yZF0ITKWGjyxXt8gTd
9cWN9OSRWzxcjch6Xv3Vb1/ZtsGAgwtNhCnxoWKlV3I3baQi69wIA+D2sTnpE4Ojl61frvqW5SKS
KT4iVjP0NBhCEYDHFQWDo0x+1JwxEv0NADyxVLf7G46vPUdEFYAZSIrlQOXtrRMKm5kZam3qZPw8
Bd7I/znkNTIbZxe9uYaXGw9q8nMDT7GjanQ4PZXEGj+Gxuy6cqF6j7js9f7TAAicKVYt7bYYu9ni
RtYOjZdWHBg4b7QznDfaeLE5t+bhUFoPB5WVr77tzBDg1nOYQ7JQPDHfQhoG5xS9+yC1HMjnhZY9
ptk4Fx5DWcwFnWHI3K7nRrkSlMpUYmNIQwjSsQsIzToqeAegkL819HOsGOQ7fIRJnNfR+fxaq7qb
+BMRfKhecX/JpTpax6ZIlMec+Q5CWFRyKcsUql3AtdHue+AnluNHVhzgCIc+qdMGYsIJGjJQ7/m9
b00c/7/avJLjiQZ1ec4wsi9lWDa2VkmYZexLy2nWFHF6RNILm5dCVwfJ7x4BknGFkYHsMI77k4aX
VigH4SjxzA4hObtS+y6VgD39sFTnj8fRE523xmUjK8K50YyDxYH31BHk7MYA788sIWz8hEDaexoV
NVrpnmv+HxH6/MIMrDaZhZwhD6UK6xWKLdOSVxsMkRmQkLh6s8y0rYZ476OAvrcfk8MCIGwt40po
Pj05Dgf+nEWnsCJ+m1OypxAsfFdpPaKFon8hlkCOlUv7tsFtnCjXME/WxY0cdiLxO2cJH69NhLbv
+/0K6waUbM0KgHqoStgde8HdAhugeO3/zZanoVMZ2yOW7l1Bbp1+fUaatYyeHZBtYe37ZHFXfxL8
+Z8PfhgX3vYTqqwwl5Us6AVWkYPgXth46S/IMvmGYjAaBAID3et4JLnyArlhqruwkA3rWmM2kXnt
rSejOe0HbkGzZtl0T456lrav01ixTu7dgLY1nphskstffC9qHZCAqUzOBE5mG6W8DCC3dOpr0Bs0
kJm3L46BjjTXg7G3+fRsJAESDoEqLMqqJZ/ynLlDmqZhqGEZtuUJGU0vnwuIQzQk5OsCXwHxQrot
5Ph4i5dhXHtsX6sOkVvAAylT+LD498dp6huDBfp8CH62BXSlAaWRRPu/whT873b/easVU3ZbiqWs
ATuMevdmVfUXzqvqnZBfNHqjvPC2Z0Rq5FeZBmj0Rv91xRpcIYsJwT+T0vwws4wwsN7sWSW6a0Ev
h8Gyp89DR0THMXwUktwdeKz8y4hcIUT/hTQKX7Id9esD0bySAngwRWKow1ic3bWxjSDlL2p5RVZf
g5PdAosWlljmDYgFnHHdobJf7Esfjp5TjdkOnELBh0EfYFAXVzxvKsXTnbrOpsuhswcBNzvZeFyT
bCbThwKxGlM+uLazh4Um6gs78gw3jhtsJp9GY/tL5tA04knEFnt4KMsla9xDII+qb4UnJ1ZHI39T
L9sVxy7lFpKrtl8Wb0LeiuZcrzWY396iJKkXrFLP34F/m9yhapKd8jdHoLq6vmSvzUDcQytDrfy2
g2r1BZAKM9Op2Ywqocpm0f2Qbt3f5RJ7xz4871DJmyay6Kr88LvDh3v81mZOBHPTFQnZXgUgDKG4
UtL9thE387JFLMYaTyKiTNo3Vw1lJ/8DTMZDkO9kJbOBhVKWgC5T/wekKlAhpnIuaDarsy9HyBkJ
7CRC0RdKeh2rrUWnvwFRE9tfbi7uuJG9zFJ6CQ9XPbTcQTUNjqFJ4hwya7ZUGbhCRCxIkv1ENUyC
g4tJdBE1xj2EikE0US4KoFMQMAOcYTEoJqn8FbvHJhahVFv07Vovm49WhbKgizT7vKGl/VmdlNCV
WDn7DkrK0LnFMsKEXG4DLDuF30BJ3Al9ZdXlid6UkLNiizuuzIx35IU6Jzk48Yne8kmbaQnjFV/R
Z11ED8MWeadfsz35z/1IBctjbhCrC+B0VWNkhxIf/6ALIiHlkSCcGr/EUgQabkPl6KBN/1XPHJ6s
0UVjl4SCx98vYM/gFvvibSip+gOV+9YNBDNIL/vAkQrZE5o3om3Do/ogwK9+/GPF8qeLaEbLEBx0
qTGT3ujQyVd86gG2/a+/15TExnZuypA2754535r/LKgwwxIpIbmfC58+jDeDGFat8+vn3BuHKDIw
uyHuDPXPj1FQpz6qgyxQX9tPRJUWwNp8VvDu+FvMr+L4zus7r6vP6O9sRuSjf4Mrlql9u10/X4fM
8of+5Sn7sPHM2pl440nbFeVlru8NEeA3K6SsFULPZV+vF5PQIDyBBrPCC8hwA41/2q54GhCHim8X
0nyHPdTUbCzzwBgnOO4nYum8mmpsoOx7FyB9dZrwTn03zKzBhBMaYhK/x81SCzLIPFfO0Xa2u9s3
ZHzC5E6uen/WnVzOFvNp4EY8LSrFtgUrowZ39bbjA8WEviUFFaKgA1RSkls18sNdSGm4DIjcOZht
l6X/TLhYnzeGazZHhWRbrRkXefIsqHkHqbu4DoaWCeBxDx7mqCCP2TNuI+HY0Uc0N4QRTuDvBCIi
eXFMXUkk/J64Jzo4o8qO8WDdPLhLEvW9nYw60IbxCqgDRJ/gSCdzZiPPCb/z3uEC5yei5h6WFzs1
sw/fSZtVGu6yT4XKkdBnGDjuqFFCguS5x24WftZzaxeF/Gx3CKBfLlNtwNEhmdZo0+mXhfdRnGnt
15oqyJdaG/f95bLc1gHTwtBS7XVqohxjdDT4xfzpr6gli0pC4G+S1rXrBygsfU5Rr51XV41a2i/H
PO74W3FowtKW4z2lqGwC9mO/KYKn5BbC73XTIupVZJG8fFRMcRD3RL3RK8m6bPBtJYjeQ22HfZNJ
1AvCp1g5TZxpfqa7BOEg3jVi4esBNn2NIBFf3i9sPG4Huturwx+f+kQn0KMg717yUIsTydzsMfFc
HNNctivnuHtFxwlve//XIay4ybI+GCTqj1t7RuMu0Ouf5a+4bE+g0aMzzn3EmtpT7tqvBZmodXDI
NMjkklcS+6SyeXXGqmW9VxoXtgbkZQiNZxWjGYCtjnJKQmZ3EXk1SEjpkoOjyA8WHr+nuti3xzmM
zmVA4xwKdsljcCRY6F61lNwJd2CkAxIrrZb/TggbxSoJh3R+vpsdvx3zlU8Oijyc/NdxWY/etJ/g
nHB5M1JRXt1Ye/vJ7SqQV32z8jRShO94gHpiKSzQ07tNaen5pFZ6OVJBqLUEJo1scSxhbyK8a3BJ
VS7gio/+PYE55cf5AOhd/8AF+jRIyuq9vwDMxIPxK28w02ijnWScNIngbchqLTC40u5f15xWNuOB
Zbi57nb+SfpkH1BkB/QBQOgf9JWQIWVAp/DRzEfD4i3qScEaVzZ+v46Xsjv1jRyNS3V4qoRTZ3Ev
tqNMHgtZ3UsjPx0D5fbbHHo0mtWyoc8eniURMTGtZUZLU8lAODMWGEyTrvKMOFQvXpjjyasJd5dI
MYDE9/Snd1uP1dLR8Bm3HdD44GsDvvagATHsNmm/HYpUiT9N9edybLjJgrDUQFprCcbwRbVO2HS/
/yrEuXRYlReFrn5GNEJqC8RTftBKXFK3p8MP5ON6Sj5IMgLTwZBey4iFsDQtGWOAjke1G1MQluA3
lzK/lvVJRR9xoImv7lWi0sSJHsQjJmS1mqC91UXmQpqD8iPYlr5/J2i8fiXkrf1MrPtbUzb+SOHL
s2zQDQezWadu1nvBcSowY/gfW8WzDoVJspuBbAJRbcomZLbgaQmpoE0+wVT1hDdZAML3RzqtCfH4
+9/OJF3wEHRMLUncehfucopxQK2Uzgqt1EHm7sQIBrxYoApqrOsUDzlz/TaMrUR1lIUK5wtwrMJR
HCdD05V9GKdKwaHCD98lvdzlDbhy8VKhcH3/O6PLmA2w7pPqHRGDXHVpCSano1t+tPnDgq9z3uvP
T9lxiEbbFdwK+QLBb7WaKKjycU9eYY+Sn/Jrmm6W5CTR6A2cDHrDuMAbS+tHSxw4Pz9hk+68Yyrt
1xZwDRBVR8qovnVAWh2zddcir7zS3Sa+Ns1wVnQ0vz6ZWfAKn4ERnVfjXUYztnxevLWAyP9IZdsP
xJUh2j/Y1nfjxx0Oa9+a2ydcmq1rcu5fOpzfAzC+OUfPT1GTFVaEegxtrV88xpUt5Fzsg0JtAW5Z
s9oTKBFX6SFGCB6dFcrTt81OXKEVz9u9xNfzlK5R4L1Q9yJzbOiujAndjghhpgr9mWi+CtYcsqR4
JIdZWDB4LfagsAN9ig1h5D1nMUuYIqlsYlOO8K0m8HYaoatgek5zxBz5m7DLrxTGH19PsF2bg3Wv
W7RSzLxlUQgw34wIgwBaamxrkWlzralBmsF3hcHOZUnxwTSS2JkhsZ3Qt+UuEICFi3mKhm/Hqz4v
Hs2qFR9Uys/UeBctKhSh7PiXkkuDWwf3zSeJzuRRRiyGN8GDXREttG1XxIOPHHVsy3yXJxRYUnbZ
Ho7xGFK4RvFmRp1hGvEOBNN+taV3wOsgzPLuhlqjhG8g2XJgXpUUCR3397X0nRMk1YH6u9KT+5FW
mBxr8uY3pRJab33fiI1WzJp4v2F+U6oMUwgZsPNeslaDaZowaCe75wicy6sOqisec1dHqjk66zrs
M/Rrc9EIiFt5xkIyeUaWy2XYFmpJwNWIOhVba9Xj17eHHSGd/DiHzGcEzGfdoLSmD/e5aSn1tSZI
kxVoOJqA5q92Eevoh2Uv7lpkVS0uWUD5vb9RyPBNsig4zOzCmFvLxAQEfmmu87/KBeEofqqH1Lfv
GACNR6gLSepiahPC7v4EO0tinM+ZaJWzbwiT9UJjfomw+C0ACw6RJjBo3iA2vPgXoaJKmZzqqMRi
PheOOsI7wJl6p/Qbj5TE88hsMW77zaSCL3NrHLQJxZYJ0gz5XTCw2Nl4R4JibCzUgJT1Ipmq9okL
Os98gdmtUMZGGzJ/3XII1Hrt6bc1+lMzFHYS/5xo7gmr+bHcsbM1BmCmF+yjt8H6KYHRURU41Ng/
s3CsRa6yeuxbtJjdtb+lTF77NbeyD0v41tHSNvGpFozptJCJpkYD/ojEBCkbld0oH80znYHWWre7
lks32xyvQnLY7AO5i+jReBQWbxaze7nWSajFM9FWj3MGBfUNhkoUFVswO//lUnw5Z5yqfs/+DXpb
3C12QcthXsKQpqXBo8y4l114xA8+hUdaXKtK0JREjlboU2QOyCCe8z8VwTqQWWvDLlgpuOwmhRGx
lnyOCAP2pexAil1xWqwRFNbPzWUy5c5EtqRtl4wrVF89nRRczmr5DDOwSbaA2IGQkSW3eMZBNpyh
ruf5BwCQzCqpLTFWsrd3bIWf9gz2JvDPP5HOs+/xuYNxElDI2RPWgbnCljcrIKkJ96iKNdIuFD+0
+iZrVRhqD1BY4HjlCaEYrcqBTRLWjjftYNrlsE+dDt0h71boq5jRjQx2lB5iJ8jGe9lA4YdQ+ZXf
QKr7qEYGQmrNwDlFNF5AyQ79PVutxa/F3fcuaThdcYdnBtQcBNVX6nn7bmMwgggdtvd2TXodD5cm
JjnYFGu7JDbg8t1+4+xyJQO6FP7Oxg/xZJGKwKuI7eSytQgVmoQSs4kMUJaAyYCMaK+HaUToMCcB
maIik0J37DkFOQY3/EYgb6/VqCyFwTnbYZQLVCuJFb0PvumHO5qJtiYz/XG03+ir62Eh6cGu4btE
0xjbu7QCYnoWwRgi72CTp5ukB0aMuf5Dn0pqw94GxWYZeVPKNggSDBeMKaR8KZogQkNy/qi0+7dx
mfHXCKAEcFHvDJbQccscFy9Nl68cfXnoosAu1ri55l2kyBBxwLaRC0QFN24QV1J+ORulUOsz27+w
WhY/GYepqQlAveyCqa8sH+m/1Ud9yOCFYtX+7Eo5QNM2qD7zJMQV97U5AvZ5tZw79/ethetBlrcm
ed6aFiqPbPL2QRaH9kfcPuV6ZoA88LDizmTzUF1Zid+OQRLpVYyEjLwQ9AKDq0keJQ0J/+7u8aey
RtVOCj2FXKML+VicOJt+6HaiqEYT4ZzOhkBY4dO85bKg4bz8GhxRipWprhERfHzGxsnxeRDu96Hm
8idhw8ucTXJdE4rGFKZKvcnl5I2R2wCiyCT68lJ3+KT2ZUM/FB/EUjSjiej3axqDi/9VNDu6TjQm
W8pni5YsamrI7j/7ENripr/F1mt5oC26vNju1qwqOOQBTyNpZMK3c7q15bs4/M5gACmTmJGQMcpO
FpzWCBEaH0gkwHcsTjXaG5QU5KJCfHwf0oJ01/sczY7Fk14YA9P8rl91Lji2ovAoHDDDyBGrPUAd
qJRfVbBAc7fyftMTB9fVc1hfc7JmU3cfk4vrXmQ6JzzzxQit6I6L+Xy6HZUqSMZnY/E5t0KhOGD6
JHv2XDL64EGlJm0pMqu3QuLtQn2iCfcG42+SLfhTz7T3MzJvwovBKEo3OOemuVYy9bCeACZvjIp0
0idVCevYCYlNvp83bZgRjloZPkyzw3qng/AIbCaRq/TjiiZUuDOfLh6bAxM77KvEpGxYNL0/eYsw
o3uXv5+6DcI6m5XvPfDHsLV9YqEwCz03W1FQqg5dO5DkvCIO1FQFIdpkkKR86vKvWvBV9anoPdtt
gwX0FyMrIRNkYNofQHRhzFvJsLcE/JlIi5jX4Yae46YjrKcGFD8km6S9occfgmUJqsfsN5S/dZkj
CjWsjlR7QvOEdu4hTCRjqa3nXQdxDjdTGKITknDX0xcXSRB9gFmk+7/CSXrE0Jh46kmnRVsJ8eWN
MSrQ9zcrnDmZ8NqWwaENBZTknWtPpMbWPI2i/dxBkDHyryYucO0WJhz6ONK9EYL2xZahtQZjTkll
z4GkUOQzl9Kb1lfKuF0Q9OT3rdzIpCNjnSt4SWcsinu0tBXzo7+Nb7QcGOhDjQCypP/DvZdCQIlz
yX0D/w36UC8tYCALOxtTsQ5xkZrUZKfiU1fn16QiidvAWE2YTHzm22rye6NZKzXxXXJsXJE9o/5e
QuN8qXuQTPNZC/FQfXPGUFBhPF7z+V9di/cc7og8vf51GLx593CmIT6pqQWTW32UbkpiBDQ1cJ/Z
P7UxS+Ved11r7u8xSreAzf9rcMyU8qXTHoYRgaE485Dv5Qc5b3dKh+ZcmnJIqqXU4V+bbXHNEUl6
wN7Jf24iKCckLwiEQydidz1WEECsc1iZcyEYRqLgIxDQnt/FI85A6Ht/ttlGMBajiv5IKvhJigrD
y3PttMahniu2KEOhQq4l1rwYdOPuZW34ZP94fmMaWr+897gdrkftHEog1WD7AY4Nqbu9xYL/TlpO
Pp+U9yMlup9zEqEZ8xwQ0O8JTCT1f0Ly/wCcNmnaF78BQAIEyUhyZPYkv/l8gHok8Ez1agLLep0g
S6ca9LT+LS5Un/darYbxJlV/anvovUD4M9rV5Dt+Rrwk5xPxd5icDw6fy1sPpUaKkT0mBbnlTatk
Y+R0+jiwv+9qAV++aasiSGStZbXloUJRgGf3XpWfSmEsBAtOsEODOmJhp5vU+v4EGD7rN5Hcom6h
XM9QnAumG14tFJMh9b6MH3/rkf6adXtPUgARm9JCU+hVCGmVk6pT2vVVqaZLh5kXT/yfo1Rm+6qK
jHHe9A0EH0/MQbJZ5lYYBlqmZQM63sq3n/8R5233Bt4CYyUS9LtGmMT2SwAE4kTCEcn+k2U12k8m
WUod40za/MAZndk/Dws7OIIzXuurwWu+JORH4Q99bNr97TJCUFfIAJBui8Ae2Bou+K/EXP6dIWtS
UJKmeyXFcldS/goxyEB9k4wiQjiS/ksuVsmPHb7EnJR/QvPsH0WoTPyAMkzylGvGJitDcxTqUG2S
Y3ID3cAwDZPFPnzT6daVj32LYAxKA829kgnjuNgMxR9XvO9nZwd1aRfKR4xdRCWCEMhuDx5SIl/1
VcZHzpeU2Wtd4k7wuO+CwpRANFRE7ZBfgyXYVaPyc/i603CGYjUPRXB8VL9YsM4uWnHN7Eb/6cH9
aTpHOjIzAMpbG7KUQ5uHWJLGHlPvXQerhI7J2iEVmcpQ3InI2zvJOVOh1tJDLC68Io10IGKHfq4B
3XGdUiPcUkSg4rIKBUTkr3Avn3bapFgft37poRQyVTyQ9S+zisxyi9csAHMMPDfyjMIe3GHY0DYi
uN4ofXCmgmeTAeq279dEjVmVDFQhmnNRua2tExwxcOKoG+h/2jAtLbyGZqbt7cyEvy/ikTlEHvYr
cI81/ybTRYfpfJfUrR5y+IjD63jgJzA6XA3HrC8ovScUh3LXy+hYA0XlakbPwFuQz/IgAvPj++3M
q1suOX5ADCzEufWHT0dWqXpE4jQ/cRekPKPjw4TyLJzcfBldptx+1Fmo3TnoJ5tPYkUv03wDhoXD
NqaRota//eUaibH341X6x+fOqbkHf112wgRCwYvUK2SC7bpxo/fPSR5W6EBssqXAJj/6qoKOZRTv
5sTZhb5Hclvar+qByF8+5f1HMQoMEiamsnUpAgRbf5nOGLvKqci7ZbybYbfQ+UXxZflNKyZ1N985
vl/WNebBAksMNrEOv3NF+J9g+u0agllx6SqcHBx0W8+pd6bAHxSP0D99mjBLvNnkS3IjUs0C9x3H
OS9UCZCW6FAxALCOtorNhMtvoPyUEktpYrxNntRBo6xo7zs+MJDSmgULl2lQ4EgufPNlnx0iyy4V
7x8f+AARSaAWcSgQ+Rdk3eEsLtki+y1mvMtCAqerrqTO2c06EKekp3XLOCE+NSR4aMNS2Us4NOkg
Ms++I12jVmm64RAlVYJRDDMHezB7dAi961d6vrhG5S7WoL8UhFOLYHBl+IrwK0ZI1QROuANOtLwc
4hdjaGha9MvoWp4htGr4p/+I8wfPnRaDM0WZQi2UKKFnUjOvp5idNH5oaPQVNuoTAVAR4guBSsPC
6qYyRH7fz+QJJV2DrN7SF6QVLECkwMSsIi2QdJKcS0McM/KDEiOK3qT3kDtVzChy+1+Qm/N0ufY/
iWay1tBT+6V4Xlb+lDPUKV5HrF5PxX7/zaQvQjZECQtVi5sSEkGE9nA6Zibsv/92Q80evrSe2HZL
VR7bY/Mwym05obpsQW63Ll7CTHPt/0lhS+j4CGOL4pd30i8SBKp2Itn6UbnUfu3kSYQq2cyp4g68
FWZ98fAqxi9sU+fYDqGdtenXdOSBOd2voG9PIkxqO1RFKtLMGg4E6UOJvRw0Av3RRnLSw9on8lRA
pP3GPU40QFq8Cp/ut9xfZaoEHV03F/PmE6iM0+fUNehs3kIThBG6umctQ7l4JlOSBMqt9W9V45qH
/9+5S0unMq6ylePCGHbK1WW/u+3UjUefGxRfTkHwYrCQss4HfMOJEd7J/tSwKvhkSZ2UOsxULq8O
hKlah5EOvlgF3WThuqZtAj1myr/P00GJgrrr/jQBxzleCPqkrLZyZ+vUq9I0Y3UvFKHUIMlBTfXj
OTl9BQtz9fE2toutd2VL0oh4Xn07qBcgVbtUlIYqexG/yh788Cupy35NLxVErVMpM9hSEijfY8Yh
a992GClP8WWgHOLFjjg1gMbF9w6Jo7NrEEwZA7HUR3YXH7TjyElzGNuuZDOlgYA/rK2rW3DoCYCr
joeggjfAvyM6A2MDMgIQTaqwVA0+okpbrZNq+qlHaENawE7O8cUry6wu8GDd1h7Eizf8St3qBmQv
nq6iWBmo7MZUEY2WVC07U+6v9/KWsy82D6qcW5wXEcRqfLKTzvtuu+M/kOBoh6Tjq077+8x7Yewi
afcri3h7hMoh7As31vOJ/PSwXUvy4eW1l7PphP0zdzCJPG+KfoCTf7HJto73FATN/4wHC8PFmrMe
1AVrPdi7T9hLJBFv+4ANl8Itxa+fCHoUv9EJQtZsUrXPCZEwyrNqeGPbPsrpfdIped7Gk0DdGX0h
Pfe+6hiIY99AEGcuzpP9CuLrsVYeCV+sDZZS8j4/NJCkSUemTAGEvPRWfN3+mtRw9mEoqDf+xpGO
SUR4178idPtCwNzJeWfRGKDVnMzn4m2lmLbh2h3iHbmgCUKYgEzHNY3UqafV1AGTvT3R7PqyvBm1
eoPCJUJV0GusJMW8UDVlkb7EC0tWONq/FXBpq7xxeMf2e6fr6HnABslXv4s7EtMI8Js69YcXHHMJ
XATZ3Ui+2DVHWXx9RASQy5lK/k5UQJz+BfSWboVfB1N0hcU7XgOEAwoVd5lKM+6+tVi0CMri46mg
AYh0q2nMbemvZ2rH4a7dDUI+ju6huZysPV5Ujy94ivIHfkYSVFnrJCgXw1riOdmhjImT2n+nWJXJ
MAz2m87TdKIKH8L/6bz0XOF0Od0E5S3tJ1HztuH1NZpxDBVtoO0Pq7lXzv9QW/8N6EnhHgvG6dlV
A3EIbizORACaP7pJBJ4b68OawwFJ/xt1Z4QbU+nLMe6eSZAXSpQxKFZkiH5+7kEIRCxSrXZJ1VJk
5vlMffR2dvjzqmYpp1CRjshquXnSHkQkGqjqC0By+xh/r2ad4pZ1twBuw07yT2ROYNpVPBkN/OWz
my8St7tKyv+hmEnBaC9U01ymKFZ5jygbqTy7eiAo/THGbwBv60kYXVpx1nWWr8XWcWTLBL2zSYhe
OqohQJYKeG1nCqp3PH1iCjqI5AlCIsUpCZpqScWQQgGK5+q94tuUGTNDO5JAMKTL7+W9rPIAQ4xE
3NctTNojEK1jxmfIU9pCNFiafQPHJXa6XfslgOfs4hSGAJ3m0LJ0bqHQaiwC8F+rZJyj9inyc0rn
sBmpH6RyXPHZvasJZb4+knvyAoUFg+JPnskVCD4PEPZ/91Bdze5FVi36mD+0vx4Vs33pD56peO0k
yVUJ0hCKVeNNZLDUQt9NiByLiwl23NIrNBbkA4fNyCkb8RvwYaA6sRPAInLDNWY3zUJ9nJJtryw0
AlLp5ZRLbHYZ2X6t9sQFQi35EtwfKWagJU5KURNOMh6Bq1Ojz2RzIUhNfqFYtj1Zc4aO5pvI1iTK
592Bi5CKuZQkPXOicf9znHXYmykb2Q9U/lxmGU/ogNtHT+swzxQXYtItKB1ymT7Sw2/LJVbgwBYb
nYV4eXKFWwTA7+ZhJ/1siqrtTgsLX4fMex/e4P7UCT1mmAAWMqcBSYZZdFWEfq1AIWfT7C6VczP5
vUTMDVbHQElmkF+L3PixgHVrOnPGB+lmgjYS6raYH1q3vGugnHEHUTOM801Q0V+np+a+2oU1IEQ6
tfUDpamSioe+0j52KqKg6dbdmO8kH15iP/93TWQ3mb/+DG0NAhT9oUCFO368tzKcoYEO46/1R9Lr
F40La5hiA62h/T2B6YDZDR9yinD0lMPwudnPE0P6lTGPN/QKIP3+tI6LFGSZw2x1i4qaOvrRNYLt
+S/TYM3DF0q+nthpX3PDqy5fnjG6T5H0S8mkslX6Mk2jirvmDycA4grgU06CvMLZSBHnjqa7mcLP
6fcCxstrNhuplBjp02oTfp2X3/Yw1wN6GkKT2+YlWWHwzJjqzk1l4Gyojaoy0wfUcsulqllpD0Ku
vnQM65mD9cRpnIF28LK4SLBtmqIvEaKj7jljtRp3m0t1cNBhGTPI53Et6ihWUwtOXVdpask2GR0f
1HAT+1971tBTMNc+x9N76m+ADO4Y6QDwSm0mFFrEFTCA42mawFS4Qm/V4wdiYtZu6TRKC/Wc0x7x
yP6AEi5y35Lq5DswlqYxDpRk/bM77cT9MdT/i7SeMSr26MQPL6DwRuo8BNXsO7tYvH8dfyr28uAx
Upbyx9Eeo4YfNIGwwDs2iixaxUg7JYxQ/Z8nGiCq/84Dwlx22hwu4Ovhpcprzuof3uyeEWw89Lg9
2LQxKgHnfAFAg8/FkrVAEQ/I5//DQ96JCePY1MbmoggaSTXIlfYBUYjqWhU5HdGjUVxaGA55x2AI
uxqmNYldcmHuZ93yU4rEA2DNkmsCVGKh+TSdGaqWFht5eGUnKlyTNEcDlzC9OX7nIPNlVSAiWpQc
AA3+IV7tDIS6pOjGOGglj4c9gmObt6kX3t3i78gKwITZ9jA9aw4x5O+NBhPd2xLa7TRFFGKPt3f8
TvpN/7tsF2V86XioqJCd9rAdMLVieX0gtC6fcuSLjU1Q2+5I7VvzCKCLiNe+Nmu8PRk4l8zYH3dr
7wtEj8OFKV1eMnuezJKzwv80xSjl6JFPBOslDhpuDW1N67O0AGPmvkltspkRf3TGbRXHVayMzdZH
6zpH2v4jbbdmpFBeg7lH7LrkjiuagjoTZCOMfHDEnq02OZB/y5rmdY/vVsccktIGghhsnuy8VQx8
9zA6CmFTTt0WjgReUG5QTLVXEktGhy+5w/tBNfDyPh0CevYE89wqsKiRiuuuFC3N9/TYdFTns2ZX
LzAMuvE0AbziTd8z97ha0ZDx+x2SOU/PDz8H/BTWLo+c9cZDiPZw2kbzKTlVFwSY0ItnUdgBdwp5
kltMZ87rzJAneQvd2zXLKRHFmhbsLyRwpnkBJqaJB2LYxlqv7JVNf6STdC3eQbyQg4GEbDCP5YX1
ouu3JPGeqzztmwfgY2JijuqTXuIIn8u/Md62mZ0cKu22fXGJ0uOKoQRgnalmNX/yJh2MZ3BiXlk/
P99gO1BHb7rZcC68eLaIjaxLc3HyaZuNrOGpVsNxn8nPlBrd0Yl/pPFjjHBnLUMwvyHs759G6lkj
mwwiR9v4kJFUoT7tobnUzszK662osGQ+SgyefZaSVRD8UjbDCg8BNVpr6F1y40+3P10uUjPFZazk
7fg+3yaYaKtXu3UWyjPjKIiQtMV9yyCKaHaCk7TX+W68hKn9k6jEqVA1wLAUXOVVjTnC/PC1nUDt
bBsKLA4EImPMJBE94TIBo4Y4rwNxq3Ixw9mdQAOvIcMXmZ9GYLXrItu6VAObnkAAnd7tY2k8hpOI
BP7oz3IQ9ZvO7RVZCA5yWpm/j//QprsCdiQZedWbJcklgF5XRv9QQU0DG/zEucOziloD7fFQqKoR
ukXihs71SR7Mb/TmOsvtkpSzAnHx/jZ/785HkUEE0U5qoDmsUFJA3AoXxsvW6ju7SlnkEb7YfhFp
fJH9NEDQEyb7FbBX2BoaGJlocs8FkG+WZ6yDjIdLsr7Mu8B3XyMhfEUkL0nrJcjK55cNZccBjjTM
V9giFjmyHbzONhL3CRNOF3pYLyjOKhFXZFXyvl9F2JBESGvRImE2xVBmYbyNs0Ps1Y+YJ8xZEqz+
45mjkUnR104NCqeYW0nxHU1doB4Gw9dv2z86Emc31yvz78PNDFulvKBt4a2tr/H2WxchDiGx0iKi
MamR9pO2EeuTXERsm8pXpiEveDjcoj6EvIdyvIJIpMNEQNqyPnoQdAdKsEDpRnAgRVgeo5j51Jdc
0tHMcJjFuwDxk6lmXw/6Qq3hHirJ/bxB7RJcQo9ULAvMkU2fUcMzVa91/OpCKg7w/APYvCTvIHjW
FYxhCInytUrhk7CXkZ/MqzAS/QnVzWdg0HhrSVG0wiqxnBbPx3jR2Nc528r0Dib9XZEAWDpVOH8O
V812yiGp2PdvKeCdHBEV/VcOVXEE9nBeEvQ4+cshWibOJZJ86Z798SUulGxBv5j5dJwQQJSlfeIe
Exn6dAtPDIts3SVgaH5YzoDjF1IAgYJp4xmCjY/cnP0Nw1DBLbabwHwC/BXQ+X8WSLMApxamdiMx
bucszeHrtb3NTl4ZHafXSCJfpeKtFpBiBB8jXG8EUxwFPri52U1nBdawXpgkO2DIrGTRxMQBXLz2
Ltcy5G+RasnrENqOrk5UBWWGW7WAsg0sh6Tmkwz4So91QVZEi0YFtXXBW2xJ4OxmD+TzDvqhCiZN
/rrUjfj4wM8dgyZdSlXGbBAZTy+Rfr3HMN46ompENz2ggZiKuuqLIErBxbECONqE96Tk1J8mnqMi
JF7u/OEM4N84/+JA3IJ6MX2IcKdM48CWa2FgWTN4OYjVxNu10NaQCznwBpdvOc2cJl/7Qmaohnpl
FowcGST3qUCHfgIKjfblRVWM3SXHFOFUfRdgzgSFhieuaPXJOWL0iBXQfbLsSsYtf3Nt5Sis/A5O
Olne+qR36Vd8gtUt5TpaPt/BACvT9VPyKGmFsqweVPEonbJfdyknrFzUCn/cY3eKOMOXuk1xFuXD
j4mwJDOv/aO+hXVR784XADSrRcKva4mmpBgFN4pPo0hI+qvZ3xBcUT1MxxJNMWeyRjocu7ryeBFz
E/kuyj2oBBlQCXvZDhn9+WNWDGzLGAUKE24RA+A1M6Sr+n94xYCu5ABveflw33nP732s8wQSGIeJ
w8ivSVmSmgpn8qvuqgku4b2kcQ1x3HfrjAteAAc3ZYyoZ/D1BvdP2zFRXskyDELuGgckJZ5MTYi3
5efdwWHzCGW2X9ZwdB5pp5CBcfdh/eRCVmeCWtuuL1jEHyS1HUTWRAbjVP4bvbBWDhrJe0TaHxO0
VWpCPDnQAdmyAkJdxx2NG+rHozTNv0HgRYg4SrSDd+xINIc0Ehfo1iZFJuWTWKVWAZ+pBsFlLP2l
0+GycD2nSlDrWw5IUrxlyqkl/WTHF2nZBdCWVoDHJZZNyK0Eqf72RBJByfPLqI3t+YS7p7/9WtfR
8sM0U3r4r4Hi/5mYF48AsYCo5d2fEY+UyVnCT/ITTbtxHkry+cRfftxv/VCUjcxj5igUfzdLDQN/
SBoz6Q2400fG3y3o3vDdHtz1ar3Shq/iJrmGYetp8xOsDIcITnjK4eO22gp/v+zWbbgS72Kzyqzb
TuTqUBvisG45V0zKOcl8pHOH0Zpvte0KNEAto2iV1CCOFFHsSmhZMuaTB5VFNjHwvwxNsPOGzYNa
DwUZzesFb8THFGNn7wZ1CMRmLvWFEcEBJnzAS7bj9EbPKUYQNrbxi1j8hKjM9M+QQXJkaEegAWqs
IbhPu0KUtvsePGi7MgyAYeu8u9TF/b1qbbfgsZFTaEf5knpq8ARt8oOeW2u51V9Zlqq5sm4iocY3
dOWj1SlQTc3dekLr2Hu6E9dSXeeHOqUlOdyvDClRPpF6HHu8xk9LxkcVWtuFA4PtecJ2HiPC/Wfq
SXLSPGeVtEaZ57NSyGvYNYeSs93u3q4FRCAkYHOd5IeslDpg8RfZ3a0t0sOElHkDdlxl4sZFVIFm
KJRjh/SKM7ILIkW1+vL68jUuf3B1CXHKdowdIYxUZFVFGijt5k42Ousx58tChWB4gysumhDr/zTQ
Y3yPIv10FxOF+jh6EmOkahG4/Q+ABpPY2kiCalpiK0fFGYaeM7cB+GMd8iguQkx+6R50XaT8HCFq
XS+SO1jJN3TS1mkHTQwitXtPZZBDhBlwzn46XjZWAY6LOSXrvmci6NddAwM5ry3L7Wxprt/v3PAd
cPoka4CCFpAEybzU2OAtFE0qTgJYAz9xrIclwpWss4rTd4hmlTf2O98rk6oFP9+wJazq5M2zT3nR
TdUg5MRJHRCVJqocOvN8/8fSDO+UB5eA/2wGsxLHdxTyJSnUPVuXnezCGG9wvuVw2VdrPa3v+4Vx
xUqWqBdgofXMIOlvInpBqMTUFYovBhzuOH/nZLZHVsMUDBEuZP1+JcXRL1eC9hQ/SDI9b+zs1x++
n/deMdYwsWtMZhqKZRYMYMZQtgQKAYiw2RlVgL8b12PExLyp4iPFhqhwxaY2MsLp+NAOUvuQGoEJ
IgJVzocNOEzNXhKifBdGEgAL0+QbE47vvwtJjME0yEb/BebFXhnUVaxztkfvvWgOJF8XyVbrmn2f
H2hGcBd9WslPuyrzPEjcTduLblgbBgcva/Plut1jpOREZ36X6Wj8gzO7SttcKQSUe/mtP6zGbouK
VvGGIqaTC4VxTuS1qgsWzP5VUTm+WJtpkSnI/bICLOn5q95HEv8lpsPd8dI9Nh7xaY2zNDbuOg9b
Hy7p1Ckn0L2qzDPRU0PyHLxKlc8tEaNxyXA8WETm0noDfH8snd+rIVTVFBkzSJitLgiKywshkv83
9qQoGN3SS9hPq/mrcX5na4JPWvFjEpuA0oJUT6JLADlRTo1/3XhrArW2WlIDSQ0gvcNi2CVR0EGa
jDH5f59g7BsiJjq8ewDrfqPWWrkC94h62WAq5xj0fsmEshLGSfZ+nPxUivrca6f8pOLe3HMPEiiI
0R5lQYVXa7ZvGau9LBFOLKfZ3XOXbBk35kyWh7zNw3YOVe/T0bpMwmIxiMt/Czfj4bUol3ZR4g5A
+8ri9fEITofKGvmHV/0mcyW7F/eMwha2rBt6heUeVEUMXuIoT7bZV5d3g0m8yglOR5NSjFnE3TsU
TstzB68PGnEeoFAhNMgT1K2WpMveWljGz80d1HS0RlHPVkzPlZcrG8uOjeJzoqlErg4Yk7V5/X++
FFzM9RpHHbVPm7b9HCVqhMlJgdSzTKN7Nwa9tbOCetJHxXX+zUQ1vYLczW80h26JTO2g/DF2ANVh
HQTLVwdU8x71Y0anpwaEKNzguzfk0DyaK+RN1f6NQgz1oWzZyHIicVksStFU8COkpgZjb7PCfYX7
NAfGtNP7uF4OCS5YPESVDjYpE9bSmuXq/8k2T6EKJsZGZwTJnkJ+MLZMR/33QHxUU25iIbFN+xqY
VkVTW/pgNIEtbo/ndhAPQownY3cxcpGDmD0gXFiMovnouQkRw8uDGWrbzhY4RhQ7as4Nf9jDLLzz
frYC7jblEFs7Kip1Y6HGBKUmVXP+UPtgQ88olU2IMHVpkIAiGf4kY7Jnh6AHIH2paikX3sUhihGI
Ipi59c6vLwi5xcgevXc+vAOk0DCYs6oqVVWjGQtF/XFQo5N25lbDO4lHVky1LYnDv/BjnqJk6KOf
nvxiG0DrT5+D+gdczOsoTDp8t3uRCF0JYSd/IvI8uY+lg4z8vy/ZP49vx7FxCm+pTOeniubWW2Zn
60U79RpVNMTMXZAVrEEeT7Chc/C2OGjc00+SxZ1hKTtHa1dWWPrJ6wr1VUKBJ66GEsn2+0jTQpve
0g+Oedf/tBbn12ZGnFHYPMvre6TX+SVp9Bt8LPCXROVFh12YzWS/aN2Axn7IXwhH6gnZF0f7X24Q
X0rMEqRpfUc7AfPV+C4cebRJ3Z2buCDh/KEMisKYVDoIKpzmXK/nJgOIE+21s6DvEWVz+863AoAU
ftOSychUbKtWsPS+e7n3KMIzwlBMu7bPeqa4UAMuLzi+dfEcu3ZzXJzf4RbE/bVabYIynPDig5qS
kX+RzwgJRwHkniOJSBuyaqMcKIz92ZulCdKCSC5Y9iqrhx4TEf6y67385E3HupC1Y5hmsJIIUyhb
RspxHIUd5IvaP8nLgEqFINa5AA3U25MgznOAwMQ9PsGofPbKQNcNJGJlyK64TQsteF4jrVKvN0hT
dYkH55QNNdf4amqJrkOXYbnU3lKzcrBWYMYGvPQYt8IOYPibiKnyccd5tlYCTjhYs0oOOKHONseV
Pizih2aJEE6pJYPxwFf+HXOzBctEadCP013IsUbyL79Ovi8NPlpy73O5E9kICf2WsIooD/2sr87b
tmuf3o1TcZ3lgqDSp6X+VXrFQqK/xP+2SFXo0/WOdl2wJblHJQiBICq0yLn7j6VYfMeXbAPPD0e3
iGaLP0WokgKiz/JBBsyUvtu4Z8Ye4cOwIVHdXIrHXWKLP8pMoUVRNV2UoeeqthwFtcgj12gfdpMw
tZRywy8DgEYacM9G9jy4oo2loLrbO1DEz6qh69H13VKkPbB6Hu+s6mIFvFfEBRcJR9bMk1zPuznJ
Q4G9bGPGQbibCIVLr7oYBQCGC5GbnCE28gTXgHZgTJJvVu82iaNXZQrvZTO/Sb2FvTV+8DnS2Dfb
cgBM7AKfrufUXM0EKiKQrgK+emqTVugaUSLh3F5cVwZZKh8TdGjl4KnbLUXGQTSZAryxliju6tCD
OVrF0R12j18kU2AV+veRwkYzNeoMrPDSoLehqo/p9m0C4n6xiCyVfDU/qh2jU5SLRcb2ethCp/mP
tkhDqy6b0WzJ/I+YhWN+6uXBIoeBnH9SIuOByKBvXf57EJk82I6yjgR3zgY9KLIZnD+SNdA4NOo6
Is41HUt6Me+GNFZtiZe2A6YAP/O9uMAAl1/4y39744TQYs08nUmZKqP0cQv3RSvR9ogGbFkMrIAu
UZ3tdfNa0w/OvFDyV5a7Pe1iJmNf9KlBSprSuL7AQlTcml8+OgkUi/utNcUnTr4FRjWGaVuCpv95
NatQljS40antC2GnEZ+0NQ3jZ1nYzW2OB14CKCjrvk+levKxnC8CSInKgJm/2rGxOF8pYLPFCRrq
J87VkwQZnx2a1Tf/LiumfgswddPYEBOZuV75I/ml2raBn9dmh+t5Cp9UBDKYGvg6hb2nVykGLrFW
dpzJvjomgUO/zWwE/LEsJCsxvrHMRdptNvdB6YEpGaGqUUMnO+04ZLotxqXS888Kta60tjXU4eIb
EozbJFPwhTMBH3Sea4fu+ZJ76Nc+QnD4OsgWc0xJolyp94yLFI/n5LJxujdasgJW8N4y95Q0AGsq
oxNFPim2Dfahl83P6gURWe6eiVM+CdwvOPA1gAySfI9dwSpyt/OSaLVuNeBqhQD94ncQJE+MR4B6
lq0khOgi7thj3b6UFGAL59C7Js+JNv4HzK3QsIHAmLDrdnjapmh1elvnLIfXcBEH4bNXPh4ShXpd
zmr7/KPUTwcrb3VlyDrwbua0visi8CAeNLnwvzGXnzJ3Mtm49hW0OMJ+O0la39RxGQVxJn5WChdV
6gSE257nC2IY/wl8ROBoBNFbDWx1U/LLQ8F+wer6MaIuV11RYWpSVjSFT8diShQ6wqeolmAgCi8O
cudQyq42MdnxoY8t5u7CYQYIsRyyHbKjR14ChZCPWipa9hQf3zq/FXL0cqpRZ82BRzZI+Dzt9mlP
Y2DFC829RSSt6a/dTHPLJkuL91zzu952Rv0sbuYbt+0vaqwuAtMtoYJX7i9XGb+N4HBbsp+qnyT6
pW6KyZKn1UPQC7h5UV21tEQ3UOFC4sefKuSnuKHP0yCBBZmUc1edFFNj5RI6fGOBvAN3iPxiPNan
PPQNh+kMYHSVJMxYIx9TAsN0DQehEfIkV7D1BJ2u99fxqyIIv8TRBRwfgCRfaq6KpWGJzt8MY/1d
V6xBlJdUomU/VH3ic3q2eZ0jrGPymXELVmEwSlEDT/CPnazME3uxwlRhjQ6yAjAQzI7nM2W96fIz
uNX/re2WGeovuDhUFvZmlsXohbyZkNb+n2c9TUmSxBTNzplDdKUWAM64HE9SmS3rX741W6HdlfB7
LmbXi+lfLr9cLvyudvAbSZHF4NRm1kaMdowYQsxXNRHxxWus626bbL94/7mk2zdcbMBhfjcOjNzM
eP9hFYSbllTR7R+/dQDc+ty4eyu909w7hgSl2Oa1EnIgJLAP2dKz/UEyoT5qgi7lz2h2aPMKcn+j
1yiXpl2gyKaJTS1KJl6+Nl0LQVmNYBEZJRQ3Oer1Yo774Hd1Mudu5fVgTq6j/V5Wt4DL7wfXgPWD
2SQOSi6NqtdfKqHL9/HEeGjbx5GDbqdNZIbYxHHTACqg4t9o9i18RCheUiRnT/Ug4byE0XpCP3hQ
vn542WkRg5K9JM8OGTbDMbI3zPdUyEDbUBvYE3XAnJF+Bqep4cIxe+szHLCVnB9m/ZjsuFTjYjN/
YSLlBrWbyl9ecP95B/tN6qkRgqyLqogn6w/5s6eqTC3Cr4Maz9FbNSFaz/sAfeBLMEMhE5smYOn+
cMYjGcMHBcvEk+hM6CMzZcjJmqcB/rg1yg9hYUzL97FpT/sy/nBAGmrCQekX9gO1GDF/gBIqeX25
pquj1SaEnJM3RR4MX/GaRyj5ZRUtZ3UA9k3xvBL5aIUW0/RD/k77uP6LUTWDHwfnsoqgXaplp12c
t2BOERYJpnMyUMRzkGqJQ4pBicXkxkBG4vY7abJJ+w9rfBqmSd0xdJp7m3tp+QGrnaARi+0vX9R8
eeIa0vYU7UzsSu8aU8SGYfCKikNs35LOJ+WjtLlz8k0dlx6/qku1b+ti3eHzExImlrjmiD/Oof9i
gPkx9LmxNm+ybpb9vdgZdbDItY22yFugRTYp+eBgHXCDMnNufSptj2Xc8FqQZTstvGYiteWaB3am
KH+ogvi8gP81ngMHfiCy+jcHh9apNGmyWPySyLNNVtL8oxWr0G/270SC6LBqaH2fNuqRhgQ3IX8I
Phzo1f87V2Ci7WjOSy1+EEA0nX8bthHI1jq6+ZlIQ2X/jhYJs44Eu7Ri9RHhfVRvErUlNQN13NMY
fBhA8+OO3V5StmNGs2FKs/5mfHuxAk6VJA4EOaEHJg0lL2iYju2L+jE8lK4NlcYMMmmXh2KjsKtt
7I8EZI5yrrOvgOXCHZ2o4nJ68s/pvWp5qrDFmDFP0a+UltV9ZEVdBhFTlOpZCM58baUS9POoZqTb
hu1dFYevKdSj/JfSOflwgyB7pDn8U73J7Z3Frc5rnjO1QBy3lL3UC5FFSRtaTShUKZuZ+pickzT8
VNWvRrp9bWbIosjwrDVwUf+GbqAte20CeUEohDD1XVN87qWe6TuogQaOkQuAlcXa851VrWdeNuXd
brBqQa8lqIcZvZGD+cFj+/iVZ2n8/55f/xnY7KYKRcO0P7hqwU31LtWTdhaPxT4PHwLHXnAf/TA4
a6o0uOnqPOLlxGxGxhFzd5CWCBaB5l7TtKnrPM9Ds5VYyS6oa+Jugj0/UdlnmzEjopeNgJAYS+ty
7XQjyX7se2/1l6mRnbUfNiWJAmAZa6lTqFExzjlxJG32YdnLZMG6w9oCB46z88zYFmzPxAKUilO5
XYHdMSZ+QTc4pGZhp0IhmSazVsd2smFoGz5KDgXTqHx+aICBtHpaDNlJ8ac62zddlF8scwuNRoEV
77ceMy1/gGwFsWnfBhN4aoptJwDPcBR32BDLA9ZaGEBHdnCj9BHfKW5fENoFf67Yu3lDgOpSXlGV
PJWYmOdDGua1DN9KrQWzWbUKwhdczdmIBBnwGXSMt5q3Ae19Kly1nTbrh1jVSCXCseiam6L99Ovc
TKQAtF6ElVvgG3TXK3PRj+Yx02/RAhLp0HsHRD5Y3S8DzTQO29TmQOMNOIRGJTbUXONpGpfaho3e
3oTdm0RcrneP0JALYg4oll3Z/i9cgWtufIGSyJgniRUZCyFs5SjWBvSahcl5NGxDgK4xqTHELEBp
T2gdKIaqqZkRSpbRlNOq0xbapT20bk3xCOysqT9xRM968lMc+mVeCEj8L97CiehRo99SFAG+BrgH
CS6Gc5LYCKHyeMRnLYse/G29wmmJEBpXzh4lOHDYUuo4/JjTHEBu86lFQwuvWh9hqJ1ZGo+z6tj+
v7g9O4CEBwD1SFegqimboiM+dOEM+2GxJ7/azrFpO040D1SzfaxzWDbncIZ5g5bWZWSxrjyiKSf5
/MWTINOZcleY1uxOuSMxMnmoUkDMmnAiXGLQoXkBMnquSShpd3a5DcPdcw2hR3qxjMSl3F62x5lw
v44EGTpVKIVPvgXIOGYeFiZtW63MqgzOnWN68hVKgLIGaIKHOaXtlB+xHJPudv7NBu9w1o0RD3rn
AHi1MAEo0AGUh8ZARUi4RNf2/oJmmwVRgSKnIBZBqKfwflw05HcI2T2NVJ5W8egMiqw2mUz0V6M1
T+KEeAP0K6GgbhjuHqBrP+iVvbqosezViK5d2IE6ALRkcwhaIRxs76pu4ldVFTYIS9Pq5ENCswDi
58U0cjXHiK3kA97fBrltAa2kf8aAY8agFew9vW6Wj4jEX/YeYwLsAqXaIGqeaqmMxZCApFAtwmTP
cSTrLpehS9+MmiYVGb1shAhdGzGz/AduY7G+zo/dsvkw7JeeJrkEkw+pdI7Adme6/+7c8IEnF2U1
tAmzgQQvocgmzPFYIH+o+dZs2nmzY/UaDp24vQhQXOD5IqkD7yfWT8GxgvN2QnqO2Al2XfR0xQHe
Dlk1azmyGZ+QI6rf+v51VpOsVzEguOOFrSggzxwE4c3p0kCULuMX+yeGwAufFuU8kIWuEGp0YlnI
vLk7zzsstPPFfkch2PWqAU/53beLbiSpAjbKmUGY028zoD9skUo6Hepf0a+tFTW8Or6J0qlXz217
jl7qgT62oAQTlgdE/Ln78O92DUQFp9ILzVEipicPvEgMy2Bx8OxY7keuBGitUWYoD52eWiH1IQSB
H8+gyJ9GfVJIx3iF3ABfdBshZnePjSsysO0KgmNRYh1onkElbhrGBTNTTdkN75tT44KdTf9UY+A3
dxDGBgnMSjwWJo74hB5wow7DSYfnneqyfJzR6EcViPy2e/Ya7KUbHTLYncVU0WCE5E0ylKqgsa7l
3wZAix7A7epwzBx8DWO9vbHF+i3prH6UPadE0C55y/CKCGKTjlIc1sFqF9zWWr6cJAEZ6a+Ls5tb
LpmvLay4BVGjPgNGBO9CVEJef+mgm9NK71Usk63LNPeUjbCp3OR+EsBpyI38PvlMCKgb3npe9+ot
fSJhdXD6FhJ7Mv7BIsZf6w2V7O6BBKsM5chNI5WeLOoZbMDQ7xRgTBigxVxkTPwHcecV9uWzHLpb
PU+msPdycndJsk38T+Ds1LGRLEqoy1WwkOJsvo4oGFVEqVpEDxQF6l8/YqrEtdX4dFBnTDsRMGE1
EIW07fH6IJzNoyEEoZqHydswYP/nOenJA2wxHVO+fOcaP10Mh/zzRLJYRI6Pq5HjkeCseqyz9DLa
2mOL5pYzp4u6AIK8UcRThFyvAjdBMXN4lX/gAA5oswgJbWopAqqsxXAwGwQ1xr2tTo/UrhR99UgV
GIq2qC4L6XHw5pogWyzgaArtE0TZnRJInayvfvcxXDAyV+lqNLAm2QT83Tznbcb1sKKVTTj6Tol5
q6F/FOL1uBnj8mnS+zikeuAH/DdTuJdKPW4rg3MzHYZ2DKVrwZKaDV0zH4Dq6E/yJjy6BebfVEd5
/EoDKhFPNqdECGbWZ2gtai3w53s0/M2GuX1qOrn1hIVCryZgOtiWMdVJbKW5367osy6lxaCvWkPH
hi72LCgKClZDNMBmqLcV4MH3HTDFoz0Mh1WgiBZQ1Ke+ywMRRHdFusvz6JSR2wihdUs9J0IKomqC
6AfkCcqd5cjF5gijRNTUSFtOnSBHyebSq3lUINSvascKqMFwcXxJMeNyUpirpV3mEZpSbyImQzGA
b1ab000v0hxLp57fZBW2XONoh8eXoOyZnqRDv7f4ubU7M+3ANHPegA5O+fq+Y9W1zVrDrKfWavQT
6EK5Z4fLJn0rUG2lfGtwgvQOCAOOkitVJQ0yut9xWZN5ZizmtYBfWSkIjIN25TaoE6jFt2vSVlMr
kIsw8k0oJg4valVXTCqk9ttrXL0ST7iNs6gQe3DzSoop5TLpK8sVoDFSWJvPKrKahXkfg7DY2bIG
ZMRE5GJ0Z2U5GY0d0KOaVVHGnytudrYwaTpWp5nFQiR18A5f0N7cb+YDQQzEU4uwT2Y2oojbQnMl
tCTwMtF3ppZYa06Rvn8m1+1iQ79U+7I9PbJMWzOsklEw1djO+TF0VnqnJj9khUZwdJF2ktPRhKdo
myoUqzQtKVlyR/jTC29gGklLnP9j/eo7sB6A4BRFbx0xj5tlhgLGxCvEgp5PE9eUSEqYg6ZVu+TK
REQ8jHpAj3/rtfBEmP8rJg+0i7EF6+QiItVqBHxs0WBYWuNBaMMKA8M0nHrvYjEr8Jy7paZ6gXAp
LjWG0REAHQfLO9IvNLvLYkpEnfN2+0Q2ub3MwBC1UA19BhvBFqt8uThSElUXYe2Xiw/TtB5tDu29
HVdcWP5VtLFQwHprYz/LJQYa5oS+lW3zu5tBLB2gF3NBbd4SR1XdeEVhBPxU6WiEPceiUWZuYeQ6
XsNtgzs0X4D9Ds2/ujKlK/Dhdl8t2gsoqacOlWqf9BhPEyEZDIFfwfiUoYk8Nctr0joEqIOJExTP
NIfn4wUWj0VX+m21jdU35Pk4N804++V5mMrz0ExnHJS9tUQSV1LMQpq9HJ69Qy/QbOr8IOSHPIPA
R47mAq2ZEJDIFPqDUXgl4/UWSWCqpWe79DeV4hS+FYhb0DvOipI2qSkrN51baNYJpQzpEPEBTsZ7
wl85LPhB2bz/b5tdK6HuoUQvfJIlIy6fVaN3j7B/U4wsLsE1zC32Em1LY9TD6eK/lh8sQI+kpbuw
Or8Cq8QgrloJTQG0fHYcnEBCiyG82XcKHcPdMYjWvPKyN4BV8hsCeLfD7koVkHLt1VrDYoTUysdl
MFS1ppax4Gi1zZ1hCyKsqOqTMaQSXo36karx4+FeqKL3Ho9QankyZNFm3eRTDsLKDq0eFIJr/edR
WubR6gPzX6MEjP/BJyz5G3cezWZ1L20vfLicYvz7A6SBriKOZXRrecc45l80/18wpyfotgArIanB
ixuYLIgdFmoAvGfxXkp0mgae2eN1Zv2yF7BNYs8Xz1OoyElRKe4n9XjG7wT4sp6Rrs+fXbQhl4n9
0o1Q3UzKV1VnF02QGIdTmL+SDHmGkZz9JfVMJ4HQkHou2iIRBg9a+KG2xp7mVNM1JasKRKyhMWrG
GeHzkp7b3qZDygzKtsN7L6/kpHw87AWk9Rqnl5ovNwV8mMEFGtqP4AduUJF9Z7IsuxnWHlgqZyoX
uOalt64sTVtov5Puo8dW2QUyL5z+JVjeO9JOsCnbspO5hoP5nTFJPY4w/QmZ5CLETlTKIJF6aeIj
XKFL1lddhIOSssmS68NeacBmBw3IYhGUbjlXXBtvlyzxMV0GNQIEqP5pZbJeorNzFcs2Qy73SRoA
jqPkpoyTyytCyNxfCR4ZyecSumUEa4stf+0mUlyo3aTpdN7SPC70B8tcJ/5uVzsVFcNUuodbKQZO
zCcaDwrUa53JD2+gczOOCce6vU+CY7nV3LlKlzNZIX6XIKaZ1K48LmhJtsuK1qF0lddNwIAo809g
yg/65h7IHjNzVCEJpszUKidmUcTwMxMXAgQ3iQbD+uDo9d+pODngdEn/AWmb5D4NAsQmcf7AfmGP
bVkeVEPNNp09mMnZfOV0gG7YpBKGQsVv8L6e7Pykc5ZnaeAqVhJimlviyUm42igXFknqBNZrHtCI
XUsWRQEG1LNOPGv0ImzhL7IcTj1DR8P6Xs0CkP2C86opmA7hhKDZrr1nX9Q4KfXoUX4SMsOR5a/h
rb/k5Rb/qUW1LGWfP57zIJGzzWWgQtEzlrXvAGM46tJHmhCHJGtqxC9HwGjVXZ2OHJ3mupx0EHq5
F6PVlDwjbMsQdm8vhNqMM+PamhHPpfxqJl/SgqDMs6V5yHq9cqb3iVcJKOxnDoCPZd1hExX6qy66
jUwBgmYg6TRD3UwrG+yGZEvTPVHPN7g3EjGdlx/nc7HIva4eEHJA7XVubz/OukcvGCyeLoZRineG
ReUc34J4J0IN+TsOnwk0kjLdduu7JO+ebGaBd4Awa+D2QSRl0d49UAgmF3YcCyj/CMdmj8jDr4qx
0ojM+zpSARxbSnIugnlWW1NT0iGk2oVEXUOtSHXGD2bUspY5axiQW5dqml/dyZ3/ChTrL009zIJL
RuZ2kA+3NZNlge4PUvB641t30F0p7AKoHloGS7BYNvZEKiD5bHL7qTMO7CUVMe5LnVOOXJDGJR/B
fOacduW/nXMYiijE647VM4xqWCsy7JoH4B4TORmxwhoh8u17C8d7eKqU7ZCPFaRuenQzUmz5+4pw
l3BQQ9+TlpClXAQE39Vn7PHNuzSuhUDeUTiooH3dHYCBnBio3cucB5RdI+y17GlX3t20komSntHK
UmEqhLwBBQrjusa4Yl8IvwW4dKkwX7NmEJfiueIeBYv4XOmYsnRpJtt+89ppBFdigW+Cr0x0Jqp0
Meu8GQ2LuKK5bGdgAHZVfaGZj6SHhdUchh4kJb8whDJ6p9Mog2EZr0SVuPWC5mxV37D4iQZxFBI6
b2obZsMAzwaR1sMJzdYLCoFVnItu4j49MR655TCaAxwxho++QmqAwLat6d4B8fYrjGI2HJ7ixHky
FHOP2P7Noz5IuMR2uJF7a6FVizEDwF5Wn8LvaX2S1fSqpwMmR3CTvMa0msKSA9fXS5+3qgxWZG2x
sSScTFanPyhuGCDp3qJkpfEOCbSh6XmAiw/Xw1pKKGWym1vuE8QB8JWIK+ke0qu4wWHqDKrISyAF
xj2FzVxN51NajuJ1ODSL9ZPuML7ite1naz/rzwW7XzaY8Glkefz0X969ig3gnocgicddpLWHet7V
MDSyULR3GUmYO/SR9DOgL3cuN3WQ/CBE5RIsc/chvXgb0LGuQZLlcUq8a7L4JK6+IIGIJxaN9kqb
nhfj6LfZ6KiZK8Xf5V4mWVgLpPBZ/VDSNePzX+vBMpixCgmoBKQegVYOtEnNHj39WIWQ5ms3385B
xMXtYszdJHsYkEOpxCkvT5Rwnda/kyUlEI5XGVilglmFuSn+iE7ma3hN61h8TDD5LSOtLX2AHbzI
00ZkL3PgCdiKGi3gi66gWfdlMtgorW0+vljpCIOLf3BGAOA413gs2RKwmiLjX5QPROOnPUWEKNPR
CKy0fbuHzHifpDJiX11HvRCaHNthFhLtOJCYPvXU29T71l3MtLPcMXqPR0bRPmCcxuKgpIwo8mB+
saVPan9zB90rAECxq7EvS21TwNPs4ukk1Jni19/G3ZtcnjA6An/RmnQr4X0hEFDRNdBVeiJNUvhA
LfD/YBdLoo74zH9N+7LDKC/0U5FMKYffFTEg+6BlpXXYEs5j6aBrhWEUjEy7olwkUKCrpUuUs9+V
YUaTL1h0Mhv4YETlSnfAem4T42uV+ZvEAl+QJouiqYNktrggL3zg/ZtII/+UaKTykpbhotR/GZJo
nT27FLnMS7rAe7uqOtnQFIliIxO3U0k/WdEf+K5HSzAResORFOxcFFOSXuFb7+CbqHRixhQqpiGy
/gKXQZXz82sFORQXqqWyftOCdV6L7aiCVZLg1jjnN15QsCQHHczsC3rXf96oBMHCMjgiJbqyUrrM
bTFVRfBMWVG92FrDwtcC9d4RXw5aW8AGng0b0QdgX5CkWWfJEAjNXpA0EBCV4OpERzo6pjeuU54j
HxZCu0La7574IGXVst+GuHOeIR2ka2hnYVeYmRJZdudZJbe1qDgEoirtV/tjEAviQ6kEl6hZ2c+z
/N+gEvanEXpCsAaWjWZY7yIAouZPaYTERsJSqerbzIF2qa59HXdHDmQ9KaoaPDGpp/RghairehUV
KrjH0M8sucrDI9vWpJFP29TbNkuHYoiJPBe4CYnKDEwoUm3oKQY2Dvwi/GHV9BtA6mOZWuMMmXCI
MYmQ0tSlKOlXH88CrxakK9JeyeREIbbjqS8ElxpHBv4barqWkLxBC2j77BORStUvmcEEB98QHlYR
SYAXDt4/DuMl1MgH9Cbpz4k+HMyW4CYmYFlytCu2veGh9THet+O7hek1QTYqxC1LC2bEpNnPP/W2
n2DT+an1B/MSt/9UlSiPM18DODHURqoumATdgmFfMnEt899dnbCPk4ISNWGYA4TDz79BtVDNga4D
lD0QxNz9aCWq5l+S5EUN4aZRbHafXongba38NY1Pv+uuoeQ5Uxg8cK8jjuceoF30GtGC6v/QZB98
HuROYQ9Xlae3Rf7/2skgDDk9w9O0dc+5bYoQOw2a3y9tt1DyHNE0e5rSp/s/9vSEvDrRICjHxOI9
0agAe8TA36IrgAMBcXW9rqhvsOyk1zfVC54xtfPW9U/pvl9hiAjiKRJDBTCDp+Lg5acbn0+cAA4N
leh6wohcchoxUELOzk7KBgFsJ+RVKwKsVABJWx8R/A9L+G6XLEIYhh0fcGC00t8FAStZ2Qv92bPB
0+zraho0T8qSO6KyBuStkBsUQgmBw+WH45Espqi4IvcCyn9LsbfNAiOol8dvAZNYvnX8NN6dF/WZ
4p7hH9f2yBhhBb55Vx/CTy21Esd5aoAtCziisxCtFfhPbda+bn1rOVHD6/XGmmAM0cWmFFCNXvZK
aJJm6B0NJ6u4C9hAFA9vpL1mDk75GJQ1POsxncbSLz3ZJexDCJZmMC9vSqHNkjwObLt8mD0LynmI
JwRzL/YwMq1QIWgyE6kMaLKVOwNO0Nxrd+BGv/WU6g4YKMpoPLGtpajrLUceniFhMGFTAugTuZb9
QLMW20j/x8E6wOKd9o40ZBwlrAtGBKr0++ez9ikQIaZplvK3796MnNXCFw2yxNfarp9oYQgaCZre
EcQBKZhuZMGKCFiAQ0b+nbDhe4k2G7PbmFS6pdTIzC7flp4jDfzYjx/8zIUfY4PhXy+SkgJJrYfH
CUWp/9BK0LJQZprkcenDk2rVfGZwYitTyifK/nc32I22N8gqgf0s0VAekwSHbjbpQZz67EBaYVnO
a4IvzgXpPIxWMe6Q/BVvTNeie7FM40y0Vaax3FnqLdrl4LKGRxy71ejIz/RFawG4+9Q2x04wS1wk
9qKnGiKyJhtiHPh1SB1MkrSqebiWp9+jbw5ax0lyC4x8Rf3Gd4svivi/8C7EwfjVpqAGd5GAm5R9
75Yg9gxqbw3WB9A7oqpePTHI6lUmKM8zHeOe9swKvHA3EPBdejdtA+EUN621CedDoL6RQ6VZ5x/R
AVSoUk2EcAjLxssAWRgcEZHQZ6erlqbp31AVhKPvpd+KxG31F/eyCNchCuDRs0Qf+JQbM6Wbsit1
LjamvEmtmEAuljMPuLKjafRHyRBJ+5jA6YLuYZLIweQPBiCFAFrSpZukcquyujPjFcSCpkwPNqIY
5+1OuZMVs5m0VTVVhaBJUXNtTBhxQP8bQny6PgYjhxVYE671HXt2/pVJ2lv/X1LwyuO/drCCuL4u
m02/tNh5u8EZwTHUn7fE09Qqm81CVAYSHr7PJVfpxqbWlMz7o10e31XTcYrliQF5jEfcTxbS+vCv
4BjhBAR4TfzTITzhFP0cJ1Sa9uyu1wO93P2Lno7zZOQSZ9+7HWCHrynBEWJQmEB1SPMoQ2Bcr7JN
A6YPgOoJUzBRfPtzBX7+KDHZcm5JxwMnkD6ukcU81FnNHM8BXe+BFIW0qRngqEtok7jifuGUDFgF
54mjwDBzPoiqmuoDRsw4Bp899EqObf+oSXkyp9vZsvmReJf4NcXmzUMnZSGLQnNZMSqMiKLYA9m2
H4ilQMtXuspxpV2Ud9RVDz1TJJHZZ9IYziHKEUCxlS++ALhbvpiOW+GUFtkv7FmjYXoLbQY7El3k
R9JNPwFUrv8v+qEVuhCbxxqUYKgZ0PzaHR7HZYLJD9D4Ut7h6lFGXOdtAO/xLr0gSZLYS/HKuqR1
UouJ4XonT3iqY7n0VH7UBkxDgDCZGI0bNqvoS9JxeuXAynKwQiTqm6HXyeUQvqABfvDVS7SrD/jv
S+IDnUs9pCs1qL5laDirbwKbHnouxsGjCtgmjKUisJUYRyoT+S2yOmuDOMluBn6Dm2RK90Yn/bzR
tfv+7LXDNgVhbsNhIJm7z03teX2KPJx5DWdqZNPczrRBWHKYESoC18uwAvHN82Rm5E2JL4nGc2r1
76JjgwJCvlGvjjFsBBI4I8kxndmkqhfbIQ78SDxJbSGnkiRR3sjrnvGkPmD0uUfpmBmu/B1okS2y
iGn5k372PY7kbMhs7yByMqqQjz5zJ5+YswySD1G0J0BsuLaVJvJ8KbTTJfFJzTgPmG71nkvQsR9z
UBH6rkPRdkH6p3oCHaXwle2FHXNPNQvpeyxWt801ib1TDRMD575okOdsMYMXWm6wcazj2DcHvbvk
dVP9UDuBa80xRDfUBrA8zyfU3xbMs8l7ndzSjkvbrrPfHrxDWVRP+wJxHTMRWCumHU6MrbeyZ/oW
jEJL7UVOA4tmP8VtQRy+UdyMGG0jc/aRIipYTjf7KG72WMjm9Wx/MK6D/i7u2EGGl6oyJMVFeNTl
VSASULdJHYtzj/amQYpAfNdRC4oBEWtj8Rq9pVdq01v9LQb3d0RBhcGZTQRfND4KElDcA/LjLLpv
itRb0GTrwgmSQb6RUH0sXSu88SN1Q3hCXcM+kN524xot2Xef7tE7U3JUhbAPChtAAmvfsjeRbuWu
cYQHrrUpsPL33TKmoNi+6ovy2mDvY6UstoeEvPbQYxYDMRcJG/KgGKJn2eBwLzxFj7NdwBjYbFDj
+rw3yMHrcQh1AxOoyUwftYn7cphCWilmH+HjDE7qhDkogHsiEICZk8NRJNhRCkz7ySWW49cGX2v5
nkeSvTzhbfxDiIl28hfKfICZT6TOVynAIKT3l2r//UjUWCFcTSVBLegGxejwn4JElmEpBffeQyGa
iwid2QpRzaQS4YjXjCMuGulAigR+yhoagUL6KcynUDLiN5fBpOjhFaoX8zKzn1p+kOiQJh95vpQl
8hvW4O21dSvzc0hLzSsfCKzZz3SZi/3LqbeUD0UWke9PPWL6ji+b5cJ6ACW9u7pCx6Gd8FzAOLKq
ICZkrLfIbDPv6FpqpNQZR9YRLbhaxKiS3l4AsEIOahNH2BsOIiMELmwbhHJLzFtSS+M0KnCMtHhd
c/qtB47Fuhj2jQPKHwUFGcwDf+JcVNbGK8rN78Jq0FoRg8PrVX2zF7FUAQHA30BJSLAxAMGShkG+
Ws4bNj2QQI3rGUNAt7yXtrlKUQF0w86tJuf1zAOinG2ump//j43me4XoYzVdVcB11LIkI3sxtef8
vNGqxK7PRMpMf1vgXvLvOcEa4J00KrHui3mflsfFk7CdsPvlPVehQP5EGkGnsNdQgQecZ6xOw9bN
xArY4WWsqEvV3fPJEBYsWzuBQnsDNn8GrfVfiCtIGxoFnlo6XDQLO+5yAQiEEVubvE5y9bl+q0FG
syRYf/ov7SwAwV01PpPhRkJLY107zMIudhLiD/Z0I72JrkGjBJrP14h6Y73NazC1f6JwxluUOZiE
ObDPiuuyPundTkGsaUvv2OqHzR6GF7z9uGPH4to4Y6hbrEBp0Q5W5m2nhm+5XZw+3VBE+DNq5y9J
LPXYuJnlu0bNppTcCALdtPD/V1HZ6kNTd6Y9vJFlJMyImWsywJ0otUlMNTy6XfLS884nuaOT8eDn
lxWM3sdM3d+QKHSWG318Pw7YPYJIfg3k0RjIseHuCJzDeD+kNSzfXdoPl13EMIccSEBijI1gJ6DJ
wqPYR3kzlSPXb8HtddG0ysYGCjklLu3OqABS6S8h8iUlyDajBR+/J+ZuPLo3LzancfLMR4KzJJcE
bUjI12+ywmVOcrYCvcF89s2UKfKN9YlpiF2NWiMyxQUmYN83ClA+qr8VB6HGW2MmdN5q6QqWyUEh
ZNhmfNWESFhvVix7qbHvN9L9rmsgR410AfZNuGetuYQqA2PkWpjAA2mmJ4WIRyGHwSK3i0Zd6u8O
zl5SWWFLIHtjUk9Zc/Vph/1Y23giz5NkOvLGnBfLwtYDczQaeRJOXcjQHX+iqs87k7+/KBsmh2YJ
C1CnbQQRu6btI0NtFSKf2/UO9FLVNY4dRmn+EZ3VrK6xX5/YvjGGDhb65cTmR2MY7fLQs4RAkNT4
Mp6GRpKMg3bGeQBWgL7Agl5l75jhqjhWDHUHuCvEWFGHfdG6Nv+6pT/GP5913tkUqSLZa2F6VehE
kxbrR+UVuC4MkKG0/q6CsZcEhRxegj2Z/o/zsujAs+oYnPRD1HCFMhAhkZqF3cRKLIcbr/sfSKEh
cj1Cffdv1Hxwt7hc/s29Tburu5vuXZCmkCDVQ9R78xgvdAE+nJCLZyqpx9sieTRw4AB96XBW4CI8
4dQaurm5ecY0Lu6m3jVygcIVhES9vCAmv8Wpzkd0ha0DB13sfu2Nh+lBE1rf4yudtfL8L7CbmCa0
oreE6kDJvHqIHxhiW92+hoFk4cnWori+4vN6+TPoHN3fHMUepy30ML6yXNFdKNj3xutuV/gfoCL7
t9MI1dq0ZEiKEiDAV7NLUCqPavajq2Eyqdl2eA2p3wXT7ESsQbX8mzDkVid9e8Gc4cm20wrWWDRP
rOSpQxx6PW2ryzGXRMam+yRI1m/NymgalFKcgYSTF8uZuY0EV0a9FWk/gQl0dzF2qKo8HPj99+ZZ
dtLOlX8Pbk13wsdclCiKCYjkCFhJbF4xWLZTM3OMv0jg3+xp4kyQI0ZiqDsKDmCnBgfcTj0gL7Y7
7jIEYbWnmWGDd1IUKQH4fLiuRUzZ+z8lzQEzxDFXYgiPtR1YtBLLIFDmbvr8wE7lg/ueA+6VUclV
o1202ddiXaggycggKqfCNtRAkHp4XFICL6KKsuDBT4z6ASHK/YoOc00SFj3WJuvyHpk6iHO7NOZg
TpGfGIAAnkdhdKPqVlzF39vqdYwskxXWaNNG2LeiTeKL/MA8z/2mtGOhDIdZ5mS0GzED53eaCrYw
5XgTGVE/b7uOpvgFrQJeE4PmfeRr5Nx3/8eY1CLghGS4olBAQQoQUzgQmTmbBX9XiV57Nd8TTZPU
APdj6jfuc94OMhhkWY4g8wm5QKzXyHaWOpxGTbboX/gSOzEnUtkwrWfSkYPTG5jHCsamO53zZ48W
Mx9ODVuE3mugCa4ZKa+BkEtUSmaQOIrhkCwv4M5u9veJ5iH9AlE5yYQBfz6Z8htXDnSmJytD/LJG
+KdD1xIc8PiqoSKLSreQAMhHkSuTOTobZl5etNT4IhbYaB1PDRDWdOkroZbzt9aQxYJoDSNNg1hq
Z/4+CHQWr+y4qNhcQSiKvrowBfosuJccl57TuQALe2wWH+7nt1gQ7V8L835dEhNQjOf2UhbmaAiH
FLHpovNNrL4/argJqit/JKv68wbyL1ZpYJP0wfeihYow/aqz/eidoQyikZ7lgZ5O9tqLJjfb1O44
1zS0lGv4M71vShBDXb9nGhZDY5JE8NSQa5k/IlcwF23isk48mhr/8ftY3QbSMhoh5Xr37ZEHRpup
KOP241vY6mzvUhMt3jUbXZ1js39zZRhOiIO4a+yWi7HkM07KHTbhFH2Vh5ifwjhZQyX8lyo+UgZX
mqddIR/eeDwdUPtM2wMirk7LFibk9BPekQ+DghV6jHfb8L34Nv1HFT8aYmfA00UjM9H7RppQKdW9
EL/Acy1Zv2LP6a+gf5SvVLHXBplXTOHuwUNcPvdk3shZUXNzVwcMUDeYYKfhFHeV2bmoljGKEofg
4JNax7wZ+9Xy6lWd2ZV5xwCWA3ehkhOUpgfJoeWWeZ4unqvP+P6coY+hV+vWBBcqa2c7rP3PBcxd
PC2/AvGCSxu92OcknYw8mrOxLJYhiP+Mbf214i1pbkPOstJgoxnj0c6qJeJCw5VfPvdUg36KeLQP
5RgBFbx0MfSEU/XOcr2P58JbvOFmAyu+RqSPvzeRyPlv4JIUByOLMA87PeIeSsiZaJ/vd9wEyYfz
LFL0HebavzsLQjRHkV/+HnN7vc6E4ZPO5DrzYoNWZJWn4yXwOhoKsqmpQzj1uDkXiECOwAjrtUe8
RSfIIAPHgqhNRjAwuHwbKadjRfocGHZTWvpo5hD95b6jwjbkkLaEGJdT8b2LhzfVXgIIkxlhU57N
LDAUAQdWFCg0RIvxI1RS/GBYCjTxjWukouSYteSIg2g54o/PklS0CHaJbmc73KOhibYsfeG8kVXQ
NG9E6yhAcwj5gzzZu1smZX6jhGb/Dnslcv9xlKdOnpQiNqsaQHh4p/qcwcwUFnIRCIqEq6FMttvb
hPeC0rGqlwllB/wtJzXvYkZb1yTHW9byrpQgoPZ09KMAz2pywePJpryvGf7JlIeZa/hBkakjE7lH
SdOckohFFrf2SiPjD9wPQXy6AbauC6ZBNM+AIXP1CShC0pfKRGCV9gRfIcK/nd/n0R/VI+xHK0Gh
LRBrqQPE/hmwmtWXQwiDNcRP2fWfztyuO2rTh6Z3UwUz+9hsia9j5IBh9MKxGaxqFC97pmw2x7cW
WRbEmvUFSvENa59OqAF5T0CI9jm1KdQCti3HBN+/EzE2uubEA0klThN5C06zQZfAFmlwlHirpBS2
S4YL4YaQ4SgbEcAXcUFkmBWQxOSV5Ercl4zDU6fl8Lj1/fH05qBSjEQg41mI52cdfwVCAujRv6vh
jsPrB142Tbj6EK6KJppRaVHmP9KSJ5k/i1KnlGUyVX1n3uZB+pKwwHERA8bmhTWI2/kuhFhpIuvs
fHUIPLK9X3GtVIZR/FNuqR7AGmCam2uJse0ks0WwMR/00CZEadGQXXplQbczZBg4s0qV1ieqUAw6
YVcn300zLmu6PW2I6xx/Q3BglxetSNpMh85If9QjK0sY4EzVeURLl/MAqJHpQlI2of5BRZ2UnE/D
2EoA47i2qTxcBftYVQPew3YlmD9v70VcGjbNdvT2PUdAbbcQoqSB8QBc74iAFcPU7baMZZtgck+4
PmLYfPL2qZRDICJhBfLI5DiaMKndX+idB1TNgReo2SD3nS6dOa7bKST6Yd/TydiBNrnYdmb+6IfA
YjT5GRreS2EtZRqwLasZbe4tCkvLIv072qQzw6MI2i+XKHHXECgwp5oaAvr9UDwE8AP6P4YxHr3x
/XBL7YwLNERIQvCTvq7mxT2gI8Y9aW2QgMcScGs+GFYljn7fvv4MwFjWaigsIUkA44RQFYZinb97
a/NTPgXbQQUYfooc8JnWanmW7g2/H03h99a6sYtro/xYZOx2diEqurAH9OPiRJzidIYzCoG+XmMN
bmXktOceHzmDB7egxtIlKgCLq/8FPr8RVMr7ULlkBoQa7WQoNqawr48dl1LJOeX/yWXYU6bcaMm9
bQz+qWyEF6rj7d7JqO81GSp8huGT7kH5hQMQKbRpJtaZsyfWCxTMbZBqS2fqrn01i9WXr+zHrMla
o/wXcH/qcPi4Mg+MiK56ndSfRkHBv7WkfMgoJOl1EdKFwdcCWib4yJjhRuJPcLEMipLqjN19Ag76
jFP/4bltfVyNeHOSrxaBt0Pgoj5LI1AGIW21Xt7pdzx42SW2F/zYt68RWwyWRbisrONa6s+f1dU5
STRul8c+c5HyB3+/tBwqKMPmJPC1mnqMj2c+SBXlIV9qdEp0bQh7dVSMXN1YmTVhWDtDe7fUk9yS
vcETpmDVdXLh/+iEboDFT7oqrDE6EO7BX2Jatf7KO5fMkQ5SynyzRxuuxvtSgmtvzhvVWGLDM3FZ
mO3OL2dZky66boxzXbiBHWg6ZBA8tqCIy9zhHBOQRS3zw1Yx2sTw5ZrGTO3V9n2C2iNluaQNlmdK
v/83B/2RNxOKDsvzC4jNsl6B4h3xYzbxfBglHn/xz5YlNG+dU1VsRl5Er9HeN20h2MriiUE0Ym9G
5fK/HoIRur21GskMTiqnGxzxsXu328fApb8c0P6AYYOwetAp2/+t4VcAiSnFrU9F33a67o5DdSca
y3qR8nEmnUdhIs2F1PtwQwlvQLTo6ECT2+bgJ6fXAgspvMbg+LvJyjD6Cz4DcNak72ghLaDje+wI
5FYPT3nEJBvfa7QhsZlJySZOeKxihaJNTSyTbPE/JsZYBnZulNcO4/LvwU409+DgwA88tFHOh3lG
wHAKOm7Vsq9L3q8/b2+egUXtyEwPC4mTpP4n1kAnFErWAR1Og0pwn4jO1rCUCeCYFIEGBMY1TDkM
fLt+pgWHxCTUTZJJsu+X560HUne1rEI4Dc3xz1St2biqDY2T2k9MY+gHLXOST0NWD5pJLDQhxipN
iWc+mA/oyVSMfblLPwmzgufFxiciX92DcRdNT185N5Y4Xfy+62fMD/kaPbADTX3e5SAYtT+y2jkO
HfpE0AY5a2F20FKQXbwYE8P836jZ5h1cEeLmXe0pSB4d1jZsYFxv4gseFYebEHg2zVDB0d6By5Bg
HFkM052n4EmDsYYm2/VwjmWjZiTJREnM2gIKpRsc3YH/R3NwyX4kL9y0wthH4cUWuEBjIJMH3Jvz
rSYN2yxY2eZD+MMcALrGd2mxVIdQLx0OLY1KgGnaC/sSv4VeWOktw7Cz/Y0WbOIj9YIg3TAVIOxE
2VxPNK80n/r7zg+d1Wnu3c5WOREm3pMfSn/m1xPK2+pV2OdPgJ89xQY/Gvjnj9/DOgxS0EZNJ3pT
M1EKdiuD9XtDE6hikgPL8S5jAAWlp358qAzGTXCV8s8Rir6rg0XspFCwROrkJcz5BxO0VRMUnvyy
m/TEhw4NPmqai7KG7/56S/FAFAh455niU7hFhoyuJrsjJXX6A4OEpXScBu1xraVohLoEG8IFvdMD
5Sl/xSDNr5I+9lt8pLduBqUT+ur5FiqAFGzCbdbCCgjIqdrl3FW2cwXkbfb3D/RlSRWH8qgUdhXn
feovyp1VSMoA1FEK0jjr+gA/R+M5r3bFFB3Rc0U3q9Nf7k4v2uG/IEDL2gzkwWJl+VqKNPSGCII1
p/tTq2aoHZqxHMJHOWmUaYqWcGlrILY1d8dC4WQUOwhF0GPScr0tdVtPuzArwGPti+ZblzvmWpQF
Q5TpdS25I5heXbEZQXcTzfABl7Tp7c4Ne3oeMkJRRLi5FVoel+5EYaFLWM4jcdC7R2Xyykxb8Nwo
XKF9vqRqICFIGE3jUdu+8UrMYSGSYpSVtpWdIOste8QPwnL0QGZGtehxR7F53QuGcohgtRW/Oqvn
mkZ1+tlqfBif+ZB9/oeENjhWKZfddaT2I+YeUyV2hZv2q7PRocBjCYJHVQv8bUyEPeXWR4j3v9YW
HnMRmq1VuFFRFC2c5VGk5lJieVhgr7YnbVNRoO4Ixoazkhl0JdD5fI8fdYlu9RnGjM0i5oBT+6F5
5cgfYr16Z7r2dPakAvqk9fbpg135+w6CUbmoEvwQQpiyr7FhoHr6nLDomQ1Pgl+3Nity89pu+mJw
37ikBbrLIX5Leh8xa9wZsO0QQ/Sbaazg3ezXppO8d1BE9VqjxALh1NQhiCI/Cswc61EbQRNrsWv6
qbNH+lRAT8zRfNVz60M+VnqOHs5jOD228+mqo8Aj2hbh/yAK41AS33P95qa2WKDJK0AYNcz7PLn1
dPPcqwFh1Q3ZFMSasiq6/62MdpKtD0iEmvWHdua1C+CU6Bkn7vgj5GuyVKKQ27VB3FUWUwjtOM/N
nYzGA4C+fx8gI41iqcdnUc883gSy5HGJ9HMey3OTHGHXsoa0lDz319qSLl5D+L3/k8FYC6HcWGas
ejTrTOHVINhjnHfQ5IluIPHQ26Xc/gxIwFi4gUMPDqgDXnndHLjwjaHG/uSqLYWKsKpboyfNvCs/
t4ayiy+G5cfOODFJwXlGcuph01dgAvcJ8krVS/0H12mXi3OOtoOCPXjfaMQjUCH/GDQ9fNFdPPdv
J7T7qgMqKO+33P68TMvn5vXxWXak/+J0YQoEoAv5RrYdMTT88jNiY5nNmjKx0YaazJWXmOzn/79V
JN8fNHBBwTQFub9rEFtMEvvJMeVWgQ55ldyRbg4pvaJkTshKjyHe0X+f+Ifu1+Y2sEFttaxzwzCZ
4Ltb/cb0qEZCzE8GNNk/MoyDnI71ARvisUhoiaNlqEPXjPz0TtvjJUfXdaxKzjkGO+bBOfARmUvD
AyBVpbd4rUtdZtxjFb7fykIjmbccEERdknmfTZeqF14kMHfvz2dw5ZezvAUDkI5VlLhOsuql/uuf
QURb2Ni62dsIIkL5rgWSBV9Lgg09qGaasa7Wo9dNDD4DKkB9y7UzkPeF7mKtZ/7d4270UEt1CXjE
LhJKnHdoEuRmDzsvJHCjUVvOw3CkwoxX4uVEVbsdR3DpljklY8ctHijf4LN/dhAtnJJweohpAkeo
XKI4TQo/7OaElkF5wVpgCjMVvyKDrdzY2RoNuTUMbiMVvhqFcNzFvyHbYtNG5XPWW1aXxWsjymp6
NBOE3/G4FZV66eib2hHQt1HoiYaeBuEU3PB6zCdk/8HYntQhXARB2oeus0dbe3D5btdNevc4USGh
5jGVYlc1w8rxyxQyfBS5dJYzKAhcf8NX7AZC0aT1As9LVf/SEgdD7WmNJlxpbLUwE27klPrZGlrI
vN0kSshyOZJeYm/51GmOe5wWwdtvC1NW0TmZvv+2+NUS3VRpkatfyJ7nqrB7CXgHU5mOV51+UYIo
e2wepdHTBTtpg8hyQX5TP516QPICadJHyQaUu9BOsbntjSnnhjJzQpf9VdvVwzQXx/ZFIAJiDP0v
MVekuy4IRrpSnyTIk5jDe7XaGKFdwgnAlg/z4DUgtMCIb7g8HDMyM8OOLrKaTIbKXJ5FpYXfYXk0
GIF/EMc4E2gsqp2SWfW+LKDT7tcLUfjGuSor7+4zdJKO0LXyHmFYWgE4lq30kg3Hy5Yzb/Ljkbzr
ZLMQXC5xTMnQnnUKZuoe9v7rmockjvqX4ZlUiXx2vVnE9WD8vnTtcosFefHtcFAICC89PunLb1Sr
a0d5VmH3T7NDrF29aMsJyvt6gGfvJeScVN+zQFT8Y+K0EQq/+aw9eu8QQIUjmJlGByolKg22GvTP
xPGK6ZZwECixPh3Jd3+HfxA4wg0ycu7n9D1RxistNIOwp9xXXHdA+bFuED0Mt3SE7Sq984zCXtt9
7Jkw4nCtp0GudHC6cdwimqfR1PpYmRRJBrR6kohmgv/LaTdDlkmHZ4NUYKoQH1BQSJiRvgy5XLlw
o9NzKaWba4oV2DgGOYtz1lC6CGn7Ama16dBM46EUe0T6qmOmyQvdDwtQK4hjfcU41UoJ69BCOcto
LlAAASh33Ek8mnowR79Y8spRv0jHhUXjYM++cN+xt9wE13XEOClvNBZQD8Z8Jz0kZt3OHtLTUVs9
//9fB/SJ5lcmUQctb5UcCqidBXOl0/4bXDB2XwiflWVaS8PmlEBKBcLQKkdIDNsvPXW0bOPF6MU6
CXOadAKJ37czjFSmzV3Sm7ra4RRfZUD5E1Wxv8W2vzaTJxD6YgQEmzuyPMRTFXddEojLsGQ+/jN0
oH8xTxKfh0jKlFdiFiiGe6TxQANu6dOCkkc2yxJH5tXHon93FIcKZXhiQ+pbMZ7GQAjfLo8kmIj4
xKiyvk4YNdR+Wte9/HhbztvaROfunxyl2xQVoJGxxUjDv3fW6s3oCYRdRtvtzQ0k81UwzsTSDp5X
BRqwJZJIhNq9URpw3hJcJoC4mLfAq3eD4PYSnoAhpCIoy3MoifMKtA11V59MGR/1yQoPr+q+Spf/
8wwtlTcG3T+By9jkx/f1pFNA39y17U8rsZdE/PJQh5SbusKFCbNuSXAIb8FMUO4BNioE/KEeEbev
GiVeZA5oaRCTuD1KVHaRjepjBUaHxQX72zyM0slWpUFBKA3iI/HL4Id/S2SDK+RLBN2rkzKwpbm9
RtgBUDU+UyLo/LB182EXHZ0Gi3WJHbwSwvhNHiSeAZ+S3oC0UTS42BkhPLDjZ14ULCkz+lX9IgHM
s2mjIAoLs9cyPu8hbYvi4GPc2EV3M1lbk2KP1HtaWfV22v1vg9b3vm1NywQLxKH3CBHbivtHmlMl
IWhqiQgT6cY857S4ANZd57Y5lWWc8sXCN/LEL1wEoH8viz1f51QqFWh91gUOxTVD4DFnXWScuQ2a
20KSZNV/HEOUW1/zkW720toq+cXgP5Pe3wwaAalXMUcikX8tYf+W15gEGCaqAoeeIjIlYVXB9e3R
JTKySgVRwIKiz+8mPHZmcvuMv8iFbyoAhAMXqjYNiAFJRrh1xkQ5+hoxZIcbOJwrzV/5zOsV0Zhk
y8bvN8OJzN/8QYTqorvEJB9Bv2aTwQ+lmnhyKxlT8oTA/n0WrK/FW6o9DG0S+RtZ8t64Px8QvBVq
2YvvnQsqhnQOKYFZvcsFDDCPNOk+qsNBOKJhEf8bOllNODKCIxSfjR148+HYYof/Vt0MtWvrRTmw
N33lhiNPpV5Eny6SsKiLGro+pewsBPCcU1xYl39E//WfIJ2iiTY0pi6eXjziCabq+jgeTcTNdEPc
P7l0Lq3jossgXPIdvmK8xNsb7PLxaD/cyXKAcktwnqJT9D1Q3d8A9oQH/pPciaG8qlLMdfEd7t6A
bUjA2xYqh6YdoT7z6XJAik0Axn8D7FDdRgn43EcnsoBeHxpPqC5mn52lCqbdgR71wd2GMON0pzGy
JEbVjngY/2mJn6w9CyTCampQcCjt6uslfP1uEBgM/15AmiJwy7Ga3Z7ZewB+9RkQFqPsmFrHMLoZ
ecItmLjwOu1O7j4/LnpAH3lIaEeYvAdUHjVgc2S+ILZylVtrkjCNUsIYRkQhgYQxcwloIaY2UrFs
uAZ9XW0WKlArnfycPgSbehgAqzDFUE9jUG0zabGPYvqpUSQp6KrOMStK5oU27EZsMdhgxICzxVQW
n3NzZLbS+uTj4TDbt2sR7kZnEBWw+CldEGJawlAFcubmsntgH90wjbwN5PLnyf+0KdcsJqA8/RNC
PM+lLLIX+pyNvLISRvgiMVTF9TzHdmun6xttGPampbrkqk7BZUeQOkipCzkgVgiSgLtgR7k8jSJ3
jiULoCto9mk3P1PfD7ueIbDWoUmJtR5gzmIS0UIQGd1WX3IhyPg7ia4tJYD9h5/KKHVyv8mqxyZK
kCHUmLp/GNV2XYgHXW2y8L9fQU6CGWF+i+8X1VQV5/ZjeO/aYDoj2V0HjBA8U/gHIecAt9ZHGOAC
tZHfGm3+JbyPPFrmZdYmArJZxCl8RI/FPTIO7CbpK52F09DDB2HcDacwsjIVfx/vfFuWUv4vKWD+
MWT59Zjf2TpIRohY/HbPjPb5TLQVD370BrzXeq3WWowyfE7v2FZGd5J7q7HZ6ymqk+CQeuiNS4uj
+3OX72DoStYTgEq24Id80fqerpJQQAq8vZ/ot5el32iwYpSECoVaAMCw7SjWWgwAcehNEE/LI2wv
KI6a1yqvaCWTfo1do+uq5NnOJHnDVZUG51izE/4KlQSY09oHEx7FnwO611H+RMQCxvRSt5sRnclu
tygZWFFfClt5yyqwXD3ZCqpJo/OzJ+3l8lcVYSL96M0Ams5g8jVtPWxqaIQocjkEouKj4L/pAEch
Af+1nFzj0Knp4+BpCauXjui51mRo5rX2YUU3dLMji/zllv/lN4WLvDrAstAOTt4Fo28kxw1yNqvz
WuO06jDDk1HvZ1MB7My6FhwBZHQTcPForys2XkdidFtwSVH/6xLo8/+1GaQEJYEE8pJDYBCVKIi/
3pcJc2MJw0ibLwvEABCqmcEu++wF6wNWNoMcgeTdJ00zTVsWgFE2P6S1QfBj67MEWunI1y/0QjYm
aCLENXJ0cvvAWkiWEQn6O78rpTNaiyEKXMtHTqZ8ASyaBHKZdc+77/ewp7Lt7uEEy7mIx64SZCVL
j8ODtKfXEobAwTXOiFdKr1eGXYoLEd0NPThWp7Wfq2S0RtE2M42ctOYmWNXOYzeGfXd3mzNgbugq
AoNzA7vcpJZizC68YQ6RXmSd/COmzKFnMQK5rxr0EYb8kpPW4TTfhwIFfIgabDfsfykBI2ghB9eW
gHUgRIq9z4tEuJU7oq38yCgeDFt7ROdBwpMAtko+7pF0U6IkqVyikf2sx2ZnpaFiKR0NmlinbihD
M6YMEP9WUujiSzlm/gXeDny//Haf3lA3+crgsOSKkO9WVnTk0Cfaue4TgTF7Mln5p8ZUF82tzcBC
gKN7HK3rbkda/qGVFMO9QruszMG0ok32WPfXNcYjSOSsgsoXTw9TcZEVbeScy7Jbn/dlqBDP22EO
JL5X6SLZte8i8u6VlZwIAt0KV/AkI9KzyUXlLridUNV7la/eWeXdirXkHXPfE7ytX4bK9CWolRAg
2spc4TZ4qvTYWFlxL3YguY5CkrflpYgzyXEGduNCW4iK8hUA00HC9v7Cqs95lsKGlIYl3VkWaZRh
6gmjlKZGhFIaV62EKLoiPKOXVGawsAazSo0H+JeVAkpUeY/+PD9VMO1O74qtIUcAoB/tO9EQXWbn
pL2+hbxpptv+b4WK6vnpfNlcg8beUmvlqmfOEdr4Ko71Uy06aDkkcg0pY8vwnbw3zAvIiACFqXmX
DFhXZTSjlvnW1pZ8ksZgjcnWC5/WJ8oR5kBwXxl//ZiL+YL5Ujvl3QtR2mRHeWb4tOrw32xsMHzY
REiClYVG8gY4skfIvHkPkZ5w+9LK3YCoikahy+4uKaOrcUIxWEZXqOabhtsrGrArbpblumfc0jf3
+dZRASadh8pbW3vlK3+9IrMHDOiW2dSE71+JQa92iEDigX5JCDiJT8OjlADs2ke5Gls3jHmRPDTG
PSaheR/AhfIUsLRjyVkXTa9ghr+T3psnJk78+mJ9QW7zsPVP2Uq9nVCL2KntcUuCdQNAAv3+vwFd
NkuLa9uvNiab9HOebYlaAfJh6wRBMBCd6c8tI47uaUpRm/i+rArN+2kmBOXE+tArSW0vts/2E1DO
WbuIegMUERTOcxX/GN87VTuxOJxeZV1CRxmYIXAf8yAeMu7GEdzE0C0Nm0thG7xVtH7BosjzZh1n
i9EIaJOTzuN5JaiXdOxTudOjTXoa4aJr5jPrgodFbu5bPjJuIxSnZlC/ZX4uEXtQ84y8OuJbw2UC
odUNdJzYhHN/7e36rd1fL7L+9LDgeUg/xkcgW5mS8549VPqZVfNRQQNZcyj8UdBAirA26xu/+m5K
1+kJrq0q4zIe5xHKOEpdVHB4lueolHccgP+vEKTYHcb4CrrJO2ruIaiqpDc7jUQgsPmwYoW6D/tj
/hPGe2hmTa/cZp5y0VHzJsEz3pVrtPvPPjW8oPOczGucuI1SDeWmytusRhOTfQYN6T38izVU941Q
Ig+2VV4Ytm7BSTucY1PM5TJVhfcj/sETuA2yM0kqHONjznSEkI+8e37IoxvkwgiJHmjKIQgvrrSo
TcA87pYA+fPQ1sOwIsAwUQmW1rwZ8rkAHfs/2Ch2sE3dQAFuYdt/Htjkxitiz14GcFRG7BegHDo2
pl74ushL5DjzDfRtjbqJT+q7ZlMlIf++rrmS6ErIeipYaNHVas/7juxRDFVydfyZ28lGRg+xaSDD
swqEaBDnEpaq1wjYEmZ5sFIRv2Oo0pRrFOk9g0NUCQOpEQQ7vwT+WgfQh8HtzvLhVB9m2tJkG1zq
SwibjlPUsaekEDYzGOs2fvuBKKd5D8ColGrAo46d7FzfCSgP+OLwpXIy6EE0RxBwQhdiBB/7PcHk
v2/D7+UQb+P5IBsSuQMww4QqFLeORqaZQisJVOwGjno1VgIDIeuA5y5Z+lPK5oiDW4so/RHkJ/Da
fH/n4l18U3gjAD9woOvxV6zTR0qjnWBZGnGJMkyatHQWfd1g2dn4zWW3maHWFVtu0cKzhaPkNfUu
NK5ox3+0ajnpEkXrI6R53zJz1gnXKsXYO7PxaoazFzJ99h895TouhPeluPmhbmNctkZSBuJngoDe
UYrvgOVVCfL61gLPgBc9YoloFS8vQ5JDFif0ww+709RThA/SIDeTBTFUMfKIgPhaAF5ms7oCquvq
z3iRc+ocvOX6I2LII4xjSbkZIGln2Q0lM8QbIdcSqvBkrroKBTVKQi5sPa92ZNXNEjbulBGpHyhv
qB1p7CK1ET/PgZui2EIX1tdjOzmOiyWfCenxG/TxMi7J3/b0nabw25e6dZIaJ6U4so1z3Cb5nWPj
0oM4cSuxrG80zuhoHQp0LxeZ8TTarQ4OXOAn4gd14mB+pz/EU++cihYqfkfKbfJW7T8uylS0G7Rr
JlNQuYm6NfXzPRfvJCo/xeaPl45+kCwt198pQ6ZGb9kkyrCrMw9O97Cz14hpsaba8UhMXelcORDw
8aHoqo/+Jm7dB/oi/y4LDYNxSKJQ4tfKqM9FtdRyQmolOBJ2nmuL0FdhQ0CAFvbFW8BVmOmGuMwF
UwWkgZOT1eYSy5owKwj/KbqAmoCuSDVhnuVDE+lIIJnfirDRtQMoLMQpRC5UGl3cG/Rwp6vrLRba
egflq2tq2uDObKdV9FDlvDLo7u/++M62jtkqE+KQYVyhzJrratWOC06XknorZPJBHUhpYM670Kbi
6qKmSNuCaMVFzGDF1BNrI+weGkP1Ae8mKwK4fJdu4OX0NkOdQcaAIf+kjDPq6i/QjVIGafPhKom6
pZ2abN76Hj8ArG9ivrqtIB0/iyyUFHz17m/gJO6sCYjvVfu6UJ50EPB9iaQou3VRYqAs7HnBp6+S
30D/RaWF37qONo6pDw9K2MsulRaz4x0gzhsj+ULjJWwMHVxa5A1WDhp0tHXo/j1eoZ16ik7i8dHL
+Se8tS6ALX9wF7Bp5SDrjN17Ctl8EB+OpJKMDKV5Q2T+AXm/VWB3RK/55VVFfT3T5FgwlRS9uhbF
el3pLOazkijsNErCCmq3RqRI9yQ02KCPBuIIN4iX6q4rxGWqEDuRr5NiAPuWoy/s8rk38S2XLMqY
1hocc/x+j90NtuXpwTxmdH1xnuGtjbogPtgZTAdt4QyIGTwoaGftxXEG0JFld7DNfb1/ws8aImgT
yujPdaF2B9ZCq3scCBuwxLdaGcr09SpGTwThjXu8sT6mNpI2OKlGVjcmb4ctM+p+tO8awPxayWcD
tUHCgL9hCumQ0Jz4UINP9AHRkaZH02tl6CbMqz/6napclqcKYAkgHVXK8Ff6eqghj1dy0IEu/9Rf
mAjOU2Ne51M3frmM4Y5j7lxwR9L6dKfeg5LUuMGC9T7gfh0sJnbd4ZYHYzdCZAMiCfILmIDWWQT7
hHKHvxid6o3kbE1F84gIYGn4+rQdQspKquhicnicR5/J77VOhDy/GZuFC3SdEIT6eLUycdiOeJw1
0f0dg5aY0eyeV3HvqlEFk7q0Z3pYV94IFcLo0XCdyKq9KYO4lgjfDY+JNwxJ5nfXVjLA9ifB0xcq
j0bayLNEwMUqpab7i1zqX4kgI6NZ9w3StckbZkUwjxg5dZJLhPMyqYmsptcYR0g5Vg1RtRnjdeCs
XhKQqz8x72luLko9+3jC2+t7OMcxByQOKZCFb2E21UijUsioDt5mlm9l7tFmbWqO+h5Kp2kd9xOK
5uzUcE8wikbHWg7EiLmj05e37elzIUlluowxjahFiRaWm0ZLj4lJSlqz9NcKCIbA6wgHiecX68by
XkrTzpU9AtoIeqMK1/3fjAiCAwUPxW1ZV+mNs8JZavwahKKYg9/ULMR/xFGbQKiJLBaHysHLsJH7
lZRW0JKl2RcrggUPmjPihxku7rD49tw4jFtg53lkCx303HjgUqOFF5SkZi8GIeTrNSd7rd14rCtr
Gfm5Ozc79dlgpHgjQbQtlek3+xX1A+TEwPGOb25p3gnLYFvp7NT3dEqqoCf3d+qeAVgNjDxPHxfU
WcJT//h8GtZZyxmFuJkmcNYoYanxevNEt/elckWZB6GNAi7LsQthfpCuXjw/3iWCXxTxuc8QKIGw
mZrbjxhXHE4mkVptEOV9mcKRLilQPMG0S4P/McMQdpwevhzIDzIaz28XcqSKEYOvHZtzafA4R3NO
7hOXl0xJf7EAkCITEGcty4mmz1z0pHMA5DYvDSIt5QWGcCW4ujxlpx8TMtCtNNr+F03or7/O4ge5
oZK+7Ky9RN9+RP9vcRoVbtlqiljyrAf4Vaf+37Alvvs4vONdXubw23qkQKzxXfbapaAsZ2p9ssYu
pUWaNvnQmiSr40pm80UER21tFe497pSkpTJdb/12xiftcqPMtI/zzSdlxwrlQ6XghGPYCTzwpni/
O3wMkNSYQQbkrxUreljMaKOvvH0J2aXXrKj73afarrqe+IjeB7KQQHxE1l6ffame0ewjTnXpSjo7
u4S55LTeFS+ayeckUvi0E5yuQ1GFUxuU7GbU0pffsSA9pl+t1eqn8fGjTYVBMqrs1LgHLTZDikA7
YkPXknE9fRSbFZcABEkj1F904yiNetqqezl35DJYcLQicO0ZhDwzAKPW4r6LrOm6rNwoNTJ51H1Q
qyN05RSPgcLm59HT5opq0Mq4vbT7yoFrUAanfUc9zzfX+alrx9Bg7KjwodgOUiLwCzrJJ6ovnMPh
JHXocoirp9IOstSvHmBj6KAVUVD4CYPpYh/tih1UA8QpF/MqrsTXsZG3aF1zcF1hQ4fAdyFaCTTP
g41Mrjq8Auz+3syNs5mTL2iNGCHA4nVLMAQAqRamvFkU2KbUhWnueI0vASAUeix6b5d/QCCXqPz4
AVCOW2pn5eQfEAA3Rl4nc9+hW4UnPBFCjM82yu2EAUWHK6CS4QAu9mkFe92QUn3nGrSA6nssZzGD
miN0VgjWgX7Ejm7n0CXVNFNZ5vOARG/9mdymFrRLznVV8zEYri34uSczgO7Yc0TSyUO1LPM3KXuG
FPI1PCfQa9gH1PqZQnaw3joruJ+rHaXFNR0rIeTRueJWH19vF7MR0aux9axzlqRJiPwISzb2DUIH
7PuJuPiEnJeVvc4o+nXZ3FX0dT0AIqjqnpxZxzpybz6nrZ62AL7+vHYHMfBiALs9rrIKPqn34ceC
pagoxXW5ywzB4O+pjvPqBwgHagV5tL3XVi+Lf19CY5sCyCCVFb0lemsV3AoYiMZ/eIhICYAznA+i
7cBg3zJ0/8k0YrlT+dED2IrX+97hVCquPsa1UjV3LF8r54MFrQNp7C6KcvfJjdPNS7QDELiblaGR
BKaDQcZLj21qh2bVi/lBOLbpm4zBwwx9GeQYEUcHsm9AldHxPPySB1mJSaQ11dIU6ohks7vEiQ5n
yLSJEBmt7ej0DJCgvT9OadQUtlAIV7uTeuJ4Wp0tm/0IPLojDY22BMmg2N9x3USHt1512Xn0pCV1
Hq8o7z1OFtcxrUVpKdUQgA3A2z6CzeJSKNpNl3Vje6V4n97xYMWRvTBW873wb5Vju+u1MJGdPhNt
DrRmaPC6o64E2+Po0sb84qMzxs1QCKoZESFI2Ufzz++gdHpnXYp5BozIcXuxSMefxLTGBJK8jy31
OmHxb1pDf3uEV5ur0PtWgsvMuS/5fS+ovjiiWwHFIV3tl3YQ3VFFDquFz+HJxBsBaZVjhMyGpvC1
EFiWQs3USRTj2UOjxjqOx0Ugb/HXuNboH09i7pyBQwQi0Bm3nSUrbP+Ns6h/vyFJVhoKEN/2lhJ4
c6iwBb7pSaFTm1WU0Jx1DCrTn+iTx1sj/8ENlplynCXoR/P6+joG6OG3osPuPai/iCDcRv7rm2Sd
6NhtZ9HeDGI9LgFVbxqI64aY31zWYPbVLTFyqBPizVyp1vdX+JRU2Lnw9UPpkSVdAXS9dj9rwRkU
281uYizPIaxAACZt2Cuqtssm95IEsF1K1wFkUI5KUt7Ve1qkB9sr5TJjbDusotfOifldr0Ljz+sV
bkhn7fnJX/Hv3MHR486DmSNkoDeGpjOibCiHf0MQXwdslqy3WMxJ84tZxLnX8K/y0Iy2oDrUYV+t
Lu0Ecrg7khxrdB3Y+RJb5gU074ep4MiuZyXEGrgudyvO84MWdfxXWuyaXUSaBh2r2y8n04lZYrWE
36KZTOGdAlUbbYGICtjadoULulZdBDYxyTxU/m8vOQZTazzpgPGsUU3oJ4IIRRcHmjopwQ1f3Uge
SwU+k0rYZZQn5Pe+UzxZEgRTYL8bvZ4lCCqlpIA4sh+8jGsl5vNY/NRdnwKdESPuhOA0FViiWTi0
W1wsUqFOAYd1V9tFqE/nTfpaGDshIxHnYtIvdjTTiYvBTd3eVOwzPM0cHGW1rGzhFJcrdCZKVQOC
0JQjr5h5cZvpkUjMFQgeSX7xThv0szbefcmuVRvwuNYTigSRhNsYYeFrTnlg+WQggJQCsq3mnix7
04yML28lHn4nHfXL2ac9LSljR0aa5tj0dHyDHfW68SItBHrIIL4LomGiXqVR9/Ta1QZCe3AkZQUa
Yyd6gYJebi2CcEV2+P+Ba5RX8WJq/4eWRXfwhhYGI7IlMXnawghqWFIe+25xhc4u52AA2JTLVJ+i
ya/+oMyxfXVrpe+83dx1ZWN+CSBZrPYFmqIcaZlxKTQvIDv7aWsEGCJ1TvwQgGps5B0W0iyKstPc
SZl/Fg73BdYuFgfXQOnAe0ixl5BEQJoWhK0lTy6qZuoKH9MSY1hw1Uj8xu8Eplbl12leGV8x3Q5m
o2VfcS5xwtseSHf37QtHnMF+pLWGEHulmcYMP5OmDOhCCcG7+9CJfHDm1Z1MGrL6kcGd3qx2/JzE
ejY72UzcEoxt3f6niAJRKvNC5tA9/PoyvlYln/+CpywF62jc8Iaay7a4MzEygVuPVEJfUpMg8mln
qNNcq4yiv5RKMoBBWmM/cGvM5xMuZxnlsBty5hY/BSp2DoVzGXH1YjEYq99bLIyJjWOEm4T2wli/
Vz0ZioKq/Ph6TNDGWcViytOk1By1zuGl9gM/2VbonJQC4MZjHuJfOLDqKF0z9WwuRteFpRWXaoJ+
jxngwhVHTN9L9G+wPGoRhFO56YkiKXgqet0ZyVlGQRCGcik042ox2NEF45UitYDU7Tw40FSINHPn
pE/1usvrPTmcMTx9wc83D3MTv1Hd3YcFOxm1y6x4020XgqNyLvll9n79NjPexH3TLIukuWiXKbiE
C7sOZlE+6KwzbS9lW5hHIP6BE2bksr7x9N1LiTmROtr6Ng/lw5BTbDIhYzUuG7hLTrzu7j3VbxSI
hONWqcbBt8RhZmeE4vjjTHaLBs8RA369Y7IcPgjpG1CXDPNCnCDMbEtVbZWBvSfgVG45PTnXcUaN
ZIa3Df8pQU6W+fZCI6ga8RrkIjNVxrMRxVuaZUbmu2zebL2jSpYTh8yN8b9JZM9thfS0iHK+4rsP
bI75o/Tln/M+B/e6iUmqWgkEsC7iLlNw0txpOGV+uvtLv46CIAtU5C50E/GybEWaqc8raIpvqzAN
39/F83vwOOVg9D/PY97bJH8c16VOKPbMrWeiqPmED3lU94mac1s+axlfB8SIWVpDdYPkgxED85aJ
5JS1T8G9wtgysglTzHH6A1b1B50eto9I221s27U8oKPexKYMT8qsjr7ovhipQQpsJPl2x0lISxdC
M9T4y3Yg2zr+2H9ozijNuH9Qbc0uX9Ea4LVRutC9+o0RYnyrYXY2651DlEvEV6JLEsBXoxqFYvEz
8RyoG70XxDLB0BeC0wLR4JORljcfqldr/aBfWw/3keMiGJ/FaRV+wv+fI1/FFQoeATdtbdrYWQRq
bqM++5CmM6w88g4wmA3w05NGSEWVoxYpflmT2/dmyDdBc3B+5Knv2AIWI04/gqzTKcC0mOCfYXok
FkEOTHJrnlFM2qvv8QgUQNMPOebHWlDVJ0usuvioRV6k8hx/mQJK05NQfy6m5Zq8yVV9UGNrsTtM
1DVuQ7NsP4fj1yXGlderTB9V1561OwyTsL1rGVq0O5HZ7+VuD94msC/dCftIiqzvZ/G/QlXdcurZ
EimLumWOlV4ww6rbqf+tLFKtwiBCKEQYbHua+AxN1s0GqaneTdaq0Kn4MBUHDNYAMywIa2UYbrOL
Id7Z34OS141xvDefPh5aZ8iJvNfv5AKvA8Bi6Wn7llxNgHjuWgP+0h3WMiUZGNC9nA1IapwobKJG
8Cd/jRfr5e5kxGd3OX4o2E3ypSAxTyRgmdToYJ79qcmbDiG2EAXOxkjtybtUwCBZ9KaDi91PCoGd
rgfJXzb3W8SVw+2VrjadaOL9yeyjc3FNx7+XmyB9i7quhQwF/Lnx8VNhU0TjoLXxzjp0Poj5cAdP
/yhDSxKcYVpdwwMjmt/zbcgcHDJ3j94ZWicP5iT3YF06eRxPpn8QZdWUcdYRYNiK36ncatbBWs1+
uEZ4+dPhuKEDiNsAfUn1TtHHeDR6I6dGMNovi9RYguNRpA7h8Pt79jVtoRfHF40XkwozG2XvivA2
ROa4mlyL7Vf89PFbmUMouvdTA7cNpGZS18WKsrA8vN8n65ht/anAh8i0/udtxk2fYXUkAj7zHY2x
YGrhdieqlRyaEszYIzzPrfKOFTgvya6t4HWD+MVb0VyMmXBOZkLXv7iP6cXcH2kqyDiVJdeRA7uY
vIw+IQ+VqBzuRKqg+bA4aqAsr6SYvAYKiaaKpPzo42uMovS01lA1m7pyor3PDdn4CQF76vIpZlPA
4sqcdUZfWSEJe8845fuVynEPDRkGut6tB5HL5tZt8Qm+er8ki0Q5xKI8wPYOqxXk/T7ZeuLMfg22
ynQI7wXFVZeE4eLvYWRmQbQpLy1/ja+uzs0/+ltQV6+IUsForb+tRSSBMKXoKU61gePlpJuLZ0oe
w+Ix/1H1qQ71VfWlBiOxsX5uibviGJKotO8TY94/MsGrtYWtff3KZ24xLGbfRcnpSYGRJqJMWAji
nNX9BXgH40Q8SPdqB110hqfzHJ6Yoz++wJSwEFgcGCm7trRUbDxq0c+mAYoS+aFA/oq4ArWB/fFR
vyrsGjNZRNFBdsZMoRpdx7YBVpYIwYZp2vEC9nmnBHHoDhOJydrNpBN1qsS1tdhI0GZaV5srRcs7
hdNL2OMtrf+ygi71yR95ugEzB12rkrWJzododKP1WkiuqSw3/ZOslcVA6QJx1lM1zPO1zsqNzXK3
OBpuFMQB8yN+9djjwM/FBL8TFRK5lDudNTnvGH95VDM/EbOgdAluHaeslTXo0NZ/YliY7ISGueX2
70hYeU0nDMxa4m1sp3jUA9BggVSIQ6sMbCIXG012040ZOYXAARrxb/Eu9QdJ4aBtxvXv6XxS45YM
sfjCZYUy91u57n1Y1xvbanCGDT9el36+c6ntvotsa+gwzdZHQeNBf7NfSrxmVvFmBrLmdrz1Msim
CfjlcVmm80M7l360wOttWfhL8vZLbgaexi9+aviLTkPPh0/TXi0fF85d1s4zZkS1Jf78o/2X79tO
dF0UbLxsHr/IEXX+xptseKm+A8VcaHTUcsh8CUezbY4BvyXzjfOT12FJ7gbVACskCKFtIBesyM0z
CkfdU2svy6vhtaMPUi4zSlI5SY610hOPlBLDf12/UJfAozUweyBjblLyFthRrH0Q4LuKB5W0YCs8
rS+d0I5nr7sL4x6m4ifcn9yvTtbr6ULxArUzKdBWyr9R2TqPOWpditIfLZ25c3DK6cFSUFUQIAEG
34n9rswjPHGFpoWxYdHZlMMqH0hjbfqfgguNVjpM5vpMTbgahNp9fllDUp3+nOCRg5fEQE8FMWPq
N+xTuy1puijDIJ4ZrrA5W1IYR4qVJCxjAg90CYXkjqP93EFchjG6B/PJouoUn5pwNx7n29aAsC32
MDxgdLTd3FAKp14pyceQOiLNOM4D/dA/Fdtw1HNmXTlPnWq8B68kkpCnuIKMCb6nfR0yrkGaJNYF
pvkP3Eql6P8t5CYLCI4JxJcgpZSgXcysNsA35RAC2CST1tP7+g7uyVOH7nv1TDPaEmwqPd+rfaUf
AGo+6PwREd6NRZs/cd1DF1qV5VNoglZwjvU/dWWlpvYAElNJcs4mkGLv/Zqul+5z0mxvI6yngLyf
Q/4YOO92Ru/BspWi2fpxfGmuA5y1xEWIFky9defh5+txqNuhciCIZ/dUWhTwAwKEP2rjjkZZN8JH
t4QIOs0JkZzN1p6Iv8Ouj8Pu4pppxF7yt1el8I7CO6FLXMkvvrtAzclsbnHL6whqE1WN86ePiQyU
xCSSH4uU4xpju57OnyodkJWbpJ9nYys04LN4qWQyo9y0KidSZ9U9pQDd57ZBJg+MRKJSVLwBMNJh
WHA+Vr8w0OSgSZX20U5USivX1IlE8CM1Au8adir9uacjX2czs7bDknJqIwYPXPC1r05aPFAV7axv
icJPIRNFWqcuTwcKhOJqbbGj1Oo6v62iBET885IUf/Xmo0pEgQK3ynRm1isO0vfVdWibF3hFBc7B
aWafzLWGvIIpVZ4O9p420lY4TY0kALYXWGxAI+0DZPy7BLHz8VZicJORoHky6w0l3SHuSz3YMidH
Ts6NpfXqorL4q9WYCoMMZaUPssebJvu9KnFmCsXdWo3qoWEHIYfKQhVgvxFr4/0lBXHaXpTqTAp9
PVkP/GidSuja/y4HZjzNK3fexLoYq21GukErJ0sKNuMiUuRiW1AqJLJZIixPKR460PKjy+DDqtK9
lHmc/JvfDRYLii6+UsQmLqsL2iLCgSpbfBLisBzN8xyYMxGiChcXTFCO16Ryi5h9bQBeLl2kxtUL
r6ZRyoZGDRv0zwzOlru9Lv6Tu/UixpN8PfeSSSqOpLeq2W8XICt03i+m8Xyde8No0XGOzqzKnUzi
R14bNRgVHXQkUDc3eR+TVqQoKvyyNC5RteT7vy/XMpqVfKM85Wjl04g84MMPlyrzwT5a80XY5bEg
B6P+1Hu2ItFtrQInA45rx40YZCz2NjyF4Tu9CSwwZfD6R65N+Db3Iw7ZzqszYFn+525k9cTr0jMF
7AaOkW41MLmrtnW4Z1+F2G+W5pmb0G9BInwq1K6U3NU/WFUiOA2GX3XgTcrW0RjfY8OveP5vV9nJ
2iDjmIUU/j94rUrWJcHc9A7CQTVscHxDNOUeBp0rEQ/2D4pPHAuSU7nukKJXe0d9SZnpNOg2WpZv
4jYJgWU9MNPZP+spKYO9199Cj7Itjug2VMKCrjXYktBm8sWzhK5jcLdo+G2HE0kSSBZ06uVxIxaW
g7W2bapa57sFCiX+l76+Bhr0kgcAaydDUBqV76jX3juvs0ALerTx4ZgxqHdNRWSuYwhizgW0zwo4
A0A2AqnNUYJllC6iUgPXtErLTeujTaOWS1ocPqG0CewkLjEmIsCl/K9diPpXgP/kzn9URWHiaTNb
UKwDX1T/rakjK6gz9M23Lmub0wSiqAlGAsJQ6ORx360nm4GcWx64oUiP1ZvHl1jkxtMRInpYiXl2
OWZ0NrhBCObyuA2jYspDAgKbbjZ8R5gZlA3kXENrWLkCPeYg4VVA5iuTHZ3p+tq1BdK8H0j+IO2t
K+5w2gSobhOoFDy1FsYLiniSXz9YGHr+8rOuPlG2CFuduIq6Y1fgl/VHViknz8TOBy4QaVbk7BKR
DD9I4frsi3G8YamToOiFExlW2XYiZaVeC6r+AjUY6iUivNxDJBD3ziX8YMJGXz8q7lC1n6NEOUj3
o517cxwg1Np/w6iQTmKxmon4o8APhkEDiKAQ3XUHH3CB0ljCB1WS/ng5Tc4S4KUIzeww2ZA7eWPh
iD8nuex0eUJIYkZcdln6zoVKTNpyvam0qmo5WqddWqMcEg3M1h5js7usvcupr8K/IdA6KSU65w/I
YJKy5VkuOofvI0LiSeBY65ChilvZcRnOFVArrn58MmEqBby1O8jhpWgMJRnUkwiO78KCFVbd/AmH
5fN/XxYsxrJgME2B6EUDGvlVVQ+KOnyQHQHxoFcRFJL7H0RGLYl8JmIaqs0cpHow6eg5OukeLXsx
mFaAqxjAyAS9Q3bKvUa3CpKj4+NQ5UL3WDPAqinjIhZ1QBaltCs9wbo4kuNEEUEM/ST/AwUnoCFj
SXrnOtKJoYu77svd7qYVds9gTAcs4wi/6COdA3s/uyVWvu0bqOeFEgHaGFO9wtoGFIw+9WVgouU6
FSpqn6I0pJAxItw/e0WyQ4wEqmI3rbwpzFAQmaWmkjTkKxBICayjbPvJ6v/e63aXVSzrYEmQiL2w
Hbt6WQNLzpuThGsziHDwa/ge/4vZG76VBj5sCOGeQgEbg1Ao0tI9jPNzo5JN4u3CMGcCmoIjDGFM
iI4SoxDC+GVEKI1+vrsscB0ziGPZ1Awvl99FlDRlfLh2fUJ8nOx96jOaL+4E7VE1Tc7mEsZTI0zI
ylmxkA1lCY5XEVrQwNsh4cW+4lJ4o13zP3ucucqZLvVW8h1ajjp2wLpK2f3DpQbemRDWJOUn14P6
VyjkqoWqz0CV5MZxKfPckimTrrjfRxDfmvRhFyihu5qkIjgLeUC15RK/O4yrG6TAt+D4giBOmzV9
wSrq+u3pp5ilgbLJKLx5bxW1xLo5Mg58WouJKK3TM/aqN8Z0SCZA9aIZxIylujCjYW4B48SW6HGr
9bj04V/s6z1R5hwLjbgKB4pol/sk22SfReh8VpYidsWMup7ElY6a1X+uX/ZI0qJFdDEupCYj7JHV
FZy+nZBSGRICmX7rQngz2zWhd9qCxo8wHa8ItgJLrwo+g2FUfUaBYg0TQY7VfWaZ7F5iLsPbZ2qS
CgdorABvM3gzOKNhloe7JsB+ul/uH8JegqHrfc5mFB//sHsHb5XbKanbvSFDV5uXSvqsSzjoXaPL
xYbNjSIrHRt0ZEGveW2qnCx7DTDxpbTmkdnKvfcT+iwc13QpqsZgIh3p+XpAB2LU8CoZCrD0J8zS
x72f6IumHvGnC0VLtJr/YuwVO9HIkPVp/ZvUppDULd9hKuimN9X8L2SFkKA8YX79Qlc4yhAgCcEW
jRmXIjmdyLMtWrZuqMlNBMPeiCazIrCGKRg1+u25YALhooGcVbPKb2dUBwvHDLbcWUSX50RkNJEX
aDgIXms/oJPlDgbTUFAV/Jo/C5IsHwh5WCY727bhrGD8N2rAZbnFogv1l4v+jvDBrKgNdJ7rxU6M
7l0zx01QyYvvGlJ0GWTLwX2nuHMx110AvIf00ywQZp3DGxf0C9ecVBLLVsjjs9qW7TaY5BRb2C51
2uTN5Y1BF2ykLUGLkXNI3A9JbnY2a8i66Ni/zV/+DB9T5EHskLP3APsUOypS5Evn9XzDAsZ0RwC1
2O15vVp/Xpz0515GiTLtRAPfWUNiDWH3cZlxDI987+00KbheYwC0xTASwZYSSA+pOJuPSFtG6c/8
E5lU61XQDoxq0un5lWQt43LoUgF3GkNQW7hXMpTxwsw4pqXt5l2AuowxJp0115MmfD9/YnL2CQvw
1oA5feQqIKjR80r5gxym9MDNaNLPdfts/t2PSpLn6/t/tYHIhoFv3d8zpnah5K12i5n3T43NthZ5
sfpjvg10awJQMneGYbRoiA+eGa9ZmjG3ow8g2K+73E6R/WvdCqAnmjZzd+UCPmLSWI1XRd1S4DVe
VIQRHHT8WoarFkubBV0MUWiUuj+GWrnGVIr5uAQwc6KaYON1R9z1tswKmgABX3NbuQcUMOtKWi1n
zXzM/RKRiJlzvFAB8Twu3ohb4U5DTWc8cNHX6zpV1ydWU+/lPxtm5rOcyfWQ3MOYZKBuXCb6O92q
vVm5K0jBa+Xx4r4qek4rbgsGAth1ddl3rY6nsTqH2NJAECIlRmoj9W/lBUg8N7AeqzcOWdJ0pvFc
hDiUc4ki4Jb9NSbHCw/HwbDq1L6S92vPunaGiN5VO8rUzFBn+nx+HfcsNXyuX8p9zk8hmv/91pSc
KIQaiRvN8vHkZiHb3Em215kZ0QhYhgTvJ2pms0uYEuaACsLsjqSIv2xQnJb5vQR1Zf3wB8yeVW5S
G19f1eDtOzvEgzl4Rbcj+jfJtWZ6SMIlXbwX6jtX5OF+XwGJNTGsrxLrlGEXirymfbp5tDgc6tPi
G7gflIXnLQPJFb6+BhFcFGGw7JJAl7DbOLsApaHKz8FOzC5xTUfjKmRUJLm4GrCiXoPRjltvGtec
Kwn/5B/dsF6AZR86S0guW2CAs9afN0AnoKxOIFP52bIVj7SIzgRlsVSgBtALXdUh2zVy14HhRRnH
WR372GegGuGdLvWd6yZF2kvCOEannI6xL8v2dYlv5q35Y4LQb+ATxJ4NzdM5zBm+70j7uTNlNe1P
iH6ebRgfaLyZQnY9h2Zx4iW5kB2BrPWEWJsCUAxtkm7HrIVuRRPuApyraAZUZkIcdGR9FbdvW7Y2
pEttYa72idbPQbGjxWJZ7TZceTpxwZ5J24GYq7chL6V3ce+V0qVarPayi0Z5dKtO5nxOVJYxVaYi
87sj+xWVvoTq4mUCeaQTWrR3wzxWiEsJCHq19Q0XW3qM7t4fpIKitEdaLLhKvCRJKgfp28nBhKeX
633ePEdbmur2/eycGtqYovx1XYQuRJjqjewy8V9/vF5A6Z5XNEeGjjs072D+lJ2eqB1ezFiZEViR
LyTEQg0KehoeHHz5FMSd4WPygj7Ov/+Tk1h/BAcQ5D+LhY+456GbJd0S3f03/353ES5prGw0gIcg
YWfvWE61BJyGqeRI1US0p9xCReD6u/F/BrZVHSK4RLjSfixD3vLWnUX557IB2K9zdD6lALolkpBD
KRNwszpgy+Stm0yrqJs7vXNpxhrqJbZdounM4+CeN3VI0hZvrsHjINScOCtMHCYrCA9Bl2oQeH7A
F8Z7OYxgx19kIy5VzRhq7aIb1jhMk5Ji+I7t3DLlMOQx47A/GKakSwoUr0JyAHX75yZ47mrYUcLI
WP1Gvz8Yn7vQvfSi/4wlOwOkpCOXJBKZbZpxImAtXkwL6Z1XBtkYslfjaOUpdMHPo/2/9E4HuKLw
muKotEJcEwQAKQ7YIryDm9Mn9ESsC7Zdd+QyV2I4IyP9ftGL+q68wXmi+suFRMfvtNTDIAf0koHL
DcAZ3uitcVy4lDSYhEQcNY0KHEbt59W7g9/z8EdVDMZa/2vcn9BmC9rXMMhIQq3GpMqmHmP4giGK
WCFKvGu/YQxvQYSXW8K93b/CaAqY3O53TbX9tjWbVc9JWMAPs0w1pFXt4KDPKk7UDaoHrDRO0Vx1
gWP///sLc9bMW6ukaCs6I+ijxLMir3i03P6U2J/Da1M4eZSgqFSw7Dc9oKySASsi3NrWqB6/Ewly
H7iB17Xf8KxR2iKplhfTyCo+hYrhe5DEZQMpH397JLp7pMvY4h6S18rD1zKAKIlP2Xf49qb6S9Y8
SMO3zEnuN3x9LSACWrn1vc4EcgNZ4aEz7SUwVdAS8t2Q1eGjv/L0W5SGnmAfcggg/f4MOgm1BiGA
PESXaPG7JICktSZ5xM61AuFZxCsI31fanLBqplOEiqCS2Io1HeDjKIFESuE1zEo78xElb8Zneoqk
QSBLem/qgVB95ITjJNErSmf0pAyURXe4sMtEfBhClKyB+y20ZLevfZOaTEg/BGT9ql5Ky5aP814M
OXpDX56mEh6Cgm4nHGazFHVR8mGf/Bu769+9ovjuMgCFrAfKEbPMUGH3Y1kI43uCs6NrVz9I5GOy
E4wV7JW1QMAF3W0FCovvw9jmSWvt4xAM/oS5916yHx4qdLDRxzsvK/Y07mbYDEagy0QzeYZU5ZDc
WNXKarmxR27tfpoDgmXkkIgocSK0MzsA+oQ7bshjZCuvqQ2JUcmpe30FhtGbdIb1vNbqwfCgnvPd
22taXdpyOtTD6kCSWBmNd7UjV03FZsg9RxhRauqWmrWWPofERU8EQOAlWlsLTJtwoZwtcx6ZflO+
V/AVYYv3DRv/oaYNFtn+7Yl03eFvajlHtb2GcPEIKvL1jKaD48cpTDFehEZQStx3HoAsbv5TqiSG
ugJdLe8bEWcI2AdRYHWt5yyynadA2QFaszo3zOXvb7wLGcCICejCq3bo86CIDdJvon1PM1Oa2Ebt
75imAUeu3AlSKfhGBsm996ojsPrPa17VA7kIouHnqpgXKcc9EFYYPrCBPpQdRs1h3hezEatr24n+
Sp9GBBPoUzsSQb/B57TivRH3I0Us9GooHodoiP4tbK50S1LVkOjXoCPoQ+WT2rmHOwye67oycloj
ZfYyPohW39LVT/1Iuw9brxx72uLf1oGSwPL4vecYVoLVaJWu5yrrlmtxF2VZ3QwHp11pArHCfYVe
CKjmJ2XWCm/RRg6wbk02z2H5pAPf+a6DuXpJun7RX/LrG/YxPMpWWdoDSoMthnvvdno/Fw1qux/s
+CCY15vXfhFuqLm8x0NMeip4zp23eaSqa1e27xk/ifafGS+5E/iu+cdmocEz3rN6m7G7JqJsItHl
cH39IRUZMyQDk9DbfxPjFbdWoqFYM2ULkkExHxHfhV385Sxnc8KYchixMrfDt8kwn/dn3TpbaJpO
LJqnrVRkybcv4ZuweKyU8zrt2Bo2JNrqYsPmWX050bH08l97c5hmq1BYgE+rxXDreckWBy6YEKii
37AjTapPaGk0RSwpQcZPflJswh3pyQ9258qMFNrEzLxJnjB/mdZ3tjh7Ap6qaXuXCwwBJMEBdWdY
/F4TabsKSyPQhZ5+D7xDEo6h2v7aAETneA/hq/Fr1KlA6zIB0aThicDcSulOume07LCmFhzyWj80
jTi3TWnGEz5iTkWEl+Lw9QOeH76C6QWr0g0cZ3AY53pohUUZy1BMnSLrxdSngu3cAniAVmmOOHog
EK5UN1IK+JQt3m30R9QeMP6BJ/qpZa8ZQ/32rezb6vyRlh647QIXZId3JF3fEpBOrH1Q+viOqgLF
0k2tuahUTieIhFfdAAEyxcF6IDbArnoo4DL/PvN8OML7nsaf5gLRRcA57o0xrkXDYbZutOE8fP55
OBHiUPk+Xa4CInewzprhYvRTTD+LAV3CV4m+umjarwuDs6YUzLKoc7jzPGYVZjCJT6ltBtwVlrWQ
oGsAyQ9kLQTRXJg1XzKv0L6vtmXAchHIGahvzHtpqGXsc+SavSxB8qvW1Q77+PcOXCK1iODoOrC/
/D35fJXYWa2XmtPAA2mrNfyyCBqC1PcU9Sd2fPuY8BqJSROoY+CDF+M8sIusiGr3DLyA5+kqZ5y8
dMGVnew3RvJJmn2nZ9v1Q1SvmbwSlInMyW/SI1S0dR29NdYL5n4KD94Hmf7xwDRmae6BSsHswmRd
1lACzRYNpWUi607d+lgYpS/8xMquOwXFu1dll7TqTPZN/FpfF2bWmC8twdKyDK735GiJeuI54mf/
CWAp5SIBgaMfjGGIoJjL8r72qPzXZfKW8g5wmi3WKLiWslO3hB9KpNQM1Z+qYR+r7Mi6cd6Bkb8A
lqJTUyDR4xtiImEk46hFviwJXmIbzuvHkxzlIVP9A9Z8xYB5EHyAzU3zqSrpyjjgkBJT7rgawXOq
K8DKcuv92IK+MMzmV/HMVB5RXAq4BKOABMX5e+BfB25vb289jeE2acODVB011huUtmicceNfxPh9
rh8XYGdRx/5QPPshMoDnityAA1lArpJOQIcI04eOavGnjukYD0YEDkqT9lUPRs+/C6DXYk+LdvB7
BDPg2kZbr7tlWq214mDlhYMjitA6HXsJnsO2YAh/SvEApCjKBNDqm/4MSjXezaUJ1i3YgGDZOFs5
G1dt7SHaUbjAN8nLkAjzkjiX5hrjKpwPptyVgRFIC5ngD5C8ZJc/OyuwIDBGMTe4+5xwinWxuCER
VfcLJ8BFGZyqyKk/lcQPG5Q30KKBDg34gfk2OvfIA0EnhNBYnLZPtBGs3NB5hstzB60tvqV+jGDF
3V0SHphchGYoqkdnN7lO9dzBrWn5XSNX7qDdJPQAZ1dC54B5XC3uspkmJQe6B2gRu+bnTZMrfmXr
F/WNMyWGSiyKHFZCVcOzFIbv3m8Phx/b36LDvRkDQh0bJgf4JVKvhFhROxZQpeHg02+lkDLdE+NB
g3D1uiHD3nUymUG20xG9n+8HLV5lABSfVA9WDE8YbNTmWawpmzYev+WjH7p/CprTUWsHV1zIiKuU
OmCLFaJOq7WvfaMnGICoBAoPKM8NLWu3I9BhK8ziblig4/AhqToQhOR8e+uLnZ5vGbwDId3AlcM/
RhxDqzOFqDe3622NkJxlaZ9UXA0AGZBRdFJmuVqZWkTnbWsHcaApEB/ZLdSOaPmrUU5hNjIA432E
1uUY/F+Rh6ALfWOUTLXkSPmdy9CyDiCo4ZgmUp9uzgx6ygyoF8O7eBAK37ZVj2tfHM61WyLnXJmC
N+jApr0RkaPYgPXfup7jIvHbQ8HMxcWzAbvyA6La9F9Onme5nl++Z0GTD7vhoKxzncfjhbYljbgK
tN5SnOzSK+Ec/R+hFUxjz2s6xp4moFGGcIJXyXfL4o+ZAye+o6cmT4NIH1Bk8CFOmf5dEKKeGbPU
D0YMLf09g+erXg85vW8Pm4YoIIv9DxYyA4oVx+akicG1VJBUfpnBvI7Kqis2NoJoW+UbwxB3SaS4
c1kQtdF7Is25R4sTyuY950h1AVTrhX9vPdm89FxtctoLAP21AkezicWVQ6yB+UBmTo3csC3iBPZt
gs+KL4zLTr69UEpS+8YCej8aJZ0Yqj9XU36zVYeX4izhWc57xxJD7liESbDOxkDPZ3l3syqfBP1e
jWmKvIqzgwZB2G1r5J8VsknjKBIA5PcYHZgnqnw6hlFFbNRyzzdV9MxNs+GcqiveZRmrtTLeFqKn
9IWhRu5YVCiR/z65dZxdOEtYbFVnTd6sVc5Qc1oTGEVkryR0O9T7yL2RUMHgYZIEHIaevZg0kGUT
X+BqFYpV46NLXoP0KeGzxJccD6Id5Lkk0tCCkSkfesna7IfKtW48j4ye8RgjLM/Tk6CXtuhDlboW
mCjJba2rPYpUV3mOl0IzgxOhpDaZM5wNTZUtTN13OVWkSCI8aGlnkx9MSgEh7Oe1xf8w3DApRgpe
Afg5BeOIJbCod9iYgynZvHhgU9yNH8mhbTG/tt9Ak7w1vVj3whR2KRdPepGUE5hqsaIFle4JB06P
NZJtB9BUAR1fn7HY+RyPvd53ZxwG668qqzesOJGtv0D8Fxg0yBi45f9nX0K5GwbeDZ3UAqi70jEL
SpCQSuqmWuB3pKroUmyTSLlz35dlrQwFi50/dF6mQwtTU4cDSq3DUviXpDpyYH/9fP3wkbCfDCxv
a5FfXZVPAgNo1/a7Ax85ktMTtcK9/6ew7/BVd7GokITAb702XMwrd1F+mnynNuANjblvQg0ykC20
CWXH/Poi9xCXzafWmgiES+NoTQbB73U6TzCg2/+Dk48N0bng+qXykmGAeR4p8+YE0zqOcYq4ef/X
gQDMfDIg50eLcgN+R8dF7vwXkhxr9qOKpT4k4X1h8/xRTcnZI1MpeLvRzE2PmhOvRyIfh4Mw16h3
ol6zrKfWaZsRWC/35ccbvGgrIoNepeLR1arG2ytAAUuPsgYqZDclJiX9Sgah3q6r7DUwyEaKvXX+
WjPGfzP50rj/c5zUnLb1gHY7g8cBn/6SUGR5p+GWYEqsoryRWzZ/sP131priOGVpxgx4PoLyqDyG
YA86kV+JxCBSW9EtjOYXS9X19gzHUQg480A0ik1hessYWpOJh4QOOHcTf5Lo+M1Pul5WuE9gOZtp
g1mj3y5VXeo1IidzB/9xhNbF3SyAZEU5aEOlV4DuHtfP5g0YWBHLihj5t4WoZdJiLsCi70H1OH3v
+Wvp3NFKt+iOmYbXFKBmg5cCfX5iy6kudHZ4vFBdqDwO0rr2FN+xfRf646ImIWHcTMNhhH1EgmC8
EmGxCfT5ZY4mHZWgNoItw/Yiy3LgFvaPKThCXuKU13gCfI3voGYDq43aiu1gZvHejBhIYvwuPD9s
t7gNXoAukpYKx/C3ic+41BZcWKpnOQcGFLFTyvWXv6vqATBSpUItUOLjs5TWmd/14fLIq0JnR5v2
wGVYWf9SYOL9lDGHFLDeteI6aNYZHHqUJcq1FnEwsaUPSDZVNDgZp50RzrXF1z/yTYd7GTr6kF77
ffiAOjkDOdwn+0CwVUByNOBXRtjS0zHC1bR7uO8uviUjLSFvyJgjNMdcqPKop8ftbEVQTUi+cgkz
px+R5ZLQV9VdQufBH4aMM/Czj/kNdI2nw8sVUZ/KW5BUFNONce56NbQaDa1poRZbzDfBPVZCgDb8
7y1i3UBYjj2fjAXgXuFZdbpVov6SPi6sahUhYCwN6dzM0TTVhGRXTACnTfb7+fbWLI+sP2jtCg2m
w/Yhuh7Bl+lTXP7bod1Sa01TVDaTfh40fEZnlyWTyHhrf7R9u2fshM10Qy1j7nWplt59DScGWnwZ
HaaXCkhP7c4xIdAInmSTIEVoYtUHO0yeWtZjmNSUjNlCAt1O4587Ysv/0+Kj3l3seCRby620+aZx
qCRQ1zIPa2WQ3/9HbfvCeBbrNaT63ZBYVMBvCtQVlZqrNpHDA6juwJIbCSlunMh0oGkO+eP8S8h6
c/m4m1wSKM3U4IvM4CKTrS9eAn/SyRTwrpT3+byj+/EIBprVplFnXBYua552xvhEQmHEokLQJxym
xsARhq/6DMcGulMX4j+bnuISQlvZl0V6Pg9o4HYjoK2IDDoFKq49heY9JN41WibJWiVmjW+vHdK5
djXGxPIEAk42LjKxgHf59kn5nFd5L1/RPl9+2fvtAlpOBm2mLbenjSHiiwdN6lKPmqTubzZPcArQ
v9OGqpkU5XaK6cXVmy6LqH2vl3rgh/hU6UmB0P+tIDDMB78ysE88AcANzKQLXpUEmDL3BER0BNp+
GgrJIuGxdbIruRz66swCHFyg3baTlGHQ5qXCX/1y8WS9FfxEe6Clbr0/3Ho/yX3JDTuZ1YpoUHbW
VTVBUKCxUDaLRDnw9SsBfRNe/NtR8gm6SBlvp0H163liEVDIvT2pn4nPAUEFGC+N3of0bzzK6mxA
rTJMkP44Takjg48VG0WDyKsId1XeR+anBlBUWilrz4AV78x9Bh+VK5qbE+RJVSCvniWp42b8VHKs
IMLyhBylCjdFpiQn8kaQMQH3AGFv140ved6kby6+dhEm/DC3GMt5PFzp4i612TGWUDk3saVf+DMn
97XKzD9VGYPJcuUP606Qw09sgzw0FZyhE1Shk1q/OJFvefK9NsL7rlZH3xDBYp19v+SE3Pxx4HJP
BJ5xXVw97iKxQDZOK2BRYgk+kQCk3OdhthM2YBziVQvl4vpKxlJAQJK3zaPVJXWTm4rs0q8x3cql
7lhsxxuY1ZBGT6anYfcn+etOYTg3sMkYGaGH4apXCyg2Qz+DwRdWiBd973YIc+I7N89bIQvkl+ja
nc2jLn9UjhTYcfxDLyA2yrzUurphh6l2Owv7ydw6PlP3B0KOZOT25qvYnUzf86ZGBc0wuxHDYTG3
n02sOeuJaO4yRF/gPr3/q5l81RweG1rx4HDzMqLOFYQc8A+pQ9G/+TUpKe/CBy/s4QfE0WD+qb99
mLsSvBBfbpkQGdw9UL0iJohR4QcO85dqd2JbctFlA3B0Xoxbn6E8zDokemCdFREl3XTxPXC0Cljg
o+KmRuUm+t5rudI3kONVcEOT6mwPqHUCxiInSjhBt9ZaxE7rrGXVzKob4rg+STkkdCFQ2kWsm0P7
LKtRT1rYMQktgDLNjQkubu+1/GHjIiy7MmgAWWGvLA7ynfSdq2BbjTZlelopQGePwvglnOARfXoy
/js4qEpo8aiI4jKX8/IxmkoAIq34RXxdGTfP9t0t7pQUrnonEanxiM3oPL4o9GPcw9o6Cu/MEPn1
6Xde2R70XiYGOr4JjGPo5+0aMTc9bJtThGMrDmFPgDmHnPMzBnraOPvRO7EjYLRNhsnkb38EC5Ws
OnWoLYLO/8Ku5li8BzOVejmlFD2XLdn5L8BfMgLkiXzS+znQkSq3zPy09GWw58VmVJ1BVpxUZD3T
NyuXR2DkzcMH51xk70+pjAXg/6DARg9SjFl6M4vRF8OSCRrGciLPkvZHPuZZuupitabx7gxL9Ask
nE+4LJxQX6UnPF9gi+eg7GwkF4YAp37/MaJ2ae7mkacn9s7OI5bgmtUrbvvXqoCufI8RLfVzuMDE
+If3fxHQ4dgQuRm7ffBbQnfVvjLevnPKKVBJ0wYzwvYOVQDSZjZnuU76awMmttuijhDKuZ17DahN
CFW7q/oTj6suMtYnPowTNk0JRwVhPaSYtcXNE5/iJZX9RyxpNXS8vGRmhJ6P3lJabA29+ugsjeef
dJEgRwTg+JdaSsjAR/jOvH/wztMZ7cls4VT92C+CLP6kSV143oUyKWyQNPjU2YVxkzY4C4bo3VDO
l1BAlPesbCXu8dJHQ2N1rf4PAp+HCmfjwxftlIKgx/i4oQbplSM3agPZniSLBTPwZSo5B7UkFqQs
WwGDXYRIBCnPpz5wWP9/X7WXw0NBMZmU3FMyhdybCKgPCKebZXKi4kWpvBtqKvRWyo0s659elqJo
CdsAS1qo2/yafW0b63L7XH4cacH3V54MNrrHzsC2Mrb4aGdo++Lx+SsI38+3R3IxLg/JTvtKrdZL
Qz97fuMRIfxAaINs8nT1NRvBdHsVRiCfvWcjzQPAR5kje/xoQwWjXNpRLE6F5lrwCJn2g6Fi1ydZ
TafzETzNlH7SxoPdJ5TG5QBa7H0IxOQUWPdsUJnetVCd57sKlLUvq0f+SK3G9Wl2/On9TrLnrW6U
vLfWOOfpRIGozMLrAAbqiAnA3W/bLWi05CLc87ldGAvUAOpU7uaZqh4Wr25Ff26yLVnr9E/Y06N4
QKntEDckWTrxXUHamMEyIqQ5i9it8OslDfnoVF7Fmi2aXG5nDSpmGh2xQBBSGke+33rIPhMp2sJa
3RFDJf0L318zFh5hIZRK92Q1KjWuCikeQZXSJKkjFctlSEthUbBPnuXZXSxHPNrDpgK3pWtZl7ov
9wUsBb2X+x65Rw4Xddsr4rOTpMxyImM8LY78fip6j9p5VrtartQkVzGw/mFaASeojBfn3KA/wG/T
gEaQ4GrQ1Aa78FxfTLCyLj5jOC33hbY5GcbRqjomXOsXMJkISevM64q1JUxWUdQdOKbdz3R2pqD1
kqqluhgxSa14OXzL7TjtGNG11S4YJjxMtMYHmRIyoDofATj4fKeM06NiHhKKe2zFYf9imZcaXZ9q
8MM8Hk4cgM50gXywoppwTHzVGPedymUd5WCE8OqacBff9uVbLp1hpTuDS8hS/GJSfw/l09KA1nPx
qYFgE5dSmyyBUHF6RzPrBdyR/m4FbBD9ULYki/sqVRMJ6QORC6/Rn6nCli+PmoXbM23c6gPKqxis
9d0O2AAu7K3FciTQ5gxDMQD5CoXkm+ckmnGknHAIG25K7eQNzoDZ0IVgQsS5S8KHA5RPZHDtPDYE
DFT0awNXmDY+zBiuXEZ6LmRoHAInraADt9yHM/y+u+f/LP0QYY5LTWOQGDVkQKvZ2TwM3NK1v7+x
y548i3w02vD4shf2rlj8PnAEm479jvUrZFC5Fjw/aULDIGY0WCpfHGYXsKIPO/TlOrf1SqyngpzX
FjDxQjK7d910J1v11UfelLQ9RfwpPblZZdpDQR5NmiWp4/5Z2rdV09SVd0o/7wvxr7gCwkGkpX0i
iBcxXYCV0cl2YozeaH5b7FxgTSyFsOMexzweuj+iC+OzG2/EV0AWes7fgJcgMx3BAQMoHmdRmAcD
H/aeYfeYShKvhZI2o4uRJ2eTf7KrINP0QUd1WzFB+Jsd8Iq6z2m1x9vV2PPAAPV+SJZXqJCQ8wr/
5m7UacRB3LGvpVCjWDuF0Ukwad6DNp5gy5FQWXnFPAXr59psxcTZexPCT1K/Q1VHxEMhdUE3Ftyn
NuVmi8dXIMF4cz28VlAt8EQ+SCb11h/kpn4pFqGj/OVSqT5Si61wlrTu6oaGW3QBK8FDKoTTWJNt
rNYxI6oCI6rR6AYMtIYeSo8pl6DyH4MpNvclkzAYUFRnoBojCNkO40PS7BtiKZlv6ejbWgr72VLj
GWZwz93oRDF9YidRQq6k+Bj9tJ6lqcLr1hnkJLKEASjUjZGlC/HpEy6l/ZuXlKNFBCRauunlrbGo
/nc3EddpYIsvJKNsqziIFbrpQ/i2JnRJNnLQa+E8aJ0hEO+buAPkSHtEtjP63r6dqLqCO3RCs13m
k5FgrBceoyt5BwFZTCBO1HUh1Gz341ZhQIcWUzM/qmIncFoFZOeERmsRydtO+hYk9zJEJcOo+Y0h
5nP6PexoAxmOqJ4t3pHbya8pE1Koif0AOSLPlR+vj2TwMufKLVXdb6e7DO1TIoDjLSEr3CXkOdQH
aCmXLW338xUjQrkK5CaNnB9os16/1JL/VVGATBry2yzxvqpwuxqNw7ZqrgJmJpvEIlR7xxXJxBPD
9Zwmjp9lDBfSlUSXh7cUcjkeym5n6q3LuEM4poKj6w8UCE7Vb5PJJCCfPDXqFO2sWMCNvrtNYyvZ
5+nxcPmMaiAVA4zeLYq7jRCyClQvarSw+J/OG8QA0HMQhGo1KLtJlaWBV89IwjrwIIMLAO6aqS1D
ZmY1tcGEoxmghxsTYqfEMSG901DlR49S9D4kasrCM8MWNJWdi7kHDoBW+bzHBupfTdUndYieVfBl
5jMPSCufg135qXOkcareL9u75iqmmVzlREBMkkBR7CcOKmCnaTPHx9L4E57C2Kyr2JZK+aeDt+60
Jg0X1O5H6JccKttkbRJCIPImn/7ELsOuFCgjEGsFHw4fJ1S2dZ75q52+iSC+KylWwM+ilRIbgZ+Z
8pzn6Lo+TsvlQL8bFIKR8xvvmewYSIQkPK6IbNPYjT6ecukIdFazVRK0DZi29U7hrLLT6HZTp5nU
7VZBK5H8eLn9FeVBpRfwjAncw8ZVZ99NBOQmqdvzUBInXRr0J9ygylO/PcOzbaXFFNEsr6MdXQrf
w5RDotSV7ERyuITaXpXkvCUpHgfF4QHFBzJZWUU52QEdwqzg29uCHpziTzDosxl/uMWQdM081K3W
ji8jTbqyRnhbHoH4fBEJiMLI3OIrEp6yK5ZxUNzN2vueGnx88sy1CTPj1Ireg8VWG7zAb0UllQFc
IZdDT2Opfph96txepNMmxqUoOsez55Ggg2TOIHBXngQhjXGTCkmzH4C3Tdqd62xG621xlP8na9NJ
K2oqK9vsNf9u1/2rBkcdqnlBCrSIT1PrTR626V5rrKLyp7IUXj1daqR0lrnSxVu1v6Q0U657g7SG
C0vC3tlMjrK9saMcuUbjoYP89PQT4YiV6fyxByzjLj3uH2ooYhzrgQcvU7zlizvUZDraEO7LGbl5
Zowjw7Gv7XPAUHg6Y7lulv8/f2raGNlFRf04AMF5YBVHiqkgG83GbqNujEBsqo9DfJnpt1z3pLhV
BBQEDYqCz6MMlw8hEPUakm4AKcNHSqoZfLVZlRB0xXzfiu6bh2LVcXLcz4KHUHStvzoBMD7TCcB7
3O55uaJKftpe2iElMZFCAxwgPp80AHAo1HA67eVYJn/nwfal8VboZQAjZrTfwnfaGKp13JWAtSZV
qqUzj71zwdrLsCSu+lB7uP3sES7PftbsZzqCdmT8l1oLrg8AVujh17vreWxAwbhq9HqvCeLnYomE
lfF9z37aZKUi0/cq8UNmTIYSc4mU9YQf0Q5qQv4XZh1nhR0uHkFvMSd0JPPJ/OrZaBw4dTpAVveT
WSWVoqL13EfV9L9xd6QQ1wplBWoqVz2wSmlgK63obH2OILArI2TmILOiuREXhsTgRlausJeaIexj
mNOJq5AmurzsshMknWvFef35ZucV0p1w2Zgst/upxN72GEeOqaBLpSE9ij4uawAvBF6uJpRJ/JXq
S8lEPAjpYFdHWPXQqXKkw1Uc2MCKCjaOJcxT4eo6GgY5dy03PTLpeWH8ltMUGsGLHI6Bp+RkhW4P
deslDwt+Wn/sM+Ri086ljbVu6xOdcSKrrLlSVzHP1+n9YHUMw0OP6UNeV3jvgqfjqDZ6asMMsQtU
3EyRQQJGyCkGMmAyw8HAFt/u6CaNzuBqSt4wFWogLmOg+gS233gx9rrXqRHrgWGSZfHbcd5dtWIj
9eE+nZ4YU8V1Sx9I/h6wKAhMiJ41zPIJxb0HZH8qbhi6pRw9IWmveg6+xgMqVmjxZcuvg5/eUmYk
eJQyxnxKwI6tLorG/lzz8NBhp5i6F19Bpkra7I6v5eoL111Us1k5CjFb01X74rU1GAbDcZBcZ2hr
j2XYsCzQEW+2PoJ5c3mjOsF6ClYJUjzbVd3wxBRO9iJDnR2wtuNmLx8ahDSQu3lc8dZrdLW7DIY8
0Qy5a6Zr0tZlvqZ+upJarFCUSrVNgewiC/ShqcWp1sDXFjhkEgyS9d7sgjCAx79WvWqvSP2Ild6q
jMk6Q4WiJS6bKD3RKw2/IgR/OoF5xcQ6xLZfdcV4oFHoyImKMGjv8mfX/OcevyO2+LkYvz5qyJH6
j7x8EWKYE3tjdUzFMhQiklvzoX2KyKNLKqmo1W9+LcAPQFvkMdCaICpqlMZnVSGpHiTJu1iDn5Pt
ERch1e6AfH1g1BhVdfOhPai0zCM62j2m1qs+SNrXrSYbPNHST8KCUXR7Y45Lhq4wbE3pInjG13ZH
RX/lHt5FedZztH6yKe7AsP7KqXLbchuKPWnSEBp7c51rtnvEdthmejtXLBgPsJzcaO6xyBkDcvV/
MGB6xLkGkbmAb0DkE54uNidCbokK+tkeOqKih6rZjPq6MD8jn3Qp8S+bvPH+8l58TYvMnqeflsD5
cmO3d8VeX9X8NjtbbU+vD9Ui4XndgFalZpuL+PG0RQQRQpKMKEYqEz6UWbSa9pFmihdk1mvq3ch1
QmliWmG+t9T0LhYfecx5qQfgkg7s6Z4bBP9nV5pb2851mw8c1JiV9KBxDIsUWgEmjuek/td5fNjG
bUWdQ+6TfzY8I+PUgZZn8ILxs3Arh+oZn1c6FiQUso8guvq7jJwMmXSlwVC6tKZr9nwQUSwoySkp
JZxr7JwMtPPxqVEkv+BE+N8TxwIXrkHKR09VQ/nsyvXOJt8iWNv35xqVwyfy4DULlaNkjvGLY3xT
mhZ0JvIQAdxMJOnb5uukAHXQ5IA8XK70+FjmXSSFxsk3jVGx3BE81c3x0tce+urFivnjuQWegRsF
hRw4A/zSkd5Dpxno6Nv5b13nBSg5Qjkl55DX1MZN9kmhKQADtukp3YfM1uW+KORWOJp/5fsKkxJG
x+RMx9B0yR5D+xIwhxi4ZBUVKEZiJdr8m9M54TIfZTWrxHkeoNAl9EyNJulUemyNgyr8sLdAJKNy
UR7FN1/IJmZFEOQUC7zhDM7Q44K5r4/rC+9Mayh8uPn83I0FSzMRq6zbvBP8+O7bm5ACKN+E2o5x
79rqb/9k0dvZQVUaddEePdRgDG2PmSDINBWqucv4F0rP5fdo32dBBaToJk2dsCmohcs4D9yK92se
+Q1DVA7ePhACR/pLyB1PzXmZWbYhXD9RwQz5HO7FI1JEWSpH0MycWJJMYubkd8lDKbBjxJV98/7G
aYAm649962DBSKdiIf27OQqDbyCkiIx//b5mMinAO77HKnfAZ79as0s59VwPIbcnEsJ2JtgbsKd0
XMx0sMrhDX6PoCSUDtsUtGleLUXZwUCVaypfdFTkxTmOiYopRGsIJHlaDGqmmgnQXSH3YHENN0PK
34hEYXmg/ZXlPMLd6Ne+/o2J3mxReLwBlFZw8UiTncyL7nL0NmhItBQruPvDhPI4f00e4XmY/Ypq
rI8OWKQVX0YQl+VMprV7ZS14puPuMe6ToHKapT9wFGi+7ZS1zGOV5yPVHepcqlXn7qaLu0uUhdtX
/l92axU8zFlyl3vUkqvK7KpgYWujZ04b3aZvlumzq/65df1hDnjUmVMVv0pqfdlrT7fVcQ276KjM
Gyh3A9uj4v9bDY98KHBVN54YwT2vbmhEYmKzkoVB+xoxhUYv15KHA0GVZF0vKwqrYbi3NdOdldUX
vPPtpg/oolO6m5RvP/4EbU/y2aOsJ0cMzWnoN9oh+1hs966+f6YcFeYRHfhFb80LCjDC/T7a8ult
dmM1p1OEN1JMsyTKxHs+inidX5Xc2yJvYux/NuT5NzeJPwg+aMUN4POe6zWluXC8iAHJo0f5x9RO
Dr55rSRahn0wCNfAuJ8iA+oBa01Rpt45NQ8mPqHUUv11lrMwy+LEHIhp1mTFfukPWsPDPxzWIedm
IhesAnQINRBRYwfxa4bHLxt1jSgli7sXaiNfMJuzk6IOnXFrIQkeXvgej1HqrTzjAa9t3I4zDlQ0
/iz8rPMD/7I+WCQVvSUmxGFn5hskd/SvhMPiXEHPefVcMLFCikq1eCOaPy11QeKSgLD0upEGp2yX
MKBnzI3/ghtQXKY8k4i46mqUirR4ZARjqMh1kCQs5lqa0Se1x0APCsuijr+dorqHFbeAKCqy3S9D
qorz7g7VEo+nQMXX4HItOEShxshkyIw5hDMoW9XqCuTRA+AvJK175OYdsALRhUwX15f094VrbInm
7/XD9cUF4oAYd9CFBYPlg4fuZAkZP8nsQgoCGCtxq3yZjwrgiy+ZR1PKCbOJBNP2xbZiWoeq+EBR
QPx+yPQXKz3wADvFJJo6ANlAvvxJOO+IX5RTUuZxYEvcWV+MK8KjlnMqoY2je9b47t4w8t79/N/1
LWtvfXTpXQQBZmQnjYYYIobKZILhm3tOLQLcuhLiMvkI64z7Q0bz82A9XoVEOrYTh6yU9WSu/uxr
AxjClwBv0Qxd0yvPda7DW5XveS8tcuijTvErgm/VgvFgeY8gw+PgnUHOoEz+cCC87zvJt59VmCVB
Fksxod7KnIP6svpV0aLzp88PioBgIdU4OQV2voY9MQQJj1X81Xj+D1zataPRFuWOqekG99mvxMBW
KFJBJSWQhkNxDJZqp7yzfxG8Po/Mlp8LjfwiitSdAFKxy+oshEHiQ+m2gTwDXNhqYhx2lEexnEmh
L+FbZrf5v8ve+tgB+8CgYDEEChO9RGFHXwGCYfI8tH4I0LHaMISHMyoTuLsSOLElYVVGFRYGDwH/
aljHHhvvhfplTgnIp+Tegp5Cg6hz05qZlqXEVfh6mJS1pAS/dqysFjDDc4FjTaEAdh32e+jpFxWZ
RhbKmVguZTW1LScp8um2cGM/EuOIUwpN4iCVZ9fWrSl51f3oUo1o0v0jD+WfU6M1+E+xsAVxs+Mu
4qiTct55Me/zeGD4jpsn96Wt+n0RUy09JeOU+zVKJgc4Kj5wolhNa7CO2fDZERf9kTZfxtKo5Hj8
wogzDDlHGKGF9VQexmKyd/hRZrylUqyxwnPTZEAozckXBNItXMofS8YTnLacpOPk5LKX3ZU2G5UI
sKhc35KO2mpCBZWja2SfzDESEtjI+Dk0upE3aG/LOsqMeQoRhqJMj4mVP/sUO2lf4+t7tRpsC9M/
Zs5qBSi/ZdrV4q4ZXN7CCom1g8OnD/blvrXhncisW7EEEEbmf4Dyw7fYsE4L2H/WUtNMlVumy4/D
iLxCkuq25k3k5x+PEKXZ+3uP6fsA63vaR24WJ+469LkxXfD6ZfXzgTocm/PMDgxip3sExlY0YcK8
whE/0xRoiT+YANXo85mRWQxqU6MaAs+g/jGPhAQjy52NtStNbZrXWsQS2Tv+N5IaSsrbum6q31p0
9aJiS4xynQ/degyX8yzWByCrB9jHjnjFvgiFI28RQZy2KZCrZSpznhr+RUEe3LSeR3F0zPnwH5sO
MEkGXfq03BtYjs6BAHryXIenArs1ig6PNtT/tjqiLmG1gKRKjWYHXQ0WqS89t7TNfBPjzbOehuRU
17Z1qdhXjuME6f9JxeyldIYN49tQlOuAhscjXqbOd7gZImlnmclbbMQSf5kALPAIDdXtVQ+RfHQf
0T8DScGyd8KQ3IR/dDZgFB+ydER8OAcfBmRPz6hQj3AYdGwDBM0DKRC90NR4s/6HeigbSeT5AzEe
RMcE41LkMH1mfCe3AJphmnHKyYynR4Qms1Tec8BVOkz59KYXOKJAGSApWlkJ9M91DDx8pQU3GnzJ
/5429RuejIAofQzM17C5enndMR3ELXIIFRFlHokNmPHP2Bfh5YSSOexTz17R3O1sjmYJd2z6SuL1
o9wjkq2QkbyJj87PNMPSxo/heRsU3Z0ZRuPU7r+BbShItwQ73aDY+FZorEUJX4FTEWRNELOw+sVn
JhvYYcPEYaEJ/DAQ/F1AVYYo+AW36YvCP2wTZ4Jz9UXOXQr6K1e2UOJyln9VEgew/wtIIEidd+y5
F89k/NGF8yT7Tu7ZiHlbdabBY7dV3cxiZzh0YfPa2S38IIZMJ/a+ACJ1SqluskGKLkR9PaykoHmD
uMV59WVlXU9hK9ACECN1qsWf8bNRM8iE8b5R3ddCKExFxTlGB1yG0UQdBBn7/JrwSNB7DxHX+DxC
7VgpzyIcaosNka7+wUhI8TsFZpvqg0dqNtoGgoB70YloUwwj87/q17qDK79LmLt+sKrN46468WD9
Qb/YbDeXmtD1H0gmhFvyZryKgfe9DSRI2Fj/wRtISa7XNWogbI1zOgX6/D5vekjV2wch8c6DhAuK
Hty8fOoWbQLvURYohesPDb3ZU/57VvA7rXthSnDwNG3MeN57D2oEW8ZK57+GnRTSNjZdLqUeGZZn
f2ZKayrTG7zLQjmmjB8lxTZq5nIiASearMmDQqRKjSBmTLTUSDpFHm2X64+NIg91FZDkpEhZd98z
q0oO/5vEW3j6j2uJqIvReYS9P3vXERtVRM0zbxGBWdObaIZbBFyx3YsnPv75F3r8EUyWlxOAfVWo
aeCrUaRgaYH9NqEEmmlfcncl1nX6Iv/piqXR1kM1HOEFBdWCwOPWbi4KLK/bgRxgvDL0P7aVEY3L
BIn0z9b911umK+HZn4r6kqk2l45ao4fJalswpkMQZQbhDpmRA01k14kdlFcyq3+5uFeW4KJqdlQo
uWKUIBNOxu8Bb6gUaFV4wtTXlK+RiyuBxlValP5v1x1nynoAw0GsrZK4op/OHmRKd4+IttWDb6/i
JFssgUqPSxNpfiMCr2pMrktYYtcNs0Q9Xx/wBjM0L8oUw5WBWmOWJDwp2h03tNr6xcyd8FuIVhxq
j13DXolcKbc81YgUXNFykHgICB1lqP6BCf7g+lQMNchLGeBJzhR76AXeVnS/VEZmCG4uZyPijg4B
+Ncdlkbq58YoKXdfVdM6nHJV2zXqbwW8DGq2ZbWXnI6C9M/GmCrBifxlirXXO1GGU7YIwF/krd4k
t3xHuBcOY5FFfX5kWgUGfaRxUzE88+Q44hqqT07hESSOOlNHFH3zghVfj15jmhGvMr45cbMae6tC
axKMMtwHVxrm0BH9zirwZCu01Tvxe0mjINf+kiWMs70o6lKZBoFNHxA9UqapAyRiLOMLylU6ntMh
hvGF3cbpaBQq1iLRxC1KduyyU+mlwSNeAy4jwxM0TjkY8vAmrPKW5QtjKBOvF2ocrPci2dLZfIun
esC/SF0DBXI4b+3f6oXgAJ/3apSLvxR8fy251xOt20KFwWMHUK1JQiXYLjsPzXIIsjlbJyUzPWlk
xCfcyVSkGch4c9QTzQ9dkO6pPLM1DQMvegdrvzVPaE9qLnrJ6QpwaiME0OXc+5yAr9119G2C+pM2
ZH4xH5QXWz9zzFsSSpslfDlIJ+X4EI0vJoDrhBMviokw91em7j7YEWTw/JqZnlqctsdpKKNXVM+X
X9uBoHQpNP7bFBEAjSX3+IoshmJR3us4wtKjlZWMNh791yWIFYaP/HjqhbwYWLN6Hv2gQ9gsV24/
qgE0RjhynRP0i1MbCgJPH2U6R13jQWJH3hqSX4ABdqWuuu8+ND9tud0Ieu/zm2OVSqmiaZ3MbUFh
IaUNkL/XuuhF1e3j3cCgPanBbJfr4PtfbnxR/ZWr5M50T9+kzPCorUj6mGWoJ8B8zMmtn1Y54jsF
7omdGYnLYeWEeD+ZaFHfrUIUjQKZAWBvEsC79+DbWIm3DAXa7hhywftWfzNbXiXMIMRPGuKzNEfP
1Pzze3YDdoO74noOYdOefV1JK0ODUBmX0wzjXeZJhOMyH2R95sqgE+6YPEMC6P6ox0mL7VjqoTP0
Ptx3S+w5k1PAbKtwXTGZIgLx5eyde61peS3Wh3vLmQ3N8P7p/Y9KFzjRcLPlPKBDp+9flbzqXgQX
u6NLVQRI5BiY8fB/OTa1zq+9P3dQ903KLDzIvn++cnaWvvQVoGBuAvUUdmcnO+93v4cL9hWzh6WU
3xWXzf12sYQkMhjL2hJDDZ2qCle82XfOVaJLG+ppmj+/8O2XChjxAxMhjVN7D2UrEmu6PtPr5K/e
MwVF5IR9cz+GcMM4/21bOoTg5sdod+clfVlNziUG1KS2tY9GQgPvnv9kKLVHKAfAicoVvh6+eRmB
QV9kMthS79uuCHKH21GH1z3XAA4gdOV8SyDlpk0bhzzGgBh5/X/9+5Cp99mJ44LpI3IvawAe3U+M
9g8a4lzkwhOicT1ZbF8yAMd0hKYsgtIZqjHgh/vE+sYKvZU1Gj43Y2dLbDYoSb/1cSEttH54+UcS
gADmOsBmocC3SgtlzmfeFLs5Yd4ERWORDNyFjCrRhh/5SUAb2S1K1iY7TafHqSI5DdOuW5is3MfQ
GP/YZIL4EHwNqvCGAoEvrZJwVnxcMvAfKLQ8cC8sAv5ATPphdoXBnG5eJtP9hT+iIvmfcpLr5Gmj
D+IxLIWldfmsEbVCfMSTQEYbz7wThSxlQaPEkULpnFmryswdco+qUcdlBjXvmMSNjo6M/Jc/br3D
zmabAocplkYEDJP76niyLohPp03NJtIpTv4Cgo9aN/e8TrJOH6VoNeVh0exzJ+UWVJjhGrUAWOYq
5sqUNVSDbbwJjIPHUZoe6l3HMyVQi+HCbKE1Q4lqURugBHz9WiBw7ag4RuSUkelpqOOnMBkQ6nsC
DZxL980zlEDH1yo22hLzQMa3bZI6vAyyu5VAFJpWSVVzMr9kWyqmR7Zu+ljq5mQyTlhSSMVPyUlX
yAE4m8lIe5ltC/MuDgtosuYbinaxkTwL36itL6SpfmFTaKI5NipvoLi9sF3tTMZhp4k58tjC5qE/
Qrvg0UNhCaxm8cLinSRCmYHO2eXOC9XZtDQ3ouRuQWxu/f1HooH3QcLqwhaExyrMXymb4hqgfHZg
k2saEYXNxpbsOZRPaOxwhCtIQq78qcqFjH+1wm4B0wtGoE0Co+q4E5r6yU6dhgheUtn7KcRoSCpw
ygyhzOzUocH7H+T5lx5zhQz1igzeEv7AWFdJkSn47SRE0aewPkrObj/uD2OYk2+NOuWGoBlZtb1B
g3UhA6LhiC7PqhPy6pxmTO8jnvSKDxl8uoj8cExrl7nz7buH3yAj2dOkr4gTzJyu84rQd6barq7k
MawZJ+EnqEq4qFmMJ/GirIbjLplswbn8cdSyJztoePSco2lDYLfNk2nyjg8E9/oH0OBjmbGXL5nb
5CJZ4Cmk450qNOS3/SgC8wFpd+gPESlZfn5BJb5rKTQZBszrzck0tbfUlQ3kTrL9zQyLuk47GaAl
S1BchYYg6MP1i6VkBRukdvwTnCUDcLqv252IN3s2X8EljmIfb7VKoZrkH+r1iSPZmUdl7yUhUMox
zb63Npxr0iD0CkP6+VsTTZgrcx/KNMokzSAhbnpl9kFGUWN+EMjC55RMr+K8cZ7GIaB6N2oOZAqX
R4WrR0qAhrSB1giVnv2ifn0h6HgkTkNel67ZZlPHC2k+WHjBkjhOhoznL+d0ch4LDMTzzDKn12xp
Zg3HboGnKwdd8Kpz/B2Mm5DKcVa6hkSmK0aFqIKxBJT7FyPpUrcdntDzTQ96Tg/fXrv9Lcz31txS
oNhNbwCq56k7Ytn9FHKfeZHmEXOyxyHKiRx10b/f+edEEEN4jSENjgahWMTIioUBoLgbT5+AV0+n
r7HLZewZbmNi3hfvnbKZ/G+Udl8WwDsbcpIWGa7j6DYm7DlNNIFfZ3H7JCIslJ5IsYurBbNVp0Yk
E1d7Fw2OSbWJt6spkl9tdEcsJp8LISb6w3FtMlZKD7bFaEQYwjrLdP/l80g6VH3Dyf+4Za+yH8W8
3yt6s9AvV3+Ovub8g2/uSSCHx0A4d+5MlTgJw260BJkgne80qMwrGxcOKDMJxPS87vlJ0hltVvIb
D+waQXCXn/auefg9lwPLBqh4uTMNPS/nzOZXTBK6ZN/ExFJ4VaGxgALc2G19omeP1B/DxP4C3Udv
E4jZq6H3XGLORluhzUkKBe5ZZ/xnckuSriVO1b+D2+8n3f8z5iKR+Enzk9NnCijBmAnaFz3TlcMi
Ju9XPT8ntx2PpmX5CSFJD55yn6bHfrtamz10sv6Qom5HN4GcpGsO8T/jylTBOeu3/zM1cHqsquLz
ALrZFZaM7D68u1NGqtU/EOmpDYIEgXmLd4dweUgxXX2JB7MbGXLiJtBDVocqCYREqpMnJ7a2kEi0
o6mShE6qqZWVxEiwNbr718t9t9eiKdgDaSS6GBiOdzyx+6vmns2TJFwK+aOiCvumHU3xdrfWkChe
B8EHHiOiukPM1WNdiggpX/bobRe38ByxSUBOSxwBeGooTCmXN+2pJxcqpFQB/qPtSzYI99CbjIV5
jmlAu/kz7IMThLOC9uKRO0q3j61siMGOoHwI8Mtew8m3ozmluckiyafPnGKAy4S+ABDF1Mz+Wko0
LmASif0MdhfftmHVSUxIiz6npnwItPJ3ZItBQUgU/642azu8dN25c81zmFhFqldJnNUY3ahTlCb1
W4cacwgxBlwXwusVnL6gtNNrXbK2LIq6fJAaN8p2NyM6vYPCTXkxNNtQPcA12G4fWHSRdkOT0//H
+QSLWANo7Ys2gh2syI1o6rqgt5mVyxPUwmrNVAA47qlGLKlKGeHMzabLTiy4/27mU1to002hfUXE
RYpvSkl0QjMpq6n4c05oUJW9M6uzifr0Q8B6kIUBfxoM4vaO8LQY9y8rlmgviF0BEiWHYDE4h7xu
Zbv6N37n83DvR/pmohLvfKnstHPidEwTL3LfdLQUfeeyVTHZ+/KoJ8qy3l/DEyK2lY4iqvrt9KYm
TPSugyACOwL08h8BlFNvdPTPiruGevMsNSdvG6QjVV5O6EBxoKDoaYRD018cp9vT4JC7QHqVu+uL
1Nc6vh6zX+crXjpsqu/5t8y6pYMICmY4xA3/uDO7RGXc3BnD4j9fUr2/QSiy3+3eFPDTgOQdSdXv
4SF9sCJ0ashKUMT1tXU0Mfy0zaPEgFzwv5ALZlyVf2lc0k0q7GEz+GbQUyeEwSXuODozP21CjQA6
iKeudI6Y4xTp9qwHZ4tD+JOUIQcGakZgrz8VBTXLHo6s7eGHAZ/UwgSL4Jgyi+TtQW4O1cgv8ooB
vu1MWe1KE3mL9RrN4Y/fwH8by8oFoZsiTACNUbVnRvtdMk2w6UcO2LB6ls76BIMHgzIZo+0SwdG5
lxNeh9/yUnj9GQILeTM3ZkfS9JzFsBpEhIbTl1Tks8x83wBOFyeNfPD4nnJ03hFtcahbtYsUDaB5
KoDab4k8+H6Pg06ijZeL3WY4iPwebasFPc0lMd3YLe/ibCLETR9LbqERkPoUX2zo/jz7UiKKVdsq
2FGYYoAgcFmm2PIqxX7lnPZ33MeprDD1P7E2kKOWrHHNchb11XcB7R1Fu2Q++trS7/OHTUuxW+0D
MnBTGWxE9O4WyuS4sIsmpZwjr8uLcVzp1GpnKnRtTYrJJ8NLjLo5+NkZWv2rsysF4t3v7/leisWF
8anLAIXSeS9U042eh4iRmKd11oovgO8Bm/ItsCzsO/YIuKI4SRYbtU2KCwQt5eNkvBe762m5h57q
tnNR5v96Df0CoLvGaYVUMb1Hz6By1J6f/GqhA/2tGDGUGrbimmSxpvqO+rKLBBvTiofOIUeZrpbQ
JJJlkrTB/xviDYKOIPkOPIf/gCQkm0MbPgvuxJttNj0qlYbAzJOpMudzcfEhIWZYf0cVbNuCmqeD
0j0lcGs5kta/g7q2qL1CXwSiJvbHPJ66Rt8DMmuuf78B8sdeJB8is6m1t1T0jh1ZMwDumLYk2YYA
Q18BA1Se+HXb5PB+tOaDYsRDv22EATnxTIvYMkA/2etpAd80gG5CVNjk7Pz/x/Dg2H4JSD6oAPh0
5iEQ5SGTokoHo2Q8WVG3xHJst1drO4vIxaFEnEx7/Zio8RFhY1mevgEA2ZhRhSzP9wfuIGHlU62W
U2cVm7QBSBcNv8Ni+2wJQmTu4kZMjrXLQgROC9LpLt7ufBZo9/oKBVSra+c34hUPLYTf80EZBmSb
fOxbxcDjdy5H6m7H6Uwsabv9ihhBGiHUjO32hDajh8UBFnZly/SZj+sAm0I7vRaa8cfb8cPsp97u
oadQwD3rHWn+YmeIxgS8nnDdkaVeGHvusysiEoE9UmFEUEDdrmlpPsKty8ro+fQN/hkd3VoQxX+N
xLh4xEs6wOA1m9GqQO6HEN8JyscdxYJccyVSAArkYjPOmQZekk4557LO7rNdDIUdAzrVbwYKUuI8
TtmPqMGn2TeFYOF6DYaksZLfNWCTDKmsFWCjm/3mHQ0YN0DEF1BXzaIaGtDliLz1wgYz6sb+zL/X
WNufpGIwtlhx8GPU3uGIAZDs3jDE4pyrhUmq1QtQh+OJ0NQHrP9HDPfDm+cD1+rm/scpPH1OmVSJ
GKGMb4AqOkq6OkI5tNnP2K0djp4PXs9mlkWi5Efq1Qo0qJoOiBlTti/1uwFjOXKRPHZ9Kl/io54V
KedK9O4GYgwLoKwB4qAhcvOJ/6z9MZVHtwl7FcphQGCIbzBw6TmsjrC9z2dR53ICUarpFoFTccEQ
4a5RKTIxSyBCrjOydS/tiNgK/84t8j7iRrPPnK3YgMUPGtHf/WmbZfGGYopSj+pciqi6F1rEkkdB
93V4EI8Tt9OqiT6CSj5pn/abpvi7HspIO/oVV9oA4I4AFMFgeH6yMHuEmFZ7JEWTyRCrIqrCtLw7
ApkChcbtDIlVQvPNNYpwFDnwnykJVzFlATFjI+AjnTa+HXAwK8yzHFwFKqtlCFptrTEFzVKxwM7S
iAn+YfqM55KMTB+eilldjiGe6MsyP5E8gRLyCSSlpRPZX807ypl+eoa3XfVhMw6pd0ls7pZ/R8z7
LLC72lECId2SAI5DmHxXtYWMq3zyIustG/XMIj0hOX5ATtJvRw0ktPBHM6fOj/IzrP1tDFyjqSWr
/ywLA9uwPd/WRR2woW0Uswu2WuMzJ6eKNFSyrs11heLSN0DJJOOJF3JFEjkftcTNsQUEmwsonwkr
8njJQI7rvfQWaCeqkk+zQ8OgII182ZELaIY+95UXz7pOjetTL8UtpDNR35aNd9Gr5ChIZCAw+KNM
jk/Ne2/usqY/qRVgpQzoF9Ef30ZkZlo4H+HOf2BlnWs4b9h9NFEhRCRhtRyWZ0/P95x2N9t7w28r
tnBQeArZusFj0hB2CkcJMRDjfFyp49zNt5n8NeVJoiTfLghYyX62q74wOqb3ZHWEJMlEiTO73M3P
j5e623wywCpxh9X5kn15wfRHpWL/3ZAEwJZMzTe3fTISlSYCZQBAOpHlOSQDzTRIXnrgMtnNo3VB
MG4zWY60qF43n126loIxY5gQ23tNxXz9NRFOgsxoNorfVCTlt79wOo5t05Bi2VEJ9g6y1TfgUj+x
Kz+6qHc2UqUK1h0hA2K0pNCeHo7iUiiBMCJIOkx9wac5AUtmtqCOWhOzV35AkDhQbBsXKwTxNx6S
wL3m9QpkI/2m1XDEA3S4i2XfAreHcfRLugnxfXR80+7GBT3z4DwaHS8Tnnr9Quzd7ZQWwkXzlCrq
LZdyqDSREbjemhP61GG1+MGq+2ASK/qvKNhfJCPXDdQLr0dQYcvu65hioCP5SOZrk6SyR5ye08fo
g97WMoRaNOEjoCNhRHciLRdtEHplWIGPGEIkUldOkFs/npj3ExohTdOmWiamcqjOo6KD6J1He7Sf
x1vXAP59mtmEIEE3i+F0oF+ZsxiRzUmZC/UVTpW5SrgMEl4ppFSkwEqJSoysPpA15zEr9x9suvqF
6IcQBzMqltYcs848SKP9alkCyYLz3iBS0l0/iDZIQ4zi2kTy88Z81NPF5S1tTC9FHWOIgx2F7iH/
ljU4ZmPAP0INGPbSfpwkDINtkYk6x95kPLSae4wmpml0GY1NedXbLuNWKItdiILZziZlTylvCz4M
I6gwVCiAowDH6ThVNGwiCMHnh2rb3LbYH7DSEZZB+WVEHEudjn1xGsyQe5GlLZyYMtuHgEo4snma
6O1fuzZxW4lb0bFqlXDY04yU4JQYVFCgFqCy2Iohn07A99CLblWTKlzA1SOh7PLFvLMU58nfrHg3
14Js9s/n8e3rZiqGQx+oyekMf//Y/WGe++R5bOGMaWEhPrcv2pSnpxNZVb1OxogrlcEvlnZWCeat
AtFQztyBtsLZSjgZXyKtF2tZ6ntyjHYO0oIS+PKt28TmVViRF/+yBr6PoQwXetO0+HIeUJLIFE8l
CJW8ZO1WmbuQnRSf+8PnJnORTfoPpp/Yhf8HxP7rG4ZTy9K4HHWKQ2Dap6ePea0efdIDkpektOH7
UBfRbjKJ0AmrPEVXJz2TPvkXL1nTWMgYF02aUaXTAF5e6+WNS6KkQbcfw28g59BvvdDXydD+c/9t
9qTmTAP975mZegA3CpsygoxUb5UygS/MnbdFh6bF4kc9T65O2p5VfzR4Rm3xKO5JgH4uNEY7IdMR
sjgfeQJrbM4nKcVKvVDhLA03EBMlGdDsdX8WXI0OeB5BA6vLY62p6OJD/lQeMAdkFFp2VoRy3Jts
XD802yMWJeQdVPtDjrVhFfsyJukbRNnakM+cvh1NVGoyZh5xJ+QrsrDqJkxXenC1q0w3h9SxUULW
ZIii2rCbh1IkVLrJfCpfhIOfr8PnOxS6SVQq8nJ8EJ4McmuEiyG5sku5e66bdcq+g2ZZBgMfwQWQ
mQ6vmmWNm2+1j+RjNCzdfVSzZhlWBL5zVKMIwQp6Ho0PeybKRc8dGMDHst3qkdECM6GZ23HJKVnV
XTtpKbA3PKA+V3Vi/kMKYmqAiIuCBkkYmWfm0MpxSG+ThZcvvxY+1Gd9a8wFpTXan11uJf8m82jU
aQ28JsGsKOEtuk5ZSuHQwJ/blXWidGAE48UPxeqtZCDoSCERB2RRKo2gZF4VQ07TJFToq/BOIDn3
UWSRhdyGVW58LAAiGAtdrfBmE+8BcNCQtRRo5OT0zaHnGIm4po9Fxc5Q4vlAmk9ixPPBV1xx4uwB
cZG30r6X01uaquqdZUTmvJeoNMcQJpbD8Dt1XvVJnwjK26WZ4iqKuEzFzw5JNUTPpDEig/vrIrLD
EROJZh8LXjKw2A+OVwQ9vQdm9oezu9ExLxaKu2P+fjaHjU037KyxYJv7m453S4sM5hOK7cRO4upc
Dt8cow0mf1Hc/k1bHDHCmxsFUi1FlP3D1c8l4O7hKASXKE3jkCO4Fh9bXctdqvU5tEHI++uKcvd0
+guvdp0P5qGVlpN54BId1Y3n/XLfNgtJ8rbCcmDKzwIJ1CRW5JQK8L+iFjurmgoWJGbSphu4vWxw
2mCr3h8bb1FypIoQ5GoIS1UXSwa87Brn/zL5sZdZAs121kglCqFgnYmq1NY6L3KpCKwPSl8sPGjn
NUg9/bZpC9M3D+BPF+zVrfqf+4+5fsQje+pEzmF6uNiru5yfExRn/jnxcx8uDPPLx/WYo4GYWg77
9RhqtbniOsFkMd93KMiOfWKdwy9P2Pl8HkjrIQei73RFp2aNnrkn4iN1OgcoG5qHluLOrLZR9GTX
xpskRiJJavyViFBsrxFNH0V4nulgM5u4fB8vrWIRcwYVdbtGl5x0lMiLgZH27xl/Kv5MrIgC0Cr9
nut47xJSn2IgfM9xvy2hKBhLqGF6JXaXGXRt606atEr9hufb/djzyUmUsWjhFJVrdiWyDretj5ey
2kFeYxywy6uWAtj88KwylOnCvuOoF2xLFkSNCl5+DgpjkdpcZkXVKCBLLYn95GMqoak9p6q0OnJs
ygtVs5Sz/nhR5xpd/ga+VnH3pzstC7HT0wPYibBJnZPibzKdqB1jH6BPn9nvfAYdF6lnVUBlLgdQ
r7VRICEr+Gzr4y0XesetwydstSSuFH2eEUZztX0IOKQuB5wY1idx5I8ZvYsW3LwoJI7AQqYF7xJ6
33pWBLsE92Ps2dlypbGgGmnmV3pnsWCIm2zfqD+6U84Jv7+8Tf7K/QS6xy6fMw1Y9ABpLNPS0qVf
ojy+S+njuNheku6ryUPOQLd4R5XUvOBHaX//IvqcflIiDT0gtTUGzXjHs6bbzf24LNEgdCEDLBvW
unPVKVH4t7/IULWDh9UlCVHcXIdUdlb4AdgxCyylaTLzBn4hJK2zQFtW8WED4H/jZJHGxlyDZ6i4
XPIIoY2YFQJNmS/ivhwLrpCBQgNeV0xFUvIV1ZuXa5bYEN75wLt9jkSaOQxrXvBgdzT3nX+I0qG0
5TSlpTKY9J7bNFerc1YkCPH9Rr8xTsfhP8Pc/BtEDwifTQ7v+8LMJgsK8fed/XvcwSpDl8OwTRH9
3wDzzXKNHnXnzRJZvFr0AjMwmLOE+E54EOCp3f8T3mMFVhgiF5JlhEUA31ioHtOjbgsWDkl5uE1G
4/QgX+0k17zisM6yX9m7DoilXSzKRDBjkp2HKAD0oetpqsjzBytkRJl8gKqIocGKDVNfcRoE4Pv/
koXy6yqxTrS4rKfyS/cLJLdQ+PnKCtE84uGoAifGjSLY1Z7amPv1CtlXC8o1/DWpaQ5ytGVu+e1J
1gmkeu0I6ZBuGD8zW+QAp6VXtjy/giTPchGYeES8LuT7yiCHs0npaDbOIaGTuHLUv0eP8ofOT8Ov
581Ik0BNs4CMiKzMx5+AqcjI0JLDuOMU13RdxcctuCERAU5y0VObQ0h9LRSbe53gl95L21A/C2FA
LjQKmJMa674aHXFBaAzB4xSoY5BKLPRV/dpYgH70VKf0ZMpT1KQ+713O+vlCnaS9QpM4TwlUcV45
PFQTI6I0Tk0Dvvnl8JaDKa8VZYs60pgllkVcmXV2q48mlW03AxxpkwEIcGhZvMGbVwAiPwjBDd/z
h76LsiNKgijHkxNeNSEo6h7mMwow07zwMjKQ6LGdWGbVTnzJN/MLm5b+1BBMze836hduJKXDS+C3
WSbJ6lfHZpzJnmMGl5TYNHLJTl6O5XI/lJ4dnziPDlUh5DDq5mfepeu9u650ijU6I9ahcN9jdj2J
jJobMsQnSIEboOCbfTjnu1NlkcVpioLjITDIEK1sTbSnNP9i2tVca7vY/Hxl8o7L7vOl3ceS3qr6
K00LdFz7HbpxFI6iiKvsJyoPSbyP5qza/U207IC0kApKqHmVv9ZkiDXGw/qhb90Q+2w0P1Pw1v7M
BiGnMVXAlDniZaVZxe00Qs7i2jld/TCag6NMkfKXJMV2S6byH+uvjhFH1iR+2+gkmF3Mws7LF/px
awLsr5sQWyVfMbBTyKllXnmJfuYry8zFa7RbnD1mrWf45dV6J1Gyho0hm4vWKmGLg3yAP3e9X1md
gboi6nCBs5nSNUvwtOIfnhgW4hqo1a8Q5U8LUhxkq725/mi4Og70YQX/z5e3+XgYgkFmT5HJcOGc
IVyDSwBi+cFtihV6z+mkSubz1eq2kI/jfpJcdtipGBEyKos9IK5MA9sE4kjoJhXo1oWdRBhP9nXH
kGm/dJ0icDKgF4Qxhc9rXvVjgx0tJnAUB9fxJibqkKaAux+KEl5iGW0B3XJKa1Hc1eozfwupOzoT
gIK8XMIx1bGG36SkzVzCGRoxmAuVu4rQSf+osD63eHeL7FXH8I/QQt3Z5UmnBMMo52AIPzFvIe+Y
5PBRtwGZzGM+Anb2HdStJ68zX4MKR33RO3Zymulvw4C+wC0QLXuuqMdewUDPvWd8h2zDpAcSGrm5
ril9s98ZSzdJvqf//W7b5i8Dfq/36A3g+PFB2WCJgHy4RDPIYkJz0zqn5CqjJb6G51IyAW4InCYi
o3zCmZ4gLXS/8xREKw4cW44goH5c+hQ2PgyECH6jMnu1l/MoRlXB1N3BkQ5gmolZ2vuf9jRuQ+qt
prOmAU1N98ZwjA8SbPEUzkFsgFy3ZLdV0yqPSJYEg9UmhkC4+M+T0riU67dII/OmcHq2PYunQDxa
I/PY+Osc2VAMnv1eIAhoLSQifbaC8RXBARVk5aP4KDK8UmTE0WXc722gAIkc1ny+VkvuAXChisCd
TOuVL3dYtvOhQdNoccuWXam85wetASqOA4aiGh1GjKsfA2gzmA8GvFWMB3ZveQqKSbrwCbK0At0y
gyLybHb0rAkj8c9qYdmJFei8kUqgP9R+BxHHcjasRzgVS9+li6XM2NI5N7OFX1lUDSdqgV536cZ/
QobSrat0+ogd7o6Es1DLzefryjotMlDmFX7aIM9ARZTgpTQN6kgHyu0/s4/3djhsIluqSMUeAUa5
5QisRP6ehQIqsiBjzJAsdCaddbqaUTcEGvnMpAJe3EuQIDmDbEHYkacrcsilPd/0pacW3G/3QDbn
TYmfdwYhtsCcoFAF+y5w2pp6sSzEKCrDDVuW6QlMHvSswGM74VwDlawynj2icMBRjNwIBJJaEcZ3
V28aC0KounO2KIs0IbglNXgYCgp9o/AgwFhHIA8ZRnhJWz6RwrxuvKI7Q5qh8cjxhrEOG0HO1xbe
mujit/fDkT3ISy77ExuaaLGadUXgMqR8yfAxNpetKrGN724OjvUlsf0fHm8LqSHhxqDo6QG5v09Z
9fqu1eOfeleAFSBi+nNvnbUAtiGwyWf8DIk40OcgRZRdGp1fl28xsL7M9Yt4z7ddBKzXq73zDo7O
XA0e7oWn9yF0YLY5l7t3W/dkqBvkJH91iSwWQd7Zsamcwbsx4LaDNLyoc4khUaeflZ6WkFmOQnk2
+toeoXlhGhdbUCVZXQpJvp/iOkO620aci11aqGBgFiBxDP7WV/MUhfXQQoXPt2DTtT8F9O/qB4K7
T0IZlX6r5X04aYDxLVrQBWv9+/r/H21HLDZEsYZEvh1HTbyiaj0eVtsGYSVwXInl7fmSY8KayzXI
ZP9NlsObEEmRaXKk1FG6QOH/ZcdAOHRIqJcg4EBAvYkRFQfIb9xqeY7e+EOxiQcVCEUDHzpwdUgK
5SjUMoNFfxCMg8wdRhNZRu4Pln4XQ2sbaSJb9Ujhr2A/yIT17OawXO1ENvoXkH05RYd5E8UHQDcb
jU2uZwd4rs9z8lnZMKAhxpXEF8ZGGY7Q3wBVtmuz4GjfK5T/04Zn2hSD8aDX731fAIGjEaWOLAzX
XKnNdeCn1Jjbq0WeXyhPhT5lAIMpkkC/exvYYmEdnLFfi6l9u7s3VoA9HucQifQiIwi1JHz8n1R1
Iur/YolqV5X8NIcaabRzLysxoOeMfC6qcA3gsqqwfu0w/H1VOb3QUqpOV+bxaxHntYqpN/9eanTi
628lG+yjQjhqzbMcjec9LcMyKr4tSf1T22rwzjKeuWe4GiXXGCoehl/d2OKm60N55/snG+c89+DK
JycjjhaLTJZ//lqxaoGy4IjcoVmWGuSdlL2GtCK+///9NrXGhsAvIPue6bQYKkGMfMf9372AFtnB
PXHKyEYp25s6L2h0bXHbqZX2ils+VTtP1lsvUb2AZMPpU+78944kCjkwlQFEsUvAsp3NBIFwW0sm
l5/I2yaZbZQ5n+NuheHn2PkdCz2efvKIGHeYxjOW/WsR68IsozP+20R8izoXN41+awK7P6q7lrbl
fkWtck8VtSpZby5ITm57dUHj+GdOyS9ug+upxeZgiwWcU1LEBeIDbTi8mN2L4ZzNmJzAFDBNWqMw
IJ8TE2dK/lC18fW2VceJJ8hvM0JWxmXRfmicg2CsXp4u7eco1YMZWfHePY+hHAiCx3w5w4Z1Y8+I
fAYZw+DmUeYoTqvfdnCbQ4CqdN+vI9IbotiYGo8U9U89g3v2pB7Dhv9nRZRy0i1mVHZWcK9eRV4u
8utee21awu/Oc1b0NP3mNfOPTXQTjC0fMWHKuxor7eaLypTNP8/VfXNIl+nmhPSH2McNPILQAH39
QLz8kHDb/3FHJRFRlOkAGmlxq7KSIC4ZcDHGe6tqOxU6KfRuYkkRRLMTwtg20ZTNy6bjyppdxv3r
cVnMa5whWU3fdd7hgiOU+/7BGPF1q+gNTgNCBY2Z6w9gaVZRrkovDn/9vVQsBlOuexVp/4aQprbT
I7bulpEYVMydPNLwYtN45ZUygksvpHuJaf1LA/xFYUJjwtrrtrPKW9lSn2WbHtgXGOmj3kUwR1q2
17G3v1Xr/r7515leu2k7FA+D2qzSbrS0qg9ZNjT2S6dgomon3za19BKtNdGUpgh7CUZ9tAc/jkWb
abz3wZFmdE1j3tJh4H5idPFFs2gmcwhcwzL2kZzkkhzsN/+HmGOQSDYzQcZHkVYEH6oaMd2U/Zt/
kzcRWTqrTJEhermypL2Y5ihwKn+XthyHtFMZqn5MNC7Dnh3EztX2Bdgwdy7wTL89kbXyXGwrqcJX
DN8DD2RW1If1X/S8fJpWHIWNISoanvFhe9zH/R2eHnjK0MktoNwKVbUYwWM4z19puBf+2TDKprCV
zHND0VSE3FMmmwhAgOv329TTcFXXyg7PJiz/ZVQ0ZmiVAyft3ISzIRWoXaOO598271+3uPjU4qxr
LJ7AcMebZujVkHSM9kodQBM8UeHc6J6Q7vunOdbNkdYHusluMNLVoMnyOVFE5dt6yL15HGr+HMYP
lfNZy5Iho8nPQMDsuq19pjA99J4uUVJVhiN2UYIVMsUSWagjIaT2EX19ZT77Mjt5MEZ1wNmfluP5
Blv5Ql32slnGHAXHaHuUj0yPd5dZMaDbGje0V6YgEBrorDVPltVYJeu4C02auroa0NFEDwuvh7cr
yEd1vBSCVFcqaa8yT0EKuRxGnHeyObSbY75IspYbHaRw2lBJiKimof+lMV6RiG0ccby9akJNigTQ
BBTkzFgm+oMo0L38FF2lRYgGf4X5q7+NEQEaVzPV9USDDrnv97xWXnxgUIUTQjLMa6jTXDZokuz0
PBdB7z8QEv3hahCPKNiXCScspmDM3vjgMIjnQruses2dKIWIqIJx54F0CXuAyZqA1grE9puwzWWN
pvgkJb3C92Dk5ImiHbkJrYKkI0JfPlaY1PWN9ZPxkFuCO6Dw+B4+AecNtAymR09Rg6QMOGjVAYeu
Ad8gNhhDs2ge+GKgAlldTQbliIl8ppDiecoTCzdfxqodwjJbvzyalPR/saKK6mrusCZsB307nh8/
PkSvhK0DARdhKy803KNhXSsjoi8GLBjqguD5Je3uX1vbmlH6bGLwHzKoGg6Lrabk9fHsV/SQ+6K5
uBQ2TVY+LqMmAJtGUOn1ZNr4jAg3dQR7O5RR0J7H5JHcP9k7Jf1Vqct4iSM6wknohFKJOVvd81wL
Si4zylQMN88AYv+rPu3aRBQvgJ00tYfO5DFoiQG3BahI6MZ4ubsxnbZkYpv9FwiiB4uwnA/G+Z9Q
9ISe93dcznk4l+MAL5Msf/icmu7SlSl0ECHLu/jbP8fHR0roEZGVTk+MzsrvXsxlGn5kcvKT3W1C
ZDLAEFPrOYYZK6VGLjnmkuLYuS0sWyb5Cljy0dC9eDAr+ZQOawj9q+h3oe0vQslq7EBmOAdrFYUI
Qkw2EUUrU9wJJGEfNensApeL1iywI7OzUxBvj5Va2iTXG6AjmbA43lJW6NhiVUSL/ppiwz3Gnngf
4TwU8uMsWLxQx5io6ZvQJqB7+ZzZ8HF3c/9VK5F2U2XZcVvRtxVpS+3GRxi4+fyF5BeeMLSn3cN/
9YpfG+unZq//YzFMgH3CAweSLOYVZdLi2XKuvubN7mF4wlmnS8tA5y2+7cadUt+USGn3eAG9OBu0
i9JOehy+X39WaVu0pYKI1b29cj9MWI10yGgZc+a0sSqSB/27TnL41ztGkHRbaFSE6d2Ne59H7rDD
B1bVGMpmltS3PKQ+CCfgZEukU933nr4JfmefGnmh9ZDDIB20DIuzy9pnp5avELHBupicnU+ZXYbI
bdAogg/HFiAaGppJFKgER32nfcmnSQILV4M74Xy3b2/ivhNBXeeKV8aRrJDvkq7ZEZoUyAKYfoW9
ypA4fJTx5EC72NNpizIZWjNKqvNfdUfuSq4nz2wLD8JzQKm4Rw/rGmyHRpfvlhkyAKlPVhN0xYJU
0qPlGE2LVtwRCn5Tv7r1fW5u5K0bfHVSGrq/Cp3WKC0UTTZ76IOMtJ1OOGCnhK8LdFWDeS6I1Z3M
jUnK16InzVt86VnNK+GC+lXdsfqw1x87R3xdHKXKN+LxK9ZwY3mnTAyMHixVj2NXKL3mNCwj23ZB
/pG7z5voWWUxVKUTiZe4gbJB0DqmBMi/1yDYytzLXj947zMD6rzQOUgkHdr7v8Vhts1TCeQz5S3p
bRI3gT3HjQ5MLOBewhy+kymK9iG2fHA1w6IX22RXeurJIdShWJ78fwJheoYaftKhjCLvaRVXVDNk
YzRCk7bmP9EJRjr8oOq/JmBCIBD5EFN+r62UJvBsMj3NnScJ/8NwCDeVqyNYK2tly3ykZYy510XP
Ach/EpSJLHzRc03Afcy2lrTGcBftaKYMSCGKmFrPDrOsTJtLobiya12nSe+ebVjou2RaHS5+dSzA
xk8uW7uh2fay5t8e0TdxXuO46YoWV1YHycYfeaDrKQ+AlEvalk4xwLQ1f2xYhpxb99H1D3jEYlnX
iD1pcxqQlB0A5Em7PcmLnRoMRkUGdtdPxCtn1RfAd03xGbEBlP+IhW//TjEAprMGCw9hCffzEaO3
YZ2cNuBuG4LQvgEcU/59j22KrOudwPOvjpbW85nLeFsql/u3PCk8yLVx8j9VkjN5hSkzzdS8ybuR
OLN6UgAmmU+e4b7qvWo5ovpkDR839o5mgHy/W+zueoOXOQF346a962YksH/3/JFKJaVT2HMiKbo/
gPRjeHt8FmoXeBzH///aCtBdtg62ZVmxbOzWa4UDLbzxNj9NOTZPzOHusJTSylUsJ+x7N+e/6tAY
V2914nFX10TKFVTd5j51xcIbjcMs+m5HGnqofL5AMPpa7/nH69O0g7WfldobU2VyIYbcsnoWyLqi
fQxC6m44vWoFFA897nlFivRQOdv7uIz3ukluW/PWFZdYnl1fi/TbXe9mQOLzXPUuxQmDvrIVSe1/
fSel5Qt+B4Fr1XeSbn0GOz4d6JpicH9tSKxLMklc8BcavAPF1eDRauGojjOWaL2R9IIYqwdyuB6q
tz1DIrrkrO4pYBKtGK6O9nF8UqzsnDmn/IijKKbHd/K+L7W2KYXMiCbx66teFJPozfBzdblOW//0
YgazPQeeItoVuaGo79SPAaJR4pbi0PrMnvQ93AslmUp1Gb0SZbsG0UKH8aRug0m9x/NA757Upt9b
fXqIXF9KcxdqFznkl/qRxTFETdcJUiU7XSl4UodU5EvIlojKC41L18HZ/YZrvFjWsu1od9htZwhz
aCsVadLOgF2Ex4xLVt5amk60wib+RCF+tQC0dNediKZQT5f0T5PvW6JbHj1Z/UP3ddzydiEMDztP
44c5jsh2iv0UbPLV089f6y+pkC3hkFZzk1JgKMsW1oH3AqnThBlhDJszbvToDHaI3S9Jgxdglwa7
b3Fzt9n4WYRQH5T3AHbke1Dxn9QFee6mrby1nr8xt+KQC1ZTwIsWyGBSJoMiomun+1palJ8A0ciA
pwbZPLf5rPembXsOeYpG2hzxL7ZEfsFFAcnyb58OS9CmmJstqLY2vIpwrtv2Mlwb657K0a6juQ9m
8Yxf2LwzYo1GrSBMQ4d4wYGWaKb02BzFX38pKUWektn9roxGxBMjJC8nqHa+nol6c1Is4clPyMU8
tQRDo7RBOuaO7vexYUCEkEWy2EWQ+t5tqo9rvd5/9EJv011wnfIQ25DWxEOtmFOU81aPOK/yKsEl
w2kZjSMI9Qf3/UNEREa/hMlY6ZDnqTO4xly32SF51vAMtBX7j3YoZddvWaQXob8yQy3JSYWXOKtm
EaRBMxtDz8ugepMN03W5gSrE8XdnT4IvB5vWPu0q/dgqvKrxLkFOa+VCVr2mC1b8UqEY0xE0l83d
AXVp/1RJPCJC4ycX3roMhWf83fvr+I8GLZll27PeIauAcvVmnpJo4NCFVZIBgB03jNj7VGgzXI67
xk3NHQjwbQHgXAGqmhN+CxmsOAdcl5/CXzYemA4Hrnnbr8r4NBEDhBcqYwT+HLYkHCL0AgRtgECF
zXaBqBlWfokvOOWe07XeuE6yhI+HdPVrFyUFJG/cGTr/anMhFArEaPMHjM/Zrpv7ymDrgTK8MlsB
wq8xTWaR8MtMkt8bF+Ehpx7w5WTa9BC14zJ9plxCPLMo3SKExyxOHs9I+osDiH+vLkn2QLfRd0qn
BrVFRigo4rBc5pc56ZvoeDaYxrGprl/bjmcBV7Y2wjceBcdnUmL+U3HUz661ugWSZRClzNkpMwtE
fagpzSBxYUNyl58PAORAH0c2fDeF4N6gq+zHwfjrmlDmG9E8K5z6UXqKdIVao830cw/o3rLc2Gud
mQPmFsQypf3XU0kjIpgIWB2OhAWUOLqLoeAOYij9KRHzww0Plh8iGN101nvekAJ89vUQ20Tj2Nkr
bnPMLjsRybLaX2Sdq9Ln1+5usqlW6DB+T66dcnZhWRpgzCFKnATmyObzWwfmJGWbWq3+agPRUdT8
VM7BmVIVwYwLkmitS5APD/LeJ4Ql/D+0EbftWr5BFU48WqzgsWw73Ht/cdP0f5RucYgkjNdGnNlu
JpEvM4BhsEdQG4q+bTQDyxgxe7qDI88l8w6HPYBi62Q/7qJvZq38CnJ/qGdubqOebUEehGqw7jOc
U71seIMNW7nLP8J8Gq5KCI2Uss/sZVs37LfCPOVudqUeJQaB0xzbdYw1TadvMrEpt2vZa18NlRls
9HUIu1ZIjjmRcB7EsTB7AUyYVUSLtZdqSTLYnmtip0JgwMuxG2lvWAcs0muCgPvSZvuG0ooShTM/
X6pXxMdItBYjLhJIT5iHIYX+V+YGVTVvMhKs5mSsj78Z009eo1f7D2YAHB1Xj3GrBb6zxJ1TMqA1
oVnelS4xQTMjvTPItSwlE4cgHYsXjato7X3i+h9cTTRUPH5av5d8pOm2HQPgkfIQsSaNBQzVKg9u
pqj0UXnmbqN5qw+0PvTnGJ+ks0PJnmGNwN8s/AsFKMomYNfo6/b2M6J0ADikfT/vwcYqTGDMKbDA
D9njCx3sI8wbIFNq7PBYp04EshYNv6wJT0m8PewyYsL3BJ0xLW2HhPQ4WRncakjvkyINJsWCIpR5
d5vQkHGjdCPNi9lQBgYgfdDrgo2W7uwP9ubvOmrvYth4Q/tciPzighY99R7nV5eo/XyALdkf2UXI
Ag2YpnkVretRmjfMqjCFpoyHL/31bAJ9dP4qn3q/nFeksw4suUw/J99nMzve5csu2paUwvL1InDb
1ShslRsnuN1YofUvBdL56JgBqXxiZs0YQQrnDtaxNzaUylLg4bReZTX5D90AAQzCkfOhRKfimtNL
1Kg2gr3DMdaMdUBpUaUFRvwnInYeLB993MdFn8MaftncxzHLUpI21lbxhbCZFssSJT7kMBoxJbd2
2GwXdPuC0g10IQVQph2l8XIyowUaUe8CU8xDLoW/CcH85F0NNA0ib3uMTpAUpg38RFg+SI0863Ov
h8o6HqUrsUb8B9fr/IhZOMqg8SrWCVk29jMXAgmMr00D6b5gwqSLeIngm5RsvpkI7bYkwFPBJ+E9
1NY5ynhtF2VgokLw+65cyyi91Jn288fimHjfMOS6/yhtK18dLLXCMOwV2N9gdo6pmJDCOV6Ysmrh
Me7Ut0+EwbXoF7RcvaoNicI4hwORzerFkTqbwMJ+86qYEUoG6gX4sXlSRuNK6XElKsC9ThbHz7ga
qF4nVYyIBIsYsncj1lWMQt+LUXLl8PoF5XkW5/7bPSIiZB/OvixGXHb+Oftm9UoIpo5M0IEU1FQr
h/f6aNjL8GaiCxkYojwryLxJ7EWVt7RPfbgy/Kgxh+/5P1BLsIDr/sG1SdOsTtfDcYIo4NwTxXU0
meUAdlyDrYsJrZTpBbidTnIFu8bJIBwNgyzgElYdgskdjpxR6pfvnv91q6Ia4Uycrpj+txfKdKnm
CLhYz4qWG+FPDrpXgQbG4zFFLBU+oMe3NZDZJnNd36/CISbssLK74rUDuDeiZQN/iUEJxrGllO0y
jmGEyrbVsqY6vBG2wXILCuwjHTgUBmZmzHVKCppAQfDCDlGvGZoQTWAEDjP+lZDvHyl8K8GEzWNi
nncC3vFdAKs6l97rdujuyt0iGDmkm/3JrZXUTgTGm65Px4N4rZHj8NPeXPnmuiXe3fUq7jsrQePc
A/M1SsXfBg8DTwY2YkJ0bpipbDijuhWutoU7+WOIcSkoyp1uJ8DA3FbZuSOTTAnUXq+pbcpELomB
9Lp37Hu8azJ8H2Hry8D+LCm9BA4z8o6hoQRZ/45ZDD1MZmwRIPKe9dkUQ5mNN98SfsfGERxmCUXx
CTEKqc3jJ9nk/olx+QRNCZ9ajSPVUQEKoB17UKaKjja5GeqRjVR2zh03WrAu76sNbRcGtQFsKC1N
Lq1SKFDzD8d+gd1K0S3EiLBLS/F1hWLBH2RAKMWqb6QVzioOJTxr6WcR0zDgYZThR1Gc3PUZavoF
Rh6f0I57UoQBI9o6GR+tWMx2bw/CTZl2H/yTlSxudB/Pg66+irdRZRFn4fTE+WYyrfh4/RVCRDeW
UQZYnKgkgK7uLw1fI5ebmSzLgZG12YC3tPkDDtnQDc3hNoLYEuwjOw3xXd/NWcHeGDRGCyERwcsh
B0B/yN4s3BqQtNHE+BuSi3k8WHVChiJiQ67sbBQ49E+TPqzUFXfzukhWcqJTy8/6ThMOsWRWhe8M
LYBOSa35R41wWmT0UciGdXN9jIsnhbMNslCVXhQ3SQmkU0JUkJYvCUsVsHeHPwOavqKYfRNPkQC6
O0wvcKVBVL+fxFABkSiWu55/QftK4h41CXFQ6XsWL6bkQaSalg9JWvKSuNipgOVzBsDFn/cASzsB
HMcqWTPmMSSTQs3F3vciKPCVnyaJUwT52eA/PC42/5PfRUvi8nHUyX91P6IPvPB6GXN1G3Y5x72n
icgKPZjiCgtutHm0pwC0UkeTWNQyrrutiv1YpPZ+uaDleDhKHeMWsq7htBdHcED829P0+Es0Tpje
UzemaIg30moaciazlYTjM6DX2yp6urhgOKRNQzol8dJ8rVTSX2tsXVawgIzNCXAhi9B8Hqilr/jr
oai5MOv5l5SbKorYC5MfXxZJg7nR4hV1MEH9WiqjuzCbjjayJ/FhxFzfIFr7rYgSjxRwjBccsXfZ
FU5C818N52CjrT97JcdbyWz36zHvnlgbrXwtjiGSEn+YZ6hpWHLdoilzjrEFDKa4w++/X1ClU7pl
/UiafBCUSjzNCBg8N0VCdKYzjwgZjqSkb+viNEcW7iO11ADi7xPlU3ZKiG84c2Mr/EgU0cN35KGq
bZzy1U7/Ow3qzpM9xbfVqnF3nNM1WHpfNMRoyKEw/UAauWa+oyC0nUFSREsvRZdxq3dto29TGkuw
SS7l1tjbuD2dRb9E6WwcQnEWE6v6kMkzjyY9JRICSMRZ5Bf4C6B7VSHpmJcXgaMjVYgtgXh6QGHP
fpKYTriar87RqpFZm5eZVZh73XGDWCSEw5skteIu20Zy/h8TBizJqt7WtyOHm8cwDSeOuWrgKchn
my/u3EyimCL7LuUusOjv/X1ZnPKmUTqRrgDohVRbn7dJvvGqpqtUaQD2p4clhvCVv+pU6tGeN9Fh
HADjs6v3T7GuB199x5RNAMoreqFaWMiYUdOGtS6paxswwGt9ZHtaUR5noxRUGbx9oGT/0EaCEMzQ
nMHh+njSsG4gRgwb19gzXSVbZB03FRz+If/MPZ6mN0A1pKJ6HwC+NZyEYLll7tjA5Cnn3S/XO5Ec
dj5F5mCdV3jKxl/zotvEkhxvSsJwLR7EkgBrnj99YQpVSkoKIcp1W27gQYq1msBEkIAdnEi0oH9D
W2ySVxrsqGTa3hfNIXUVHKBM7rXW2/KgGS5UUcX6xVp3BpOQsCdB0PzOvN0/u4ZJoLp4Mi0rZ/fq
nzAaZ2+ZwD4u3q9GYjXHzC3H1E3Hzw7tlJQKgS/v3AV3sc8vUus8dpvSPt1fj66cgXXDvHFzfXYR
SPC44f0/tY0M+unFBHVqjPeonqdVdcTWW2oqw6wWgVPVxnPp1GYwT4OwriRcuK9SoARbDbF5mZoe
5PIZzOJObFjonf9LS3Wvro+jD+rt6OPEv1pxiX/4PfWH4zRKSxwGCSWY8fSB11rB9Bcvw/aduPfI
uJGKTB4sPst6xDy+41Lf9w7dJ81X3dtBdY+m3MG8C9M7Rtsu4jzCSEqH5Xit15PlG5c5rhH+6SbT
F3ZgFj3a9r7VdFWjcqYZpZNL4dHvNfeCX1VkXvyDtP72Ex4MWqCHFY/Qlm3e/uLigpVUhKCKAjsY
8/SArfd9PSnKazuPsIAv57I7JY+IvWCkhQ9M9znYq4zgCnQkl4a+LEW1FvF6QjV6crbYdWHx/Lsk
Ahxj+sDx4cfTMcpjj1voCVi14rAY+u6tuZIj23Z13mYSecVdDE+JGr+dpFYb2npbb73AhjCkHEjU
0Wf9gP0gPpLGkwCd7eQFrj153JExNMccprI39uT2lKBtiJviejqGjo/9O87smcp+J/izqNv9/dVu
vGJyn0yx21n1iRcShbxXs/nCXn1RitgRg6G3zUthBJXtdfgaFiJBtQIRCsJGgGCbImvHYJpsj+s9
GVO7AQWNY7+n5zgaV1++6nRTaBug76dkBM/z4j/2quC5RY5WsjOn+bgFuOf8NzwTSN5sI22Mriqo
kbqO1aHZDOimvTWYdVjly4FOc8OEo5rKiXFgrRACyoIjW03RwfAG+YaM9AKZGE6iXckcfwkc2zDM
1T71TYlIHbIqutCeCEkv3tQ/AGokjrjyiZu3ilNLpuU7GvKklJwJ3LO59L9laCLQek7zZH7J/6/t
FtR4SZaNmWbooTX9X81iG1/bCAxj4OySZmXNX4NuijNax75gx3P++VY8wd8m2HFc9smZ/YCTIGUc
Hp4EALXmobmb/cLzQsvEIJJ/ukoLYMy+6vf5c7jZjDp9P3A+LQeewD+NussG1/0wqquV8CvCQjDN
LEb0x6Lho5t+wgjB25/dzNcAcWC+SaUiSGBlzzj3i031zF+dnHb6Iz4r3Lymq7M8vt7YfF5eA0mz
p9qqE12c3iuN7kaajAX4FkZaMTUXiQ8WifqrnB5bq5FoaLFxYmvCuRgj2XVcIZyUd5XNE29G1luB
4QSg0EbQEs26LC61gpxFx2YvhEbHuPSSzopcBrxCFMvxfhe9g8+LYXlzHqObg2mEFKZ6a7+YoYxN
sypaMQrJuTTnVOz2qy2IBVVEk38z2wrGD8eu8cZDajHBJaJ8u2D3Mv5085CPJKK1X2nD9PcEm76J
1dYWEtR1hHPeflx+pDAjhEQgDzXck/Ak2WqrYGyMHKQRCI2VOugXjyraeYy8zxVzx6AwgBZDela+
wdfBZeGVaXgMRb5iyba+3DaWv2/5W7JaJ21UIEHoHWUdDWRM9mMg7ZgIendVTAR3EGeGooQblcK3
ajx61YGkvee974TOuvqVz6nK01e054NEuJMhS+i3R4ep0c2sysWr1cXJXqB+78gsdAxS7wGPJDfa
W7HTDU+F3eWOA+mSxk/XirpC0ghdXofCkK7QxWfFGkrIu78sdoQ1UD2mIhPJ0dIGX+PfikRIOsp1
dj80xIKXKv1IxSXm9gfJvryepbeiqr/a4j81B/WbnDfVsuYto5nA8eLA7udbZAPxEzctbN2B/wxc
BXPIH4F5EJtoq98BkNkr4y0CCoTkIR2ySaB70d5DRmZqtWWUB58qu8VVdty3zalRaBP4jsAqKnLw
asALtfzt8btd3z00mXD+IXyTj5U1UrMkkSdZIfNzvYwapAM5enKfMFX282WDiO1SRVyH+GsKjvIQ
esJ8EKnHIliy/WSXJLsdiPbL5bRELQhRXGCEM9QaI7r68yEdheOF3o19KKhC55NxKsRX/SiGb9P1
D9SukAnk+PIPZrsrJA7cA9l61M5A9fK42fyBOpVuKm0f/sqjwDACzmPBn97nPiXxAF8E/JeObOda
EkYKmdMfR3OVu5VK33VEOhobiTOP+CWHIpKDwXjB+mOTaUc0990q/d35LqKv5KJUK+mgXfdFj6o0
FQo4XVQPFB8MPV6hpmLoqVzAXhabQ4wH/Pbq7SNmEHKi2IPSIm3J9U3YTZvIccixUC78F0pQjx3Y
zO5DREIgp3mef3vKKIEQVG0auBK7S/HgbtUqL23c71Pi/5M0xnHHHu4APlL84sLYQO0PfLZU8u14
U0I97mqFcgu2P21mLu/PMnm44rD9RqDUr7mRDhobna559QGJd0D+QLZHqUnTNm1V2nRD2EAvF9OA
glay9HT81a3E7MFWUHMwLQZFt7RPf+D1pK06lVpFMnXVWkUQQO/XyZHPqsQs5mVLM5vV++Ri9QAD
B3hte3+kr/uMgOn8jHcVyK7kr3vmPkL9Hq+6yT/fC92+5ppkycRDAmYWuwxZomNzGEb5shKsyQsK
1wUlIzsXwnb25h9a8lYAJFB5EEK/oJP1HJFa79RncscoEUY80hntyeQJzH4/Uf4UBXC442enkECq
J2bVYYGtBMhy7HHdJMw8DUs8j5sjJOjXITMZ82nVUqB/u+MZ9dt65elSfq3Crvi9eZT8eL1F2Jak
5MSsWb43ukCcB0n8VEB2vLSu8B3mdMAW+e+C8dtuSr+PWKTjIIwV1cMkmPAlgVAYTMRGhmcVRnTN
nu8bKW3RD+dFAg3olggcZdFeN5c3VCS3gcZ52aGCvlbGchWJQ8j6kZnsXgQTfEAg8dU9MW3UPD7C
i/JtaZI/WiZ/Nk7fTp76mrZLYw72N8voA8oLaquWt6ZCTfiYFYqoGdLtc5MpUGQTXQjLKQ5pqzra
3PG420xUQ1TD7c5NbspUWPj8QgiPdjcytaBwcXg3LP6ImhIIE5kRuU4GE6D+LBpwRP3WZZm+hQny
O0q0qKC4PlzGibZ44bcHkYGKebUq5E70j0iJUGxcFuQ4rli10JySgSKjHO4qKebMnQCz/CHxg2p1
NpJ1nIvFn6LJRW8E0gGAWmLxGwMIt7wVWtEvqVd+JxWD+TAc/s/jQ81fqeycQgA/CPOWLZTeknM2
T/KRR1tx3M+e5BP39GY+8/i2r3CHNBWLUffbdAcj/9jDlaI70N0Tt7o0qWsuAOfBNHeOmRqA+0td
EDyAaqR9u++7d8k7qC4BDGF4a5Ie7/TO/u4yI0LOeleoV+0OnZNLADphLg8UWhy+sVDx3s7DYqOZ
EoS+qSCake1WsaqJOHJRfXF4F9kR02+DIxIIpDAQVHYdRE+QhutGrGN6dOJ83p+kXva5VzV/nyO2
SRCMYNdtXmfjqsX5IVM3uFZEaO1gm0aAr0PEHtwzNV2gX1Vqe1PtcckaeQzn50a7SH4b31pQfbgS
eKbRYORLknLN0FBY+Zn9H2e508raho202srz8wf4SWM2nCODPME2U4JV1ZA7pnBUdpQ97+MRKeHP
Iym/N56z33p8z8cOuwHLXUBonknff5p/kilvP+l71GNUlsH3/yVsAQQ/+9LZUyF4ZcJ3y38l2f7f
sh79lk2GV7RL7a9OXgBXM1rBPpZmR2iQRS0jbLr9ttdcnWWbfbyqqT9ua063kvV71qAWcrpIESuc
DDzbFINwZxYeHqGGDkFthoAjQGrepqTpCXJSqxngRvWPxnk7v8t8u6dmb/FCs8HdU3fkb/zKXr+p
f5MKelZvSZ+R/OCxFutWsFWpEVCPHzRD7KSDDXy1szgMAXfBiWa4g+9pVGPh3XYYd1jBYN7MCSgZ
BdZpUQx7uNPxk6f9Bjg8lF4Ky3oZWGNWJx/XLD0nag7y9enR9Cg+cl6vdp8smGmLA/9fiat7epFu
gIDp1UCPfWx3l3MBZ7PQeMY2uCaUdMJQ2cW6Y8IMvAMvuuIzLtA1t6A7Zb1J/oweQOi4o85kx5+L
iL202JAgBo3Xz7OedtegPECehSAL0homJtlcYZihgGrUHcjf5O/ROZf73B8sBvs7lX+p2NUgcu01
/WKzfIKSetU/luGk/dcbWfSO5a0hW+lAwQ/ngVak0PeyvgxIGyD7STcDBTS73CSYkc6UY3OM+2FH
c0X3FU0bXl1644NMGKrJgnoCMN53ZuHmwWcUun8rJN2ULaKyFAEnhAoJ8pEk9spExbgWXC6xIVsV
z5uFdqOev1iJPeEDuFsOp3PfcSJ0IOPhVEVtB5LR23WPeaSQwkvtqwVYhttlJmkJK0NBe4ErZz9B
avl/6sfZINL95Brh2n7vGIldiwRPM+f2bFt89u7IKxDdlrDa1AaS0bYUJ63mNWoMMKAIv048zznV
hCptWYXufC34cWNFmbfB64SqVNlN8/E2h9hCPgMN5EsAMqnHZadqI5FRITikIB/80/qDmJzcB8uD
c7qb4MCAAUUYaCw6swsjFuVUDvwnWt1tvNMSR2GuNpyp3YzWuk4E4p21tKn1u1M33A2Oa7DIq4GY
XBM4iHR4tLfRTip8eLwX5we337ZEqYryaeNI/EEc6cM6PYidaLqd38ByWfzrMM7wUxZm3gazRyWm
ZrTRZt5GEz2tTI4ez75pOzphL62VDTcMKWqCcX+9ZO0yY6Le74qRt8nZCCE9ZIq31aU/e9JvPDUZ
yXtV3XeJvXXTMI39X7H/uUJFLLJtAKg6KVP5f7G4gGy/LXYI9uqeqT4fuO+Czue28nyTP1fmqRXW
bAw29JbCOoLhn7k46ZZNlgyuiCtku/o1Lsz63HnQYDqRePCyS1rZxpj5Doc2TCzf/E/QNr+8OZPd
0MjpOF/c69Twdp/aS7lQKgglVDfEffLYn/ASp7m8XZnwNJE7ZyCdoG9nvFGlT5B8b6XSFw9Z5Hvb
RNAbRQ+pu5lJStSANwEYEBNqkdqoFeAtSIJswMK/frOwvGIq1cB8XHnum3ofnt9Qen6Rz6e4Biu8
Xd77az6sQJQP0PLhWuwB4d6LVMOKaNsSvioQIpbqTsdos7oHi511Yaj7DFqKhgzpDYj/BWapg1bP
X1SbJIm4f5UyHn8KFQ600r/ziMAUg9uwsHQ6/H/4ohKeGQDcV8mmBFDtMAQKCWyDTIShYy7MzIKi
LeKvfrDXygHgBHYwizuYusJjVXz/myRue0QquQTy+pHaYjTYVTGByNAERbugE0BOIcGzvjQumfuZ
k1K8nP6my54OQinjV+K0OjeWIRq1igzsQAdUBMoy1SfrPsNquTTG16oJ3fOtHVeDUbxoHYYTDv1x
OmIhx/xm+6ylOP7E9EFktuaJrlWYbhhriBkyM9AamikhHAqQ2HLGDvUewzbiPeG2WlvWGHO1GHbK
dClQ6olGLZPk3GRjJ5/081ZtO/+3CPJW2z6I9IeJXOAz2CZS6zbrEkf/4ksGdTqFUdhAKl6Gw7dy
hcEZQhvkX23ilhmrygn/UcDFb3T8fR8oUClYYJZZTsp4VBve0gfZsjUwV9en58SoL6po6grugeGk
CIUu8KuiOfc1eCp/n6O3gIVuyKVaBE2ksygSmVIbH6PUQwTlCaWXoRXB2NLLU5yzaKXB2X9CViZ+
i/fvG2fJMXPIzY6tTLhuxr2jE3cMgyE+iMpSoK10U4+ZyRLcnWUBxYISuUR3RKKqfodNyyO1LdfW
CtXmWo0LNHHDpivkl96+8w3/htZIdP4B1FOOdNXfCMWJcNhE15AO2Xs+FH4RW7A4fXxUdgG81N6C
GTeJPGTHoxZTcgva09HX0SW+cOnIMRxOdBbBJ7IBBlfInOSb6K+KBgSnKy1aYgIAgoFirZUctWBc
M0a10M8+hfMyyuOycm17NuHmC11r1TXHA2Mygjev3zBYW+V/NPgefNN2kOqUHLJ1L1nbbR87AtT/
o/x7k80OxOG2rMJMXOXW9cte2dGxscg0FedzX5exo+ozA4urlhFtmlAVGGBP9+SS1kotmAYCNiRM
R4m8M7hiD6e52F2nO/QPeGx2JfiKXVozS/e0SUv6oslSTTMgsUw9gSQSFtm60DY9VfFohiOWBWKr
zK45+KhTS1dcOloqQVX3VG9qrE3IIpnDDn+wI+n821tIZxt36v7robzs0N9nEahPxG67UPGES6IQ
B8MLdmQATdegDFVVciwjn2gwfftsCJacr9UxSqeYeqvQaKbApihOtSUdcXW0BgLazZUzd/ly/+NQ
XJkw2nfiFytY07TqavDJ8Ygxr2eqGZuw4bsNYri8xkSnic/bMtk8MSKCmuI1EefaI1K/UNzgZYVW
C54drQJE63h+YC6sGwp3SfqOii/TL0O+q/+ecrSDw/k6uaigUet/iPyBh8HVml+vmhQt2NGebv/J
8YKC4Y3MOrGTHYXR7oqhEaTJJ/L/Z93YpnyZALeCGZMJdRFh+eWNh577E+PTbz/8o0zk/Kk7D8kO
mKQalumItNhCZdWt2CviJThgl+OrV4KZU/ekcW0ftFtbv3gH/llIXfKSyflGUdxB2mMgHhDUu2kQ
aKx41Biq5HfPkY4dCVHHY0SkD/lW1Z4AVVfjjMw6ZMg8zp0x1WISEEnjfEdPrs8oBeSJWlRXi784
uFaoxXXdv0SPpcFiqz6CW3kDe44eFaGWBelmeNtZ9Ap7ZystBBIK6xf51POKsoX83tFkr1GAM0Po
s1C3c4Cx3Ra0N/to5qd/JvjB0MzV3r/nAOFlC25zp3QgC5283yJzYH7l0wlfYaL0w/bjfqKcmDS/
qGcXb/3DbZEgaZbBqqDJ/XsE4lnTmWcRRReVaCuOWwXC9sxbHxw4CpGGClvquMjjzWpMrU8c3kBp
xVfbTHjFrNVao7H47FtzWK6OJv1oQOi42TBJjygyxtsi0vGVbD7unXl82Ndxumx9uelLJeyy3dTG
wTe+aBUYcScS60tUoXckX+M0ncEakqTqUTpyO7Ufkks+2E4gJTdUUDeatMr5gUoP+qky1iNfXB80
Wd16XFaKNlkz84tjdbirLC82YGhVnHb+lAqzUMOU9y4DH0Zpbvvou8va1BTm2xFUv89RFhHraDJr
BRI5rcSSpYhdXCAiROE3z81O4FqdZOW6JVWJrgULfIUFhKzXooey/TDZFbpWnd89NbYKhv3FdsLj
6VpAfstfgonIfaRUqmOE5fk8TP772AF357Q7EePiMY8G0vBQW40KgIhmIdukjOFTU0Vqtzx+q3MZ
+tHzS9xff8zefuLilUwgGDdL85gPAojv9ZUYOJUKnUkSvOPpy/bibMEqrg614crsyBttDTKd+6Ov
CwHjJhL+bXlD4tCAyEd0UjNen069MInThfWOAhsLuRAWlz19/U2b+uM3FO6xohoWGBnOCmxZeC7U
CCagRj0IkthPWObMUMAWQvDgWiL0aocukv+ByoBuSXqckzV4Leed8plXr4ezZeMXUN+LPY1yYCmJ
IQxzMpWMTLKn+3Gxuhz9VcyvLBnD/1E/W7qGll4lIjatCVNLH+gY200nABrh60jA1CYe7XD/FIq5
n4zK0+tyH/MGGRfjOPSp7F3UHCouK2l01yag8niRm3MbYa5usw9bNUDEPYBwnZIm1vhb1XlapW0s
LyUTTMEmHQlle2pfIqYwD9jHTIFWV8NxVHygKQt5IW1UoYcq7NQr34r+RcqbbVxp33/F0BafVps4
U2QJHi6cKoFiw4l1hoOeTWMlQ8CxcGuuOh37KllgBrAcLCGr7gPvrspMvxPTdXxifSBh7K/TnpsW
r0+9RLGU8Zk2EzzsAmA2AJj7WbE+VDkO4OrMBNcjJ9e1IyzI7tbKDciz+tPVaCM/9s0JXWcOp0Am
Oc0PZ4dkKQWKh1M4QeNPxAmHidoZsY6gqhXSUac9cOJfYBRu+EB6SKCVwGZCrRD1GW6a0zFeijH5
4jnOwywUDKldBF608lzyKz8RyjRNzggLgTTbt0olgQkKJ0m6F9PWhnr9zoPzOSq76E7m1gcxQSdF
18kZpHaMl13FtfS+GdUqzeFobwghMc4p3PCd463hMwvCVGS9lVFu81iVP3qCjmBTYKMNuEFydBb+
IIMBn2Bpi2yZJ/6HVHlRXHc+fe5z43wr+2kvn3J9X3TGbTk2cbW9NilIvzjnNOk5gq2+IOseKoBw
uRrckM09Jp5GSCUDyTrJ5EpzZyvUWiMyHBVkhOks3YSJRIX93+dPY2426vQpraZIAQtEII8H6KZ5
zRkc/0Ctie3h0S1jKktKhlMSVLNJGsAyOBYBK/W3venCrlhmlYX+c3mY1dQ65rdcR5vE9L9M8n56
PDjvYMGBwe5Zcn11W7M0cn9AL+9hQuxE42JMZbVInuR44zk/bHHsm0/IeGyWyd23GlA7d5MAIrgi
i/7KTMa/NUoEqCgBCEDp1fCsWcMhMmWQ1r5HJ1GPsOrhDcQs7F6LEBzAGgzB7FlOgMR8qP//UEWK
mT4AWl79nZDqPABlBdQoMTFZn7LVhW7iPxHJEDZQmRTdWpMkhCXVx6QG0GoDK7MUM2iv/TyhILQa
gog3tTj3/DfQ6EyRe4gjPN6cFY5c2dmMiLjoSBarA0FPJ63Ae+LskEnb8b6KTHbqDZZd3usRI+Ic
w+LLXpEispd+E8cEzbcsl01lqzcEcvQj0AbsUEMmiQgnjqWx2fEFq4EZ6vT+Z6GxhHcW6RN9Py1Z
QrBAyRccVnGYBd7wmT/mcilXetEciHOz8Gz8HwI9L1xE6iTnvGtWL95Lj3g71v/rS9bKJVi6L2nA
XwM0XiaGU46AY0i0DvOQ+iE8ceHcjfmzocMvZ+iwX5oWvs2juMnlK9cRK6VXnmtUAFhn5UyidHAz
79Oy48IgYhbwTLtHzE1HOyPzFdnB31b8e0HTwx22ZLBZ4tOb2GDLXP3HGtytTDRyT/byT0/i6ngx
9guWOQSmi6TNWZev1u756nUBUdYDezKUDFrgjw9Dw6I7oeZlSMNGp9shADyeZzvfm4YCeFKZqQH2
Hqsuj7sjMTSvbSJVo7I8IunnsjivJ2teZRrbQdxTyjwu9Ho1Pp4Fm8CZvDL6eVf8f0+ijrp80fmB
3suq1CGfDEBj82u5bASbzy052MF2EMqFXLbS32Rfe87IiiOy2Mu8zJaIyl3Krabmnslwj9fPsj6T
KE4DzoUn5m/jyOZJgSO1oM35s+QsZplrHE1KoHyxfQhF+IHXdeO32V270GoR+j9sIex8JqlbIGQA
w5KYAJLkD/Kp3pYseRLwBGUYsEsASLCgZAPn40UkcR3oyoiC1XUxVM/UNz3gb3HY9cShJFIuz5N+
nLyQuvCa1shscp+9gMuQGvkN/aEG16nc7QbdK1LjDfwyDxINKxW57eMcpKFy+7I+TE0qDiLihpso
hX2cKDhg+GP4wpt6saiEHP21GjO9kcXw31N/R3G9KyGShet5UbWY/UyAZ6YXpmJSQpGLoKNaRJnK
OvKB1Q63decIn3OwaTF76zCsqcof6PdPE7UCjy8NXfjhVlrIandKQbWZVwaovPBoKFQfajzkIcnP
LVlnOYG5ykmz8h15r/kCe+cc1zOv4wJ8SmeFrrVP7CKqwzMy3v/NgrJTwqmINt+NzDN7bCcqwiZz
x0VJcDSfbe1/RETalk4JRb8Set2QDQqzrOu0aDxJLtxM31zsaO/LagAQYQTQtdELlqp6lUVJPivZ
uvqiqC7gTRSuGbdSvzDRYZXwwp88eU5Tn2jQA5X1XWzZECzZmm1I2w2tMTiYXvKfs6MiD3mDqX/z
LouEOf4YbWBw/bf3B0cCf/WZo3Ikbdja098WnIkOxKV2h9JtxlF1Q8tKRG18E5/L+zw1ZKTLbpHR
5juBHS0NDj+vq9XST3XQMOCJOLFVGPWtnA0oXHCEtZCk/ElXfnGg7tx1NNrsx26g2Vv83QFYe6lc
0VMTVqeelNSGclMCJLfIPpMgAr5yPigpfj40McnOy9rI/6wmRWseoOatnGqaiUx1RHh48QdLUdAI
BCsOQ438thMJrRwmtZZBN6epATeihr52KQOEI4WMT19E8otMzh/5kDcsbQw6T4AsMBEll+beMdqX
lMS/S7hx5HugwzIoop0UQtMy275qIWzRs9+g7HMaWnCQIWVVkAmp9GR8PxLshEEI8TOecXKkvkG0
/0r8Yw7Kxb8g+uGqJiBw9nhbI5dmm1D/YfVpHzzTLRov6eYcShe8CeVcbvCrQBLIX9GgJRw0fO8x
eTuxY41HlEdFif+l7DBtmpY+MtlBYkj4XoUcMmYA4dOJqbIpFqAxC+oeIPGo/kvjOtMkIhr+xtV2
nlpTDqQLq2QItzok5Mql1xMlntwvSKBdkpiSSjBHVHjnIlNwO45D5TbKl5RCiMTy7V5U6kGqDgKN
zq8VG1zfCmEhFKttSgpcrjGvCfKVBmlbAZdkTxxCBQd5Kb6Z9bYAt13A4lsg9C57jGM5ZAyjnax2
AH9RbjyVWShMLJxVmUDVvU6KnNy2VL8mzJoDwWDTnIsGQDgRRUYfAfeo2vjQTsDB1az4CBIZC+E9
S757nKgb7cFH0g//FkPD8lfTX/lCGLtaSeGnrkPHBqBwKpT76gJwtFEOHBsU7+P63CUWIVhYRzAi
vLY4z7v4WZSk2mHwuX/AM3y66xYsAv1P+VMhy83szTxv3HkyqEfgwwZTGgCNEE0A4HLPYH2qza5o
IMWtFfq78XcpSjHHmKfhJNUm+d8cKBs2A9WnnCdG1nX0nEkavRwCxpjDalJLWvg0+2tGUFtW0990
eVVg7U7BsPQMbZSR487qrF2vNh6dn0lOGg6P9JFU3XYiJJevJIHX2mhkyMFs7XfgYHTHvVCMoEqe
jGo8CXz/BmJhpubCLyTEljNyRuR7htOmjfBqPbJBl0S0wwmlCZmOji/MNEtkKBbBPULbgPkPsOcB
60JfZ2RHHyU8sRgn5xFw4UPsVhaRdMCLIHtEfBwH0O8WcsM/KOGK5J4EC3vF6hKocFISo7Us3lvQ
MHY02wjXuFdSntFXCuawaARMf0i2KLEl4inKwiFnyMFqFmp1ISW6urpp3+SLnQw64gCfd1+4s72Q
Fbhf8xjs32JTtC4XZlOINbwHc3Z08OzVKF8t/pkzI+tWwc539d5Xm/EVolfu41TTPvZkbULxAu1n
JEV6lVimEnHOQwLuDCKAB1dy/TPeayl78QW/Ig7pfi1evGRX8yIJifFZi+nIzKLhi+WCJPO2a2h+
8SrTajm4jjTi700IGv0nQqhOPVrXokV7eg304iOA2c9OVg5Y7lCOfRnLQ8NbMNBJzBn+1CV/MgTA
fNUJlP01Ygicnak3yVamSzKc546vSbjCyjj9iOLOSPx41ULL23EVuyY7w1XXji0+dLG+p3BafrnZ
z2trmppH1jyWb7uvo5bzJUTwGTuE14wR20g9EQgBcPja74dFaCQAdY1bnEzCq8SZ0NWHr2qfjsDU
DSFeBuGxLzuwBjscjQeMdBQcchKEbMtbs5XPPeM9JRKhvSdmDQ7GtfO8qMIr2DG5PqqNVKcDtxFJ
5KEJ6w93kOnmEGwmlVCpx3pKzYyDecL1rCp6gCViq8mfcuDBPYljGaUUiZeqsTte8FF1qeYyixdV
cTRZ1rnGpwChn93yiXFgLzOUGZ4NCmBX9d4dNL245UFpYNAwl/+jFSUsvKvQlkFtAV7g07dbqyeR
JqSO+lLBwr1tSt8ZKYgNUcxt8aDex915PU0jsm0NUU4xBe3iLhcA5SLSDgXi093dt4YfxAzGeNzI
ZOhJcwFoTukEQYzla2yEk4Gl5ZS4fHJEWSrY109vBaVGF1F8P8JNAEdMocCvAwofB2BgybUaIpNZ
BzajxIXZ5cIAf7WMVXO/9K5ZA4OqHyEonQMAQVDqL/Xzi8dzGg9BpkVqpyxSONwvjy5R6xPxOGx1
dEEYQUnVpD4VHG61nx51kKSOsrNAzOY7MDM8S7yJKUjA2O9spxHjCfB4EQUeZ3cNYMbh2UUplTie
RdyzXJZK64gS1rHGPIyav2jHlLYqcRtAohTdK9+cEfawVU+ELb+PD5tjpcOvUi/pnrshHAFScE0C
HGgurFfH1wdhM0WU60dzzXXIOb57AusTM86t7Zn68O/1cUcCRC/k6gJYwSnXi2dbG2hbkuOg+wbY
2KST9Ty9/reIM+4Weq5MMLlYSSJQQD6POANo45fdANiaLiX9qKx7pollur3hgReJF9oZowIz/4+i
XVrMxc3TVpcZ4k0XZSQpkAc4kcTo/3TwIv0qmbuJV1dJUiTxSB8A7O+Udpo1EwVBexNN4i8fGpcu
zo1gAGVZ4jOLC1H8QOTi+hf7QFjJ5qpJuzirBpH3THc477tnPe36x/0OwPPIWYU2QgB+2FRmdBM7
iAgEVq6ctmWHlu1Tw+7ch/EyFEPXgtGSuuLiH+4luepNT4ulmlkr6KRM0zTjXMH/sZzQG/oSAnGr
47f9x+bVLEsvg19tzVBMDZXsxSjhNbM/vgZ3gfp1SV9OJz5BKKKwXIjED/2XF7zDK3jugwqB9++G
Kz/L/BJ+OVKBOOeg6aADrbRDHXsau5RUQE9AWo6uX3J23KJM4B6ma3Bx2pU+dSYBtcEO1zxsY58x
NtTp7WNj+X+tnVciXexHa4jyk5hSFmMLQ6WtcczGhbwhGzyQlT9uH/XhfLl6gCnlZfq1Zbpc2HO6
o0i5jus/pLvMX89qfQw87+yvU2F5ifu+g+EkcISNpEmqXaUpXS05dah9RtRJCeRw/BuWqHC6q+4a
/uXuHczqI9tAXbKPc1NrOrtirFII2/zjGd8o8Y3px36ubGF637kuUAPm+N5mdS7IlsTTje3v6+qv
k2H0rxbyFu5+bCbQRsffiTwagBFRPanCBuSyfn2LqrZKT0NNJUd7Apadk0USw9xQfRUVvSQMmOQx
PncKlnIdUUdG/KpHSPW8sOYwunCutGoeXzQls36ISvsLmotPeETXkMbola9DuJO/SBWaB+5vEJBm
LAanRu6oLLSIjRlR24498jW1kXco945NRvB7DVWY23iXYLU8YWc/bseve2rP69dZcm5KtDzpJlVV
5ZZVfStCL4L8cRJxQh0FDffHCtcqJnATBNjK9sEsUEmbSP69ZcjM9/iVI11zbiDaVJ6pA7M0OYo3
DGLBpEgbcDJEa0IElUIcBredU1mZnBysBKYKVjZYbsLUb3Xs5icu1DGGwL4kU9iltIzNm6Q5FoMB
iBSvGTo+mklQkmmYbhoTrmnj+IVIg70zlztm3iebktGESUQI6hHbRr1EcIVatHbsfKM9ig5InQnC
vfR6kG3bHtKFoyH5A0FipDBGsEzQagO7BCXeVcDuOVEfo0YjPZ8FyOdqqX67u/6rYUfVA824Cup2
OyU1vcbi5jgGQzTe/aXbMo3K9ABwAvZn6CguRhmxFJcynMJF6GzKQB29dO1i4XC032enB8T/9vRS
W0JvscC0r0JfETVWOl2QebNmW5XpGqNClrgxJ3X1PsdicZwOX1J4zb7Uxy2g4tjtrcCVhdm9O8/7
V9z0VWdaUxOJE7H29fgghnpSOOHSDt9ggqkMfKdX5+fTcLdrbohakXcD41QHHL22oHUBsemnxmRB
WxyFM3GV+2PpMLyeeqpKVepN3j8+Mwhyc85176Yvpv262NAlpvm2D/NjIoLYVpOvQ4v/JGRbiTqe
yAzTmyxzpunWssk/l1+FqTRiDWO2cZrLzWEpKh/GzXmuUqnWDj8RP/gXkbYD3XP5sxBGUHO2eDoT
vXOgWW/YTk2R5UMoE1wUFr0WLxp0SpYzg6PZiTTNkQVCD45LsE1X8pHjDduqnJfkh5V9b4P6jekz
7x0zdaEfLp30Dl8v3fVSkhYD4b0ZDC1u2EL1JnxaewQbQQh1AIUwDrwzAQB8BOSkSFeYbqWPWmC+
6+DoPfBe2m5YW3FqqcUa5lt2sS4vCQBJJhQ+JtqkvIb548HKOlGI7xmhsFN0JLILYy7CcrFAM/2t
0Cskhdt4++uvaexPQ1Vaqx3f21OnHaznvpsbdZXiOR7DqJJGU8E8b/Ch7uPpXwyyTot6o3/JsWyW
QkHJMcLh/uA//H/bE6uw03jjYn2ym/5mlZD++hQA14mspCsFB/UVf12hRqTPJTmN/Tq9ahEv22td
rJaTB48RmqRveBxmYIJfvMFZzURY2r9IHuqx5JeUVBjJVBynvYOvlJFNKKC9ZjL2HGKw1gOYn9u9
kfyjPWQS6fEkPPObHzTJeQ2qSSXcMGKmZj6ntkh+J0K8EKCfPqmDaU0fGuJbEspPRpD4Xao2KoCY
ARgvABuc9E5+arvPU+3BHRqWfTCLEvtRjEziVV6peouSpF1ulQXVBjbnmPHt7+KTOMqB4B+37Xgr
Ld7xcbY/w/WcFcpkfFiy2kgbVAYimRGqWtD9+xuMfW/2CZyDYdx+7J4QyHFGuP05zQNxiyev+H3h
dYc7P1ADgVtSMQBL55oNjzJL/5BE4JnIsHtQy6H3aQ//gAVR3g6kh32qitl+bDoj+QxSIwZgMKAu
w2+0cfifV5jxgt0fTQr84ox3R0/0ArPAp4CYfnKY2bM+WveipG8wgGV3H8SmV/z8yQqnt65u8qFC
omFAjq1Bww77z9VX/XlThD15GAwuBCqu3/28dvE0KRBupy7besed8wliH13lC7qdNmNS17FeYtEc
SYHuF2fOf/HK+G1yQHSRM9s91MokjLGufsFS/tsOaXC16w89c2/c/7ItnKPdyNmdoAmxzwNYBoPI
pEQJYcqgwaETvvnCeKpCZITSkb3GqfNaBi3TSgjopJk8Y4Gyw9maf0sIcr+TkU03QaSWXU+8SG6v
fWfQ3DrWDanz8uZizIVfcvWZtCeHtlxPeeuoyMyVdvzCMEhowkvONHIcgEzjEdAGFnAloFRgTFK7
91gsCyHlTa4dPftbWVzsKDSKLabQPwGV6mS7TldBSk3loLa/CYBM/syX6qp0yecGbq9lfFTeJ2IB
ZeuZyCVZ0u8F9cCHvOfFQEFRdcYSJE3QQgA6wWX7L5bZjiKjvOpRAC6iLmph2FVwzjybnw++WmBu
CDWOx4itvbmiOICWNxsqNChXmJv45Ixw8e9mpaegML1vK5ImtKUmxAAe7IemHx2HWmLtJv3zi9+q
2EbgF6/ypuFdtpD8xDD2HvCocMPRdqzg/1AUIgfVgjxPLu0CP6IKQwnCfVkpyQKQ5LCV/IhLMNbY
rHqvREBn+RAHQw9zD9VjkudFn443asx+uqR3RZOKyFtZ4DpIc4bAERbSLLIS0fwNj3BgmAUeUI1q
PmdBdg9a9G0AAhnEqTWD7/OlrvEk+OlZQLwTUuNvJmJolTi0TBQrVKagsNtJIvJgbxK5NB/6NjxV
jrSypJtjn4u0Qch8ov8MWoVWkMxgVVpR3nlI9Hs/PoPAtmVuUH9iDiTBWWT1dzVqSdINHl7sBlMb
fb28wBeswtLLFEfGM1j+EABFrdp5CbdV8oAo0nFew1Jg7SuAqPZdXdPvS8NBgQeJhzaT4wAXk0Uy
ohK6APDO4noQmjc/7oHbagJMeMrvn7h0hgiSrlfQn6W5QvPbhjFQVBcR7oXCTQETkStGmqnrNBNK
2BuZFpKTqR5jU47lYMJfOnMODmEyzvjcO3SWkaO0Hod8uzFjl//tNBVAl+p1jdKZFpYKIlLajKJI
fEg+3+yp5rbRiaMaZxtjgVJkdirvLxtybhxUv0dfK4AGfMWnyjv8u+YfY5rYP0brvEKiHC+Z0kNJ
u9XmCKL4kb/Aj6fdh2abVQTgGyVvvOpt/MOaHMQRL9Ws54+oDvgwMVEG44wC5eZwl68qcwm+wSMh
KauXLD0Uz9/yUa8JntWPTS3FWCb+d/tiO9rLMrRyhsWX6qng2IX2L6+WRGUPWvW9+YlpfgicA+h6
+TfS3/n5OcJ/H1VAgyclwoT4Gx6UnBbmaxav1bkHAy1Acyc6pN8Et7qnjzZ+mSryU+HnwBzJHr0G
Hjd5imsd0Olc71oyzIpda3Wy43MxHbse+g62yISI19O+YV17TR1PT6uipmWkNx+0fpCJJBGpV8DP
fTkJ0H3HUdEv1TQc2MOmAjrXAznTuMvV/Ofs1N5iDHk5yG4EZJXmg8uvj6/HHk6KjGAHvGEOuLkl
2qNQs3CK2/7fEHYmc0wQs8ysLSAASKmBWP9RLy4fhjAL4SPWxcgvmanjd0thGPcwtmR3xkB2L4ny
RZ4onxrSrsShJF3AYw0ahoIJDlz0ISplCgtD+1T9u7j6vd8y12ClCbaIfhJrdYPTVsVZKYHvBLTC
OsAbQty5jiw0nZZ86+95NcB8DjKzT3QzBv3FxnZCn1kInpFqyBrMAzSeVWkGEoM+p1pZsBq7BR5m
4IXV2+ug3UJs8xXXs6JaSQZlW3XBDz8bp7OJ8QiE3zbvVZUL14MryrXH1ElxmVJ9PVFtr6Y2ljss
KeXi8z0rFg9xQE9H4+MxJ4rxpAfX7VGhp9h14ceqI1bhaLdrNURI3nw0RTnm2eQKzKm6S6r5HIsR
0k+IpxQr9uAt+YP9LRlgjQFMmwnmqyt1kl8roBILYt+E8X3WEDhAj0JIihrsr9TnNwNRo40r8AX0
NfkcyT1pWoECY1MonOS4iCT7ocFEE+e5U4n13Qy0ZxiQB8LBTo7aPkdOnDkW6x8DGavTBI3f/7t0
kunlWAeTdNVucLzwHyQWqzTUnwqLdmGST+S/NTeAnfBYxq3xHeW17IzGHDdFhZcVw0QfTnvGHktN
hfAhU1fPWGxrb0YMYPajAW8i0noJKwf99jWuU+4MZDEAcjXmfnyYIbdDCoJ8NU26pacmpgpElCLL
XkxDzLyA8Ucs8fJymQNyLqbDnPI2CKz80dkGHBT8BwXeF9d8upn4ucFR8AigV8gc50wGjPG3hJtS
pAZpbsMKq1NSHFyeIoSm1dZnt8FDKJkT/6PXk0nkCccKXmhXj+YMiAvuOCbDvO859LK1VAwcGF/W
itcvkqgLYO/VMswhCPMU7/k/Qn3eKMY45xpmKOSWhrLVA9iGE2vnnnYOdObVu8i8aJkZ8o4dapa1
++ZC6VMsyuariKOR91pvSMObop3eWdoIqGuwmZ5QvVYW1SmWyFhmljXhUao22Zmgyh+1tfDH1QID
tHLPYgPmRlip6YXxWylSa+Jj+vkJXAFog+jysh6gs7U8dnzi78HUn3ZIOSXcUyCuB3yd65RXWORu
Xn4iTEB7JM1utND3ZIcUW/SvsbrGhH9f20WTIIbygRlLd1bozXBU3YFq01Lo7OqSv04D9FKTowzL
v57YqlpdKNls+osr7XEbsHFe/yybZ6gB1qTYjy/1lPpGAzD2xvmRJFwE8nH6FD1N7Zld80QMLKZc
5SGNJmhh250GjLZaXDBoXpr6FkzO58L7/CaNanygRSfGdW8Nu2XQ+ih5xGHjLOEVvc/+Ii2iBKbJ
MMwpWdCMKJB2xj0MQY9eAk5cg517TJIhNgYgDD+sMcGcJtpyeACc+huXRFS6401vVgmx2dtaaWVY
yirioBWh+btwbbZc5lyGZm6+L1p0IanMk3dq6iBn4znkplNpGUgSN5BnhSnQuYb8re6zfA83C5VR
5X9C8RHm+p+PatYstwwEPZi7zp09cyMBaF8ljWoO/VWooKBXR2ibmHce8PdM412KoB79/dTiX95X
64UW+SnWEJAiV1d9mG6CohY30Xziwyb6sJ9IH6CfehVOQshB48/P+b8ZY2S8c5rV6UkUwH73PWCs
tPy1cJLNsn3Vbsc+u/p32b9l84pQgsj/88l8bRvr3GmQLPyp1OckLWBR0W+rEfEntz47BZsIgS6L
1fzsbR3vJVxekw/A8ppoO1lwGdrkDO9JCiy5vEubJXKJZ5a7fwp5u2AhEBXp56inXLHt2KmLYm/E
SLETA8/4ZIAw4mFm9fzTVgLNF0KFrLFjOXoHrbYlHIzd9TmxrIWqMEKGBoxWQZ5+e1PA7B+xjg7F
HQr9J6YBQcNlgwwowwCyuaga83F/Nppa2gQjNzWKf9bmMwo2l5+KGhsYa4xCaPfoBfABQD64Bein
bUQa8645STDmKsL2lpeAbW/Mg4J7etuClxvgYYOdzV7kcDjcB6V3/1dg0fd/Jq+OtOz47KMeKQgL
HT0img1qMuU+V0sCfskshBBSp99ZSeYCvdGFrnHwJ5pGhkKSDk4yYIfbpyOvfBeLofxzF5rHYVdE
VHcivSolg+GRDh5GmuRMv5bcTKe34gB7FA/SjtFaxiCgAHS1P5L2LP7LL8AVypUVZ+x8rAyX1BGv
9JXpb218Dr/ZUK3zZCqp4RHjzcw/UI/Yf+37ggU2pOrUiKk4GBZwjvOj8EGBjg8FM8zC0DuOVPsy
KiCZuBxsHaHZZnfB8lyBP/sfIvxampeSGUQtXQ8wON3TbdiD9E10zLrKxzXTmLWarSK4xiuf4gx5
NXeTsWOwOsGKJUIShllunZ7fOj0CnPj4RvgRLWWqwS1W0r/bqY8GInR++0eHFfZr0yOk6OLZtwEt
AtJSGeUrZAvN8EKn7DmL+xnCkD/MZfizAtK4aF7oDxWYgkk2PG97Nf2/CupupFFdccRZLhQUdrrv
K5ZOZCF8CLKKsgtp7QmXe19wKP1OBqd+57qsEdquiOJRt53jeW74BFStQ6mA0IuJ2O7VODovKGHp
E9wGPwLYBfsFZnC9Ah/h0J+K4VPw5xBv1JaEZmwbdVTiD45qc9a7wQHJ051Xe5IIKaO+7sp65ANg
doU6cIpvM+ty/xL6grEVcfckTKATmZ/6DiCZ9LUj71t009OXzDOEBiQW/S+dsC4nI1C1VSh88Rmt
aBWDP+iOsUJO+v8WDVag9xsXbivWViWJGH8sdIn5Q3/G+xSL4IOr/WjmE7EVrn5eqoK7wsluN4qT
XFDYRBQT2ap5frO+jyFDwZeg97wgBW5cOexJwgzgSkWff0pqk2nbSxZyUX1cpgleejMoDfHuSsec
AAdIO4/T8gAK8FCC/rnkhHkdr2UG3LIfIBqXMcgr8Pv0r9S6KTu6tUzwqMedoelkQwSXDYHBU5E2
tMkvWNmgVkMRjqibOYC45sGkRuTR0E226r+mLE6FRcRKtGsNLWIdZFrYWrXEkfxBSDRM283ki5/y
rSBdpWdRNkoSZ+QMDn4JpPr/MTm/jbm2hBVuXz0kQvYWlCazvwpCM0M4pPVMDhh50M6a3UyiHXmC
ZEVpeI82ccytKpHZgazGG1UBYhpNA7u6Tw1PzRIjLs63ebb1VlN/Lp2vbMfFEgPZio5kQmdyiC6Z
4kdnWjHgdHUcMqxJ2P4VSAzPiCVoFyfb3ZVXQxIb4aLqYxA1MAeIjVHmYrgC1yr5Dm6rT7M3kEt5
vo62KVFrUpICrKTv3GYZnV44eM3VXGzA8nHxFtbyYe1zJ9+Cc9LIg9TDFoJVkgsdGygt0+XdUChw
Z1omc1AylDqrzsAmNGMnX6T06fvWkQCAnYBrIILDy/dvOrX48GnoRit5aC6dGYHJ/AFPX5V9V4Y2
ndxm3NVbw0Sf3UqHVPsCqjP1zPnEoVHGINRDkqmZOGY2xGduc1BZKwAv4nwk8MresjoGaw8rqrPy
xH5GOFkBIkHDD9hKTQR0q+hGEx0FUBDhac5UuBsxlw0146ZjRYRHmAyaz/Xr9cnHbb8K9wKspdUw
So1IZF0RCwJKpqsB4Yu7z96YdrvGiRwvWPeXCEwiOxQabAlUTDpR21+KPlB9NELGZ0cwKCWn4Bje
YAPTsnamX8uVA8vNUj5/eOAgLAbarE47aPFQtrunpKhLf5rhgAeu0Mi350SF4gLXnFkE6UEfkoRd
wXlP2NlOL+It3i7QL14X6Q3nObXpTE4fT1CWwNKV3RGfqn8cu/MsTxLl/fxqA7wLBnmoofrC5AiS
knIhqLTHZxV1x+g2ohUVg7WidPGyCVC9H28i4NcYc+t4c3qGAm3wlP320+xRtHsm7NMyso4yrYUU
ZQjJaWTqfCPTsVDzkzLDq46Jilh55FUYXmHsLqK5woekm2x2OFBeQJU18Yx1WNenEub6sLCHdVkl
7hrStzRJGaYSvDn8p5YTvLxI0NeegejrZMszIBp4C64ph8dgnWaX7VE4wL39vaWh/q3WLOFCxJAc
45/azvUk4rJEhS4MSUz96OCY8CRGgkocd8KKBadmNTFifxgIBCYPRsRP5FeiU+m3dVG5xyuF0nXE
TK7nlvklByaMxRxD2bF8FiJ9b57tq5/vGtZeUlLhZ8/0Ugk+V2c0mo1Io1dAVGj5Y15K/AQkTSSI
n8tTJ0Q/Zly1SekdDyZ0MOc9mYUZUGk8GFsi/pGBWhMT+oqcBXN0sHhiIsI4R8IzAY2r96I+sML5
ebZTVoUdSoYaYKpaAHoxOU/CWW9OK811hkppnTUoWiZGvIAEFsiOKIcixp9B1XniQ+6azhq23O3K
qOS7MBacyTmNgMlCCu3xf5jP5KF6h+o7t+VIKGtYq1azSxu2lKZRZ1gBFwIVy1seuwqOOlA8b8dt
UMd6jzXAwjibaT1gNEC/t3rOWI77Hr3mXHxo9Btnf4ACHBqVkwTs5tmA/NxNKJzuzb1/EXvPWN66
RnerT/qo+tivBx+qbxEuNdlyrvUFfcXcXXf9ZQ4cR7+9j/n3l2jSB0DkDlKNQ63cbD8v2kNyqgem
+iwPaeKQflPzxyf9JctxjceGQy8mfxz6zwSJnL/hScovW6hht+Hwc39OJ2gwmVvcidjYz1gGOUTs
laH6d4CTYisNP/1uHxqO/hhNHliNlV0JJhpx5Kldgje+hNluz5kF3h0+AzPk74M76pAvjtCJLeAj
AbLeVTkkM5TBYFBbRL/J7KhV1Pqok0tbOwzdnipC7QBLIpBRhMYyXFtullAhuqe71X+5+w6X0Q5Y
MvBeQgQW547NL6U67dccmVopcGCN3Fx7rRGVVvWZpnJfzFS+1PpBFwKWVvjlXxpmFsa6vQt2nWWp
MPoirG5DeicsjUIEzzOG59LbfuDPBjyXZuwf14f8tYfm148dZabkYk+HBbsxAdTabCHIVjGfdKjO
xhYzQwjX26/T3Sote8tl3LOjgOjHuR2ImywLmaO69PzbcHCpmK2/luE3iUVb5AyvjxpaYJpvhr9E
AsgVXEsv6z6J3qq9riL2+ClW24pzMgpzpwOvwweqVIjeRbWVycGcj+/OrjwQO8LvYGl+SjXvGdBp
ZZBy6p+DuE3A3GLhycMqyY9ZfD1G9whcvTC8fydPLoUk8UlKIaTmw3XvryJHLgsEcWGA8GWyjNcC
ZNc1BWkfaHg/DvdBM96ZaDETgjIovUIaEdybMIvACXlq9/27EPn2uXmlU5ehv//SBiyfLgKFT7dW
dUMhUdyJRW7sDbeESblWVjbdc1tPgoI9zMERP+G0KKfejPgkzPKIchSkq9Xwr5IstJJwWhePVC3g
5hWp0j5QsZfqh7VC402MojpWOJqIO9dfUz1agviDRW1Uj6Mrrxa+CEgjcP+ma4PjiSU5itD7ek8G
/Z+8LzgAP7pQOOwZDYghgWylY1xOpgHfx23EhVUce0a5qUm1ts6DAF/SWP+OCw483kNp1CkBlos5
hffHZ0ij7U02B+ti5P4So78SUZAzq6dwzNYz8rpdkotMRynt9sbdMHo0+iTUUDZHS9sn1Av2GUia
AoyiftjWHjtBB/+zquelyuCBkLIZAGBLlnvIFlZ9dCYnnN/PnDXK+nfVD7tgnXD87jckf1SVXYzS
xGWc5IuFlPquOrK4K7SUDI9Ms8nm9eS9PbCT4bHETTWekaHO3tpoRXx5n1R/mnnWKVqhhsbw6Pe2
lQNGAoh0xKTOiTcmUG9J0oF2a0hrKfxZ2QbVzoPCLAI7NpsUmOhD0yEQkLNPq/fwdoUbRuMG/+86
bKvZXana2SFU3IfdHrC8i5wqRqjua8xbGk8qTYoUIX9jegLqwV3NKllJymUyMTAPdzeAsxUsrsEM
khblGZIw0dOIfO0T0sBM++iVHCt4JBRMJPgEZ9zvMMhUeo2mrQ7nDpKAQgo7f6UEDNqAjh4mm5uI
lzAa3pu2Z2PmNL7ARhozSkppwyYapC9BlbC+EHfa8gp0yF14491leZgWvoGNZSV9jIegz5KxIVs8
kQRmoVuqKALzeFQTP4Xk8a1rW0+s3wFsgMYVR1BZD2K4JKGP9eJOw08K4dE+7YQRnGpGcyGs8fgj
qb9ZPLCF6gsNLU2B8lWgqf3/xVhiISWy9asv4DTbXMwLpToQhMI5IkGPSpRt9iSPFAkKXY1s7AhH
w49wrnkjFoswb9B0vqKv/aWVmo0hXn0ktSxUS8D+w9QDfJfUcc1B9DYzHbP7mm4WyABE4eswVx4B
6tNzbcBODjpvwBGEqPERCHuZC6hoYv3d6PX6phuF2E2TYgTqfW2vISV46O1Rt3ZRhH9gblU5KfCw
IMcQAxWiYU5B6xpNs7X4BMGuUVEtUVvCW85uqaB2f02IcwQE28mj+JzDMgnV0FcPVUj12eAd4LYe
wRsJBcXr+hfaa+uASBgKE+vveWWec+UwM1iRTJSSuJ1eTdELvsJpbZAJ5qgd2RmI9Amv/CxDRKy3
Ylupoqai12IwYQ6TOkofrcOv+k1/yA+NbPqNgDvyDu9mWtF77V65LSEYzgYaeCOaybLg6rwKvfgj
Gk+6VUwmG0f5btuEKA2C5xL4drxaeXIKZbJmKCR/IZ/99MTtvKSjgDWgn/bGfumPZILIoTgVVgye
yX0dgdMVxNeeOZKFu3TEaCXMd2XlNEINhliy17t6rlHLaQHwu+dI7zMFZwlkJQYyqB0hxXiL6r/e
LjHsQz2Inr+5c/RJGYIDOD8+GLbxx6vi6xzuUYXoUi1572MUyEyhjpjtb6ipNQbNw6Uye/6ToAug
Qr1crrVHxqB4FvqNA0agBv88q9JNj2MrO/f0J7h2ZpNBazUgjA5Gotb2zlP2/MH4N8AU6ag6pcPw
lClzMC4fMLLE1/RaqEbbMg6kHSCP6cZUkIrRgDObwU1zgSrutXzbUtwJZkIuXB9A3ddxtzjQWfQx
OtIZcrgR+bVKezds5iW//jXdV59SSrUAdq0pdadXSfd05x1y6aqYS2gZIQjIp0Mh8mNC02GYMwFd
8xWUEXZFhTZYN28B91cGoxawt9E35yHNW3sribsnQWxseo3FK2QdwpJDYWhuLkQSUkB3rvSUtLWU
bEkvar9jULs3cM0j7BxjRZWceJyu1K12H9VdmuhXPrBYry82xj0YzsS5Fl7hVRX9tOgozLSEaX9B
kgh1XWHurey8idk1AFOCkXdzeSVd1lLduRjFBL4mbSfuKaf6yyJaBdv+2xrT6P6O9cuwRr3+GmNI
g+5di7CmJMlVTLD//Rzk9/bZbf5L5R02HWHRjuRddgLwixo92lD1kFrpdN3q9B+1ZdB2R3so6NwU
pgDkmFRkyjBlFsr3Kvk1JMJ/iMv/OY3fhK31tnEAMd+VuQX0KVEy8htzGufG9xYbKY05sASWDSqi
knVZyaiGVvaGgSNhav/I2O2k5omyuxC1cV9idGB15Wta1SShG4gMCYK6N4XPhLFgbqChoL5FJ0BY
fKMTqaNNEYgWBprd0DiKSwFrjRbgTZRP2DZo4md8rwO1SpbyAJD5LYvkcrzG/oAg5ZwgyBMrLXZ7
hBXEpmsO6nTXaKEwdHb9tSNdtZZtmyVrO8rFB3NXHULoVZjD6enjjdN7eY4mUx7JmfN92dOofHSa
U4kdurYPc46DGlNXft/CisGlkKapnk5H7q9u0REBGggKEg6zwkHdw/UvqAkKoiVF/McSkN1s18W9
dwzG/4r3PTMSsjXNVC2LPIQ1fLeMtJsp35EuxNohmEM9V8L0JeTKTqfhCa7VxzsKPrk7anAABm4K
c3zaYQlmvMOpPzUY/7uIQQ2x/IJdanuJ6Wel/lz6d35PPi6Bvh+edgsaVv8+kSWPuhM3KjWI620n
6gJDnWf+YXD/RTIUAFFyRwC2iKhnEhZfwnEqjJuKb9hYi9kmS7UZ7QYVzZtTr3JewXz0a13G2wsb
040L6Gomiulq6S+DSg8S18Zn4X4aLJ5TrV6jA/j05p2+rAcRswnjxXKs0dj8NwXOvT/dCXKOyBNl
s0Ii5OHghnCE66LJXNqepCmmEhd6i2R2F9KgWv+3igl1gTkDrNdd03vJFuvP2LEeEc+6/hTQ++Vk
DJvBTUqO0CYPWCn8GUWkcKgy3YA4WZ8W/da0+EfPa/RGnvbzYKzo9senCsuIqq3QOkw5xuQzKzLm
4kL0/fiMIhj5LI8IkghxdXwUatli8HGTYvOlDGT8+npf13FRQ9+YzCwtCepoWm54PEvVgiSIhq8T
hh3eVywFlMTMidM5VqdsAeiHsmMc2F0f9fV0T3g7Hi9Hc24DVIeC0MF7nEl3ns1zPpY0ZEVhRCT2
11E3EBOy/RHcRYWbJV/yTuAyLl4iLwnmh5/2xa5tN5zO5iMudHn3QpIfXSt3pebb4zL5Ldye+8r8
mFue7Fahg9e9r333B9phrikpAGNLVQForC2wFRqwNlz0dA2Cto8tk0OCw3bcrq3CG49eWGTv93m4
uDEF/kCuBVlVZATJrB8z9ocWUCFeecMTPuSxXl4gsTedblIbhTIgex3AGGqhq4KDbkebwlZ/YYZr
30mUGCwrzwAFuX6i3XUDmrwM0191tDefINd/MivUy3/ACeOtDLQDXZcBmqCIs8/Vp0qxswL/wx6A
meAM294lSXGXQ82xvClUG7IobrUah/Bmu9RT88j9uE2QDPLRGTHW3jiSE+IOuZmPg0HgMJ/pqVYp
zvSvHOJ2PGUjg6vTnukFy8sXvy9AfBmXpF8zJGD2lH7r9s20dKjPVzODikKOnO3IacwqVgQo7vfe
S2D8IUMScdghtqmZtKKpdbkuI8r1yu+5325U6SM4VAcbtRUX6vzBhdGKfEr3QJ9H9f18N7qeXE05
vbf9HOUDHztbWwsKOiK/jd7kemupJYgboUplLUKR1CoV7hidKINg70+FfowC2fU/HQ4b3PEDmCgk
TxJGcdo/bYCuRshNK4b3FC1vYCVgFphN5XqxbFOddAxZotl1I47OvK1zD41z+UO+FdA8k5rOBVIo
FW+wfBAw8TnGStvlSiPSfiPxgUw5qzRS6LuAXiJOsMU79DGUVIAlZRN9jSneR0wsLduTz1ccOsJA
FyXsJx7c9Ghyh8RLdBtrzilifjcoQVTduLSWAX6x5IgiGMhP+Jve/zoOLhtRfzxZn8NukIOb930O
9lOwWrWqMkYwsgF4PV3QvmqPRnaLVJR9EUV+W+VAzigoLV523tg5lKKpnXo0tGz/LGkhuZPM+eO3
S9yPMEM3Hh7eQSC+4D+Op301KvQtzTT+lqo4iJuKb8/FJ6Al3pG02hj4eP1GUDVGWS+zxa/bRzks
5PpzJ0VJSI0mDWPvaTuzRPlfCHhh0se2QHJ1pMGMWGW9WlUWTJdnpbCk0aYzmROpsP5U4SiwJK3X
HM+tBivxWbqicNbGQtjQp/QrHjBLWx68W2Rfpe1n34zRhv3kDCGRdpKlSmRIwLhO0X59s9HVNtYc
imXDiY0NCm/usx/6M75Bz+YST8FXhqSzyNtVOZTXCCvfLPha2IP8BRZedftSAkoxC8/x+gQSp31f
zpOjxFbjOj4h5rngCFea3UDkiJUYxd5HSVSeRBtK1FAu2N5tZEN4wb2i9TIF8RMxfm8AjCIsZcLj
A2Go2vPppMuaMJo3dtaL2wQO+K/wkSJknHDTNohaiCfu88vKcmnx0Ag0cs/mNH412q3tugHP31bk
kBeNkf+unv+jdGKkt1uwiNYFpzKOW+5upoQJTYiDBJrPXCRaeBymq85j930Sa+hyv69gs799tNMM
wt/AnxamiVAl3ihrVJPuHejF1zlE27hoVobfF7ehNmWFbIiYaaruQMcZ9SGs/5vIMviQaaZcyeAL
WpYn73CzjzAffLay268kNn3Mz4XyklnWDvPm8/0NGjKgy/xGBrwlI1O6xG9QmLzj+v6bFHg9ENM9
7UJN3nVycmEuMXj7eWA31YxOaxAtq5qltEJpagy+E4QpSplmigH2CyCIjNIdCVehUq6N/stA2cSy
G+KrZ4koBgYGbr8bWfs2p5F+amCPKgzyEQn7fTMmO+hnw7CKESPe/mWXS6YDTJ5pn/QiVbN0SK1y
YLfP+BjsvTud7XET8aw4O9YsAclCO4/bgee2643OVdC7qZb1M+65rJjSbKk8ktuGrKV2U85tD9rk
Js6mIi+puw4NaXdJGikfWL3WbfX8iagU/BpN8pR/Jd/ly6grFfxk7AI8mqh2uspeN0NQB/tdevDe
dayOwRVxC9lyM6d/uy3yl6Rx427jb0GpukxxU5nLODTara+OkMewncVcQbdzbFuVfQv0AQboZy74
EwrPnurnuIuhoDwadXchJDVjpZHlipWj0wYyOcNYjadSXpvSSuJojusyWFFyO5RpZZkyAJVHW8UB
qfTcHeC4kQWtvl63QOOiGM2j2zcpmYZ7qwToChHnGBZh1yrQ+u7ho5rRV2zAAhs3ZCJqXu9TArc4
TIV47ZyNwyWyi0xZyTyfZxMd1SJv7Q5wvxPW9WKlM1eWu82cKTnTGt6HXl+rWM/HTsB9Vmz3KDJS
kBZZ4r6JhkXA0Cw1Wkc1ezBMs9FzqTvK77lQPZ/ttpuvC1Uhg6XsAx41Mm9EnCO+TgoDzprIpbDC
s+DsxTlj05IyCueOzUzltkPm8QaBK4vGHzXuwXVtDzwjwRsJqYPL5g+vf+fJ92J/bSH+gP2X0AKL
YK8lyVDW470JEij2s/5ESTNNtaz8WRkRueepg14ftNNhT8/Eb1qmKuYSoqoALNeiL47Vk8T0SvH1
fozUkbfLDnRdcUvv1JfgnuwhtNMyZ7Nyw4KsWo3bv+qMzrwsxBOywBumn66W9CgIKTbaq3gjiLcV
5wgmh8LV1NaG9k3ZRskCytbEUjoiYXSRVMA0KxNTQm4NhrUJhcM1B4+3UPUWFFestXztFmfM26dA
Lhj6JZtDbXsZyH+bQVY2ViSTJxrP5lXOMn33MxKHlAdYetOdAHVme/H5GZvjD6v85VAKBrR1I0d1
7sAxFPgPB4GtL0OvYXGAPWGiX3qv83rasn0kzmmpZ7E3PvoVUjMsYOePMDKdNgE6LwXlRGrFGrJ9
oRivr+gOLUNejjHrkERtjiJyOOEJrxxtdT0GcjzvcG895HRFhRa3SFuccHpgG4eQPFNrblYah4Cr
ZcM05bhVqdswodIvg7Kq21M8c1tMxjsGZItIpDpAhA1/G5Y9CfJ4h/ybR+kfufdMSHSCxu78DmEb
ju5C9XqJuYkZGwfm7MS97x2sHC8VYcmKC2+Uf6ifHxvnGITu60pz0Jp8Skqif0jdg2Ri0EQ4Ev6Y
6GfkRAN7KRwlZlGVAM+8tMPf1aWsVyBFv92d4bgQFIcxEK5L7dQKZo6remaHdTctH7qC8P6D9ZfC
PnWL7KaUwazlPWKxpU8SzjIYXePxb/YCxBcoACLib6bEiwCBj+9AWl6IwGdStjskq2XRBN5pQUls
+x+4jcyzEqksxPWGhVTBcGPCMQY6r/rfHII9KWoy7Q1mZRW7Cd3mp/noFL4TtAU464NsQYysEl+6
9iBQgGLAWfAlK26mDuMtgtpaeUh0x6wssMZDHzY72DttS9Pf0ocoW8ufpJbhYhG6MQhKRuEybckm
4N1QrInRCb8L+cn7YidyjFqNg7l7FGcs2u3j3O5u2lwFLjgdTohBD8CkoFwvtL8p2wb30KUVe8KU
E8TBLHiuCjN66z7aWeweeOksQxLvCO2idZctirlg9Teg01d4AtwYyDM3NY3BHBr51bC16GUco+9U
4JlpTt/upuRuXytLZ/v+x0UQGNPkcCyApE29lvb7AEmUwVwvJyv/ptWR1lSg1CEKz9UVeXAOtWfG
sUi5hEw054c/oLbvW9XAUMVm9ReQtCnVFrcfgh8Ve0l8d2Jhv8d/3WoDZLWBRQ/9w0wQCbe+0aEI
wWRNIZaPdG6bsd+UvUyuTZNfDr2Ul0yh7JtiY/iDdQJdiF/Xhmu7RdP5EIULrQR8ekNnNGR4EDEv
L9JVZi8IKcyjgo68xjJbjZz7C+lhbU9rx09t5G5LwdPMV7XiJSaPlfUPZocfDxHHnXun4pXanG3K
32Maaei2Hm4UBRoXGEHZfwsIfvvFeZXOD3+NNnFv++T1HWtVyGENefqFUeX/SNn7YqJGIrKBQr6x
zgxDAwi++OJuB+2Kl3tDTRzqt9YrC3Iy/q0LfuLlBLiQqlNjEkinZArXnOW6pTT8eIV5CM8jGFW7
JVL02kOoD74Gp9dvsuqEa9LsjtvLXuuwo5CkwAlT9y43fup3Mh90Qeizqivq9M0Po1EVd8W35jb8
XeK6ieJpnf2O6D4WPafrMxW9w97gNNoim4xEsh6frjQb/dfp8LzVaZ8E5nvPIoMdhFTUo9/M3nzU
ptBDP660LYwRyjSYvgP7OdWq/SqAAOrneKsBjP6y0w0E2IJdBlonpe2DYMRNMdOGIYesW0fDsAWk
83GnRzjqQvwzDZ5aXblFJ+iLu6lZSfOaWjLYiECve1+ldekfb959ogkC0Id90MVx9FWkLYo+v+KA
9E+l/jDjdwRBgepOV+Oi7lmju/HpqB2fRxa5XOedwiXldrX9wRpOQLBzuAJ25KNdk3gT0syEMIL/
5tKS1tzpr5LIMLDtANKnJQE575g1d8a6bKkvWT146igHyy28hoIMUtsa3sC7ct6GrMXsWDzn1caw
+ODnW27jNwve/OiKnh8GND2spg6XfI7/2OEtcu+3Qgvhy3YZN9C2zSff3szhRmnFn6NvmgEHBVMM
O75SX4WumvQN8uwC+Xu/nMi4NpL2RmONP5Qhj0uM6RQUjghtPKlEgu2Hlm/4TJoT0hxPgo2Lp5IF
AZxZbZab5xnebGLQMHIvp50iyQ5v6JCJ6ungFh7sPGcGBNLWYxT3Pc1CGaWDfaDO+H+m4z2hxu3P
S0KWN6WTLbbcrn2EfLO1wSVS9iw3Br0VlFaEkIUZen3lHFmj56Ij0eiHE3SGQaZxJY3Y1qfUfIN4
gsM8VGsD6dMy5Xo6i2/HgmC/gF9UQXT+2xbI3hXbMVrjdUg0XpPG7lW8Xl/elAVSUT912FD3hxmU
XEBEbRaa3ihyG9tp217fVaHC/ljTr+6e9dYCwsrDwQGPQvgVK7HZv/I/hkse/Cl6Ulbg5xHNu+aR
MrvnmRYAAwA34YJs4KnJxRptpLK4ScHEr5+4Yn7zezSeVcpkshBzbcas0CiCD7hWf0oSQYh0lnLC
PPACGrpZAjfnYJI28+GCZeMsx0e2H0OA+LccG+KXVAttSf9aktH1rRF/SXqs7bMWJaHYDyNxJOea
BfwRbci24swbiClHNBl6GUjQl50d6DcYcHkxlW5kxfJM2mh9pN00cOwMhGKjhc27tnBVf6QVVR4o
e2XZxk0j0VxM0GO1tr2/J0T13rdDeEfSpqrdb3iofvFlgMoLfwBdEhAamuEktjDPnzXto/HHBcbt
MzIIBKe1BGP99gJtBOE26Q3irJn/OfVdz+ERnmmyAAOrQmrRjorvtfH5RHA3vH/JUcK/euG3/2Pf
ckx3fKfO5hPOGXwebNrpL+bkBnMUGSJYxtkekWyt2KnSHbAFzZSIMaaIAxq85wTPxVRJJRDqGJH0
sNodo/Th50emq36Mbhs+gWPOwOrj4Q4IBNNHXzIVE9xLfA1dfrg0jZNE+Y9K+HIGv+SWcW+AfLuE
+KfwllDmSQMmjE+DY5h6YS8sqXm/65hZ5fNu60jPXavgQmgtKOdX9o8ji075GxvWB6nk1nxZNIit
CY2foN+qy2OyONOdF+3161GT1Eu5fsqsDkKeYj9g5sFbTKQEJ/p65PRxKzhz0bBCO1PiaKh8fdkF
Z7rYh4xVW1g5nwLft906hwmuoIJgMtXDVPi70ifVzbJ7vUx78MeAKApmXz91rS/MGSrL91NmLSmi
TSsNvlH15nBrbdpWxb8+PGCeCeFHnKaplhd7e7Y52iiBChJNZ5RQcyuLxRyljbJ82Na3zoiSszJT
T1+MaQb82gkpCJL4FmSI0IjCQkF4d7APdnbRVYHAIr19aeKTlA1DhBgz2Jt6NVG1SIKleKKrRRb6
RSDPBG09GUINTq6gyv20x0Rge4rkIsFJaqAOr/G4yxrwyDrz5aBC7lYiUcUNaegu06Z73gbDJZ56
LZSL/PmU59idwnCFrQzDwdYDMEGIJ8BOeDdaDfOtNhvVauEV9iSmjl0G7Q3thvyqhIWMY8pji9Ii
4KD9hsdau+i3VwqY74iICGfn0jNxYLX7sj2R5Nc8b19ervA8bNe53hRdkf5RLLbIQaCXx6QYa+or
5FKp9JrVVPD8/IVfKwYi81ZCndqmSFY4Y6SgfXHWIYqIi0qMAqhLTBM6i7DDJ7iW48eDvTn1zINj
ioUSO54hIqGog1bcm4jF8dFhQ+ujAq4iclWwg8cwAlIJJVgDU1PLquHKbY3wmge+lSrxjZP3CuPg
xjfRrVW8YzYka2OFdmvsd8HnhxUpiqPg3mEdAUQBzQ60aSyg//JSKB0ffhGqX8cgtDcr0saamNsA
LFNL+BImmtfkSS7j1Ytna9qBwsh3GlLmOKDrRQ6niiel7z4AK48wQaqsqL64m9Z9QTF+1EM8NcMt
ZcaE3S7x09RuHpsbkUCuAFPn5ON5WizsJ741Jgod1d22QJ1gLbTJwu4SiMstfqw0oNUx9i/Dr93F
RaALeyntjMe7hVNQnJbSr57sRzjr5KUtGiFioTaBW/84uKd4qLdqNlEAJ2ZxhSRhDMPL6up5xkb4
COSWGKbF858WbFgO3UGFPiujumWzz8PwpH81vvNT2C6wv3GXq3s2HESXekrm8CeaWUM7FkGT+rd3
cvUYxjdaIK8WEwVLFHvGIp7qHgxf/ZplUZFwtyDB5yBGfztMmqb7VOxZw2h//UhmydQzrvIKolJO
vBct4jZsAPo+g7hQKBJtAz3dQ3imGtaUvRRK/iEBy3lxXjKvax0qHGL9uJBwSAlWD5uNQQBhy94T
lF2oywhytZAaXuyK2vMkr+mdZIsK6GnTjorgaaCDaM3KQKCdvZ2zL1GzwSFXmu0nUnG4bHBtF7ve
xTNNen9meFHIcgVmt/xd/F7NeVIwwo0NPadpSQD70NK2Y2xfbnaI3D5FC+eTJPZ2e8yIzVNkWaAE
PmAyAPeiSBt21oeaIgYn7oRgcprv4SqaTskUx9xAutoNaDXD8nIPnhFTdLJUMaeo3kSJc5q7kR77
hVJt2vIkTvhbS5xCfBppxyOF+HXiRevHMK8sCHofOf1V1eDoWNTzmfhT72vXdWs6oCahBBdSkS7c
n7yBWwVi2W/OGgzI5rw8IUTxG5hTZojdhSmHSoURALjybqMyEvczoS6WpP9OdpTyIwKioAf9yXEk
ZbCu8JUO0Z9qND7W9s7gIyF56LQ6t/qjiP6qE86ZMXZGQ2X6S5J3QdkxFFFQkpwTQorMwXv6VZoE
Rn8HDxL2FMWeH5p/LODZMakQl/BBzMBWOm+6/Uo1fMUctA+sK7rBsWXBoj51InxM6Xg9SCk3plLH
/XzIrOj3rhpNcw2OeVB153DCAMrpgx7VjkUTD2nHiaFMV5E2M1cynmT8Rz2dJc1zxYSu0c0YRbwV
urQ9PN20OMGPBiFAWkbTua13iaqBmV7odlmhlebOe5gC0mzkW6XaFHijOPVwP24A4MGwa2nduhUI
Gj67tsHdXCJz6R3fCirqVxmKLEHUEXdee+M9Zvm0qX/bQbDxkIckdzANqVHetPsqG5GgqX68Sab2
Kgqgas/XDtItafjnxGalAuDxz7wGhETJOzeVmBHJIVp4lJzez51wRmEcQxiDOAWZyOXUXTz10qRo
SObdf1tYngX3Q+MYU8gUSdzJGX0jsrL2MXZX6quuD48kDGolFHk6dR0hpBZ35x8NVgzrziZ32pVK
wA7Xvkzcp96Krz1JlIIPCO9UI8B0v9qMVbmax/KQuMSBRCESMP1NkonhFs8h2+g+vhEfLAkZT5Sz
mpBaI3LzpC849h2I5ZDCYP0UkCU2Eooh4ASRMEqN8WXRjLFcYv76XVN8uNYjN+5ohTNQ/MWo2q2j
YmADPPHO5eEsS4yzRnwNL73oOZFqFTG4iXLYmJWnL+fgNK3zO0L9byOW6L2xSrokxMAGJ99heeXr
JttvfzIkN1AzwSZAVe4jKWa48wGuywuSysvHKgMYryivJjQIwM7iNxV4jslnSDYJBolddL9VyT5O
moVEKWhbx9p1/Y946pj6CDMgy7FPl8d/QZ7ptFw9EjQXudfId+V7pV3aMIY3vG7cY73RiZTvWUcU
gEHJ/pWqKDDYfmL0OwHWsiI5L69ReM6w8txn5p3LDaJBGCkN8zRDqatvCd0wjeLAFJ1RAC8i34On
n/MzQ8OpazWhrpPuGQXfOgllYrRwoi+ebHNHVQsIB+tetmBvupOkMhADHr8o8i/5gqwuHj59z7BZ
XGI7UOy9eaQMb0J+qg474bhDuo5KBLvpnRpsTN0WjWA8UyN8u0bxvtqZTuurI6ca6Q2i2gDIf66C
S2NezFvOq06xyuQUc0hWwjipIvx0JEi5B44JBND18Wj5qpps6+DIURim0rANfuYvrqwwndkiDOrY
P8qVkxPxHKBAnB+OrTybXHX1cymxAZnqo3amYSRxuQcxMJaj51O58CB0CZku3DfiSdzfjUG10RlB
uiIlJyKcLvkGkywrEF8ALw2f1pWT2LsZwB8prBhS3nAKEfFsE/qt4z5ummbHLjGjgPRnSNAFJFOY
4NdA9tDN/1KIJIimtz91zn6WiknrC8wJQB2i4oIu9qKFy40bbObiZXe+eP9KqwhtoI/fRs6m5t3x
JyXu12C2aQzBRa6m3PCyUcd6uGZdm8pPMVTDTaOoCbPFJnnJa/J38tpsP77OSkQaCtldQogpt2NV
pDZmTQsPmkV4Oe/ZUGlW3M1R56NZr3+FfXidCEQinFgOVN3rQq9UonopDMK/xOIFgVRANOBHsY+W
HpE2F2/bG0UtLn/wcg+7u9xhs0hjBba9i55hBZoBgqhrf8vr9Q09NIN3MWgZNckwNhQUT8hiFDPL
poBoCIkJ5j6JE5F7SPzfSi6vqOqAsNNgqn2fbVmMM0LbOYsL/LjBtm5kXd6tp1zAgp45gp3wWLdF
pDTH6yioI/2liwqTH3MW3N4PYuf5WzXEOc8oFpXz8jCYUhmdnbJki5jAvgW1uWW6BVrz1vbPecLX
QSIhG4lM6c7AEONwEBPJV3aKtCF04zriwqhfhyiOCkY0ekjRI5WupdzrzR9BnR7LUYzv7JRORxl7
QJ/WHmOTEfMj2mMnQGrHFvWPRfOeSjhQPwbLq06ql+wfyMM1ittxV/LxeT+h9g2/Twbewj9sv/gz
CL7Odws8rpwjjMSgg9/rZItgBJX6OdArAP9f2QPZwcvcwV1DcR49qOmFNN38KmkOB9dQ8UFcXIBr
8KqTAf2EVZXcyGttuDeDFMCKwwJly/e7uQb7iyHa/tsDMep3+DENvhu9acGfg209X/TcSZMwQP3Q
Vanfn1oVxwHBRYYZuMfxiXN2i7QVeldSEHvry4PpKJPB+YxEsYmfm5dO5j6dIT11RZXuMYeqA7Mv
jsG1TSFq9rpJdWGK0tlwKoiuI4NeTZuLhv3Sg8KKAd5UwUfyiRKyVJ2uoWrDgn0iwYgZOYnTR/R2
pbO0dnIf1ATK2tBuOjNEHxrkmg3oh00MQgr8b5TlXyNez3GD2qif/G7M9wHJCd4c25BADBihB2dO
1UztWg7CoiRhcKT3ZNbo2Bje8IHU9q0HcmsVuCZ9DC9H0U/uOjZsrzOQJgL1dFQMfvnlSx7OvSx2
yaBAuCZNat3ZuHA5bTBjSBg1K+kZu/3zR8j6981Nd2kg6iMEsKELgZjhtVsY/ctxPTpa+oN1D0ui
4C19ZQhVsQ4fCyz20tXDLANgQ6kSSOgWp6HemeVO5gvZo9o8z7Xt6aL6suFX3ZXO+XgASM/gzQky
NAuKa+uWpVVR9OO1hl6TB5APWUbo8Zmov4IlyGHSmgB+fGGPPgmF0Lulkr5jvHf+6f0bkIceBcMR
B/IWtjsTQcmU7kfl7jhI/t8yEpJENaF5ZliX4qOnFqQIfjrjEIGUCkSQ75kfjPN3w6xFA8swRrVt
h95m2SrJPK9VQg45MoYiLWn7l5fVHYNpEwDqdgWH8TO8EdycluUxpYZuOtyTXfQ066j6aZX9WcPH
jYYk7wJiZNn6yyPw5SAfo05PbcHNkn6XuDRwXSarlBKZUEgFdH7HGpWbIgMrDvohnRRgvyxLm4Wn
3ZL8FnclyZsLXyyYd6DLmntlS+QDsJ3CdmwnqMI2g/0XKnKhbK7/e66OBf+xPDUNA5BbcZJW3IIr
VItp6wyWVs/PbcwjPVFdPGKWfowfjUqgKuiAaijSA5Ce4MAgOgLVbcop6mubJOVvIwerKtf1BkGI
iJyo1WI5ytDUQZleVfkFVLxJVkFDCZdCGMJRAqWUhEUGtgttCVPyvEFvicnBo7B9h28Nvim8vyBQ
nILE+FwRYTqfY7oMxFBHzVFfg3Uwn/WOPiNKs997EytHl87cuxeNuL2/n8KK7T4vwQAJegA06ini
1F5ZNI5HXdflxEVMQx2/qRNCbE+9qd9UtaOXOq6E1NlR3eXN3hhPehoFEjR3SJoU19ARLiItoiNJ
eEBrtYbq3Vou6OMW7od0mfiu/l8CDLVlzjR7sjlKQAD4YxTBQMqdg00koMqaFUXQF9n2hBaqPUZk
jsouoqnjreQ9ZFM1+itk37G7nqXyghiDGt2cxdEk2waL+aEwVDOGcXHGwJx5afuxq9FHMjSQemRk
IAaJ7x8CXFmn9mCo3JqYjrh1DdavT7unzuOIP8Lx/NCfv2VxXF3APZ/NbU29BWc5cZCDnKCHMlu4
XnOyrEdgC/i2QOi5Gyei6nJ1z6bJt2ueUWWOe3FFIGyMCKW87f0w+wUOV/W0GoIIZcN36y/ksAED
ZoLaaG+J+0w1XRchbMPN3GczWwaYQqIIP3cZ0a4aTK274/68YmP6IIY3kwY5dkeXjkE/JhUIzHBC
aJ2ZVLj0iNbMUu+1bSrbSQj8+j/0xlOWv29tU5qubQlqanjQyha4I4ITUNFv+g1EPYou0G2x+s42
03jGfzus9jXgeemuKpmPnV2LI9X7JkvJNn89ZdIKadWuoZZUimydBQVyKlKOKLYdyk14AH1UK4jD
ub989DsJYJohGPICRlvkS7kNOCueFdF0aJZu9iAJnKE6+DUW+8kUTYnCZMrZSQD9MuNJMKRgF+Ef
DP/DCuD06uoH33qoJ7vhviA5OHAhTCEx9DGRCuFLavR4ahhbT3YaoK6fH+DkPFyTCIJeiKWuD+Su
c5Yi/m9hiKy8Lre413cZaMmtzicJaNOrruRgDOaZwcU3e5iw5aE2vjk8R6pmNaVZDUzlPgv4kNbv
s0fyN+Ju1al+WcVNMox0uqc7P98vE9Kp35S5PFW3ZE21xWYda4pyLYeH+sI3sda1WW15T7icIFpA
ABm53O5lxERMvuPp8c/39myG3JIp2fYjEpVTDAB0G4tB3K1zxuRTm0SSITIr8NDOhXl8Xgv6A0mG
PnH/U9WIvzEGQLa4AAkhNdyRiQWPF3CsshNFB6fvQPK1S1SteS97HdKwOcE/X07oK6fl3PzTB8tb
T50NehKgnzsfHfcwEuEM/rBB42pjgVP9mlpLzXPLsyhZ1EPdHzBwyjFcwXcUmQsPRLax6KXOIuQS
zJ+1pkJDzbDnVbb2QSsu0MHjscmoI2wydwKfHRBwK0Tb8P2CEo/fSljRWGqx35w7gYublZj53uLe
vSXEQFG2Ihp41h4SmM+WxMHknnMSgUTWBaQQsWNDcyGAwfYb3SmdoDAM5UDrF2S0ZnqfSCPbHjGq
xIxKKdkwl8mMGXOx10BrZ2zWXUqIxSFuJxpReeKfnApF8fzib6jiEpg1x9jBDGAlwNjLjsUDKP3D
y+AvIYomb+d5Oflk8JGQ8bCt7Qf99+qZsQgFxRsRqvnLZr59YbVIE3bz8CqytuZ3yHL9S/yLxYH5
DgySPFXpdDwEgNKuaa/bEox3SI8STVigfQNmI2lTvYtuP+XWSubrvIwP2fGIJAJsf0KUMPIlDe6H
7O5SOK+W7VT308HForYy6XspUTTI8hkMH1MqGsAhoc1EsNXTemUSiXExc1TjtFzia6t7Lotkb9KT
VFzzBS8AUqWJ6IgHN5dz0oib/ozfEAXBew0rIUw6qjIQgfrmLww2AhK7GFibtMVef7HQkljjfWTz
e5LMeAQoWKPXDHu1TtlinHlH1Hfy+Bzw0OwcSpGZFTIsmxpHhI3CtZ5pVAH/hKxdNRnLpLVrNBGY
GD0XBqpOgtVjkucDTfOJgmv/4BFQUOi5Zbmy69lklXUzADQ8ZhNRdoHlXjv2trW3h421UulgqDsw
kdPv6LhcQySp+tVaIKXHqpv0lel5N2Dhif5S0M9JY4WPr3sBuW5mkcx5jTWUGEzW7PASFIHEwGWd
O6kOnn9IxkO7g4s4gKdz7NVCOJLMYIAz+Gr8UHrrLXWGwhC1Dzkj8RQMRnfiSAFGZ4E6cGqqpbCm
2AwgzutaZP60l6iEh87n6zIGyIHQt4aSfKEGPdKOvJjIj2gVBjQkKXVCDqCd2yw5g3aNTqqkNYPd
wfi8i1a16x52XxjQI+IWnaKvFWx5SNyV4UWrcEmHJ97WxCbl0znr/FHbih5f9PGwMXK6I/m4wSqd
+ycvMJG8PEPAoS25OQZVHzHEARJI66Ub2teYYfOsqevFKUryNfinDCbgj0tz3mVm8vUUnj57upMU
0MmEFE8iXIiISM9DFGmjICm66yzcuNHxCMnWjFlL4EvUPxBG66fv2r5iFZTs1WdD6RPApYKN5TRb
YWds6Xs4aXIAeTQw0F9V2UhKsae1/EBX89nqtly7wVT3ltRCKv7ERur6ZQZgBWrjZRDgG6Fwg5HG
RJa687uWvrgkgXlvxGKxjv/exhiDniZsJDISIxOJ0wZ3q0wIgi78/07VniUttCPjsWYqdLX0+/Xe
bneoMOjzostGpLgG4O9r3fHr4x4qMWaByHqDE7s14IEsE0EdBRLo3mSYU2gAjkMG9yU8vSO71M9B
/tRnQ41/3HbfSFHS1h15y7Ded21qXMn6tgH2cmvEvtmA1v5aLmtdx+7JcPBiKVc5FQRzo1sCV0Kr
w2oAHdeBVSUIMZXk3Vqpk92m2DEssvrvF7fntJiBY1DfGXf9k9mYviYCewI1X8qXmC/diGl5sS+R
9oy9Zm/oMF32IrlnOp96iACYJF0IkHPWs2Xag2mY5mzwadEjkHsQIgsq7onfszemqpj0ppnlHnNl
bJuJ2eT1exBthM3gP1O409whgJTBJv4GR5NsequkNLwgnK2dl4M+p8dZvkwcqmKSfYvycXKFFtd8
xqrnrmst0sapKHj5//zgiIKqYry1/x2g+CgZg1ahVlJ2erNPckoxpqFFxe2v2KU564+ILGEhhX5x
AYAu9NNYxH+KU4KVssyXW6lcbzAWZFzUInOa2/2ntt4/JIu5F5kVfSIEv/dKDcaqZatL0vcf+WZX
5d5ZPyM4+jthverAHTFzLo/SoJB4SR91Lhw4OrqolnKZebP/++SE8mY+kgYazrv+kEfKhSI/RkO1
UX9yraIvtk2kZppmf+/B1wNLMpJZPltDDscFlNsateCilO6yt5dcR4gD+zyZzVsI6QYqkC0KLDDW
VpxVx2/xMsQa84LxtI4fAr1sXbt/Ju6PXY9584tx39u81SEphYsYH2kHjeJtwrIKApckIrCnww5h
mmvyWkL9c2UHpJjmR4A+5zh5K65Mr5vU/N+HDRRdhDrO6bUcU8QgITSsMSoUXAzKWbjzYWHxq+mS
QZPCRtj8oDqbM195sAKkcc9jB6EaAAxqQAZPbqG1WudL1OH7rwLmxnlOoDuAyTtgMctzKgS6K7+j
0IpCiinUOsrS1apuWg9uq7O+jmUoNYUxPcawXBu/yap6iOMRayIVIzdgGoya/Cb0Kean/cCt427D
twCQHXSembNSlGVAc6XFEBejlewkwhIhA1pe+wsmYcO5bObQ26IA7wsv7XRhsdzllaCW7IWV8Gcz
lgazkGEKWKF8l7wQi2xw3wpNYPGRlxGp3qWFIRtl3su/ByS3RUKTkchi5msqrqZc9/cfbl8BWrIC
RtVAjQyHeDjlbMORydGqUwxYZ1q3ytnE2wughSoaYFAxCNkgbVePRf59ekyT4y8lCOVQJkq6a3XJ
AXASz5yI3ABOrzMlmg+XsroRjPGvQ8eNUK6pY4ZkSSnIVAeKRWHetD73lxMB3NHhfoyy3zfTPevu
yj5kC5v6tLTMtFYy8qfdr3dMHcym5J4H7DUpTkWNlCLkKbA5Ntd3anfRc/whLmlm6wC+FaFJ+yRX
LHqe4pXtv92gy6Z6FGs9LmY5qmL78CKxsDz4znY2inOecDive4dY4TN4WqWfexH+8WNRBH1lHbsC
J8ZSusyMaXI6jtMO66EATt3eGKUDZ1sfs3NG2KhshzMfn1YcsrFj+ABZ0f914drUe45UAO1BMkl6
g5v1PEWRoQdB74jIphKGa9Pz71mSdXa9ErtSPlauOvJlp4SIvk8FiGUc6Yq3g3GWYQxftaLUjqxl
1L6CTLMz+ft0hJBeN0HT78vMUzlbCHkM4sXAXimJIqzOXZz051qlIkaRJEFSPXda69XUYkcmYUyv
0gGAgwTJCEibvbxuhB5h8j6SFJTjeiEKfNN7PSYieOhlHBnBTB7GmzzYvuaa9rkOLv/UxSI0E9/Z
/S6H/YKBOmy4XlrmFeQXrysHm8oNBexc5uOFlW55ePyac6W78dj7B37PHgE2Xur8wAxI2faZjU6/
Q07eztrlujaw//KzHgZZeLGQ0og7vVbSffwFxmcF0sQft7W3jXLKgLx4kLUaY4RH2LHigAJDQsP/
e5l425dFyO0CuGN8zZ480suWK59+L7qcPqqmSPTi7zIrLFNeY7K1hgUgN3PyNs4aBKm5g2YLRcSa
27lR3tZwUIX8hGwOk/7fTR4Jp3E9LQmtGjfTQLSdWSpuhZ10d9DSsigrUYI9L8doCJPGA+sz+Y03
U+J8H7BK2/hT8Ctj9qrqjnpkM05i5Kz9gHh5jhKUVDNdcvNDlt8dOm7qMiYw0vnzL0ZpX9PgP6jl
CTtsmMKNne+UdctUayAJpqSIUkbFEujsATjMbM+UFM6/RKaghkY1cyMei9SoU2RkoSq1kyU/Iwm/
n7NABxbsUVQbqQxMdYs18j/r2MFoLXxn2sjvNOF+kFegw6lzY17bijLqjG0cXRXhCTGjgjR5DigC
KlGqhvIqUQ65toUlzaTIXklp+Spy6hMZKNqE8j44K4dWv4kQ8qFYKwKxV/9OiyfKFJxsYrUCoGGD
I0QqiG0Q8z+2UvVZWQcUVcWWcD+GpEobr/TQbnoUpDRdcHnbX5+TSbcRficcm1ZgF+xlMJRyOaAw
y0ItPbDPwE2JdMm/Ic6GUcwcJwsaeOdRW9VG/LZYcE/uNKhm4JfLTBgL6L5RhfBFf/942qbNIu0r
tfhgZpeFfkYTO+3cBsJO6ijJ37d2eegLMgKKFmyoz5mFSw44+z4uzYH0DV3oHPWzet1b+RvCQB0u
X2Rrm9Q4MLlUgGT+9nkSgyGsPKmZzAxXZWBXn0opEvdXz7RpbQlhd8TTFYyUJAJwsb1iWuStO4f3
W6jxS0aj/3rsi1lQDJLUFEFHtp9Cd+HoGBpKP67jn266UrrJLSLjX21L4lSZJRe7VIZ35DkfkvV9
QeLW0t398mPxrZXiZLegR/1OYBFCpCi9oaz1XRmYDzibAgetyIMZSJgxAO2rfAUME3qcHYQewnFA
/zW8SAL5su/4/4Kbz6WlZhqoMTVMRDUPcO0AVGVpOwmQ+KEDD+RvfOfhvOMdpKHmz4nJmcT6/yYQ
tco6Fk3AJq7IBEjxb3NhSTQErRVuuRDIZGFey+iIa7CGNDgohP1Rczn16oWsllm+7vetBu7DwKU7
UeLkNea5M66JiBXb7YfGgqgE5zVw5bENw2hcL6buwwlV4+1HnHsyGBgWhh2PbLoaUafIOyHSzwPj
ClaEIzp2xknbGxEZtGIkOHJ9ERfzXQTi+h0MaTNx72RiIHI/9GR7xLrAhKhmZrHcH+pCSBf6drM1
ur4AqDpM8VW+hxX48JueT9k4F//fRMEbV2dwV11lqaqERD+K8S8lkntQGZp/LQlOqVsrAATC/lgF
Io7kSHPh4sD+kEZW8qdGX+zA5o1m20R59BpxSaJTAWtnUuJOcXd+3vgnC2Z+EDd5yQl5tvqSPcmS
YqrcKoxwi07RCIlL2TmG0WN0se6V7ZcpR9ER+MnuNYm+bVMmP3RAWnERdyv7ADQQOm43E49XoxdL
3FGxPMT2RpG/nfO7+UD5d1/+hb4+GGWAcEKqCygG6TeBXr1mElNBmPKMDm5DpEisXS5fob0vZobG
9o9DtUpIAqtaeh4bJJr5KDF9He3LahL8mVOS5wAnjMY1xrfpxhTvAgqfaZvK4gPCmcURsc7k5VbQ
Vd8yfSkHBNfRvr6H5YW9Gw0++DsS7Z7Yw9u//HqAt1mitADK1IBXYtGVgg0P6Is6xF6y7gvraYu2
dURdmtHSVsuzipcPweYNzzu2VM3vLYC+EyBeK1csrKdHyK9yYK89FZ6LsyfUiKJzAQVkuT2sLEZC
68mkKMMaNYmhn5Q+2jbSsnkVoO5jQwMBYFe/AZjHNnNew5NydJqerO777Lhrjhc3GHnhqoCLbIeZ
WYNTj4lBz6K5ELGGVtA1g7K+GYpQOeFG6kKsuDrQEeVsTN2PmQIEe9bsQWdiVIZdpJkV95uaLBIm
rgYMx0veQYB6H+wsfYnh6paj/Tq3UgcW+KTh4DX7zgFWmt5x2rCnbm2+FAm9hSa4yc1br8dmxbUL
znmieW3YUJWETIEqcAC/+qXEN8W5/N4rRNUvGstfUSgNlFITbv8VMoweA6vZPy4eA07d0/MhZlPw
CXgmi5SAr6qppb8M/3vGRos5UXWelzIyahbbdmXKNqULqW8mV5mLm934gEbt5DRbrOyaVUriwCDc
Jv+NO9xH4xnq0YvcwiEpnxaPymHQ3/XBlGMUcRbYWz5UKaWZnchAxVg6leK5WLHzX6FgL4pArqjM
WlqY8qxUHObvNhDoQvm02sYIP/u+SitYMxz+967vOjue8BTlHEQvj31hWVhicpHx6c15ENm1kgUm
z8eDcrW/9bvAAZUJd5D9McuNzaORgMOsAjzlDhAEwWIdhhiooWgx/r9d7X1FJVYMRvUa3ppWBcMT
YXcdsFBFHkpH+LdgpLegTgRSds3jsW0+0hObOZodu293J00LLC6+Sxiv4gWVtSS24T4VOmtkWLS7
IAQ+qOv8SbBgqxFNQjLFnWwuihhEEnAk5vsCaSmLSqQP0BDioG2CsKCRGwp+ZonHdvpKI5N5MbAA
LyZqqgEA+pMQATiY7s9Co0jtcD3JrdMSAaub+arybP6lKfz2e2+tKi7lk2ix2lDuYuDVZcIqE3YU
UEnjA2XcmRivbbNEFe020b2DG+LSpr18d8SktSu03xSbG1omAgjX+kwW0RV/lfz6DJQ9uG2kLf/L
lFV9iODF12B8K80VCozr3Gpgnht0XMh7clTJSC7rSSlgLvbQaCNGotAYw+kqo/9NWCOQTHV7vYUA
2cqUz0X5MxeHJ3+B9G2fasQzHhFseW8HQa+SVG1nynN+U1bWYOFCtpcBd+xRxjZ0AM1O1GyTIlkT
8updSBDDhglS0BEQMgu2dDXRUg1VL2X7cJGDmekyka6aUNSRsrz4xp+HqL6Z3UPe4lDxqWfojzl1
nwcvEmlSCQAAxNM9iFLqEYcbw2Ps9TjkCJkycv6gK6MbwFiyW9rknSBZCOGtiVp4iynoqQtRvOI/
ec6gQW29qV8nMcGUkL+0fq7us7CzSQ/R2dIeFZZ7pjUC7joYC1J3y6TIh6LsrucDcaZ4QiP8nSnC
tD2B/NTn8+9044NZOIGvYDTl0BNDTlZrCq56tBcvtbVsGvINoIUPIRTSd+TCxbSHZ+pj5buFUfTA
q7+mt92cRR6MADz2P9OUpQzuOPVBV7vsKoLZFAkYbgHKour3oTFwqKpLvjDwjJOrXYOjANHgJAPo
g81RnW75GElkA/wxtEFqTREdd/yKcx5KhpiVlsvAxcDNjOoOUn3ASRhFI/Mz1ozLrGOpcuOOXidR
UC/hngOL6JrbgSf3GtQm/miBJHrc8QfZlOjhnA9BOM/sgpmhi7HjoRcJN/IkA82bFoyf7hzGWgi4
dSJiVs6QaJuBHnmqW9uNdUiqlI9xDQLo085GOYDmitEHNE0XsqRcwuPKskiz9bKuybx+aOCkH2UM
FUbK5cDp0mv3Q8R64b9BcCW8cm1xe92gv4vB1BiFzjxE0rUeYUNLvdytiBf72O2+Jklrmkm+dYJt
w0DRvXZrdxS2+fVglrLGXH5sjX+0kXPs28iB4S2+Bu98VD1BpUXdhJitnNq7uratq3ruLE1YLOA/
OrbUVyCMnxociXroYBX1nqhryDAkgBwCtp6GNF9ehODZjuhEs0aCdOIv2cMIn7FIV7ffTla+Xtru
H+UxktphcsQVD5pnWA2VU0YSFcB/Hn9r3sWEjju1jm0LXMtiIt1pmtV/VT+TyBay3uNURCLFntOn
EY6IKMdUWCMWruZdkAcoXoRPm8Lr1vYP8qTX6cdhbkKSlzBXdQwEuTrbj6h7cHO0g8UZ/IDBw4+v
YsHoaoffp2eHXdCF0wNRTv/Pv5jq8Km+Owxf7z1bCTJYWmArDbhgy3ZNd80R2rKiuZ4qCmryDKUB
u16S25GG5RDy7DBSJ4EGQ5wOWlDOmnJkYWxecyQpbdWWdiYrPhWuRLuvMBoI7gfxi4KE7FwunyYo
CqlFqvtSDN76r0ap79+9Q95MC9WbXu8bB3m76BuUQhP4bD4STMWNYA/LdaxDe2N6lP2q6IRY9vDL
sp+W6jQhL+tklVO26kAFciMrdCNVYVyUeTu4nkevlQQfMjz7vHQY1Tu7gIFvzQzeQ7CNXhB5iSMm
eVaIkncO9JnoiyPYZemj/13zEW0obKOk3SMpZk1RABR+m5qAzsnkllePTfruzRRcSOyOyfuwjLp2
bYXduNXKeJTzmXnTCybBQ0eVgmWP+wplD7Ky4V4SGZL1teKwz1YiSUMB5k4q2F/tCcD945CHE0R/
1EL/fpY+NfYyzU+FR8LQQHnZZ2eRoiPDJgZbXYuyHxZPeaRBhiy9IuY5NdzmOpBJ93zkmYMINBST
ZYoqFtpCRHeg7E0sKox810sfMxn1S2rzn1Br9RD6QXil8LNrXz3oePB+85Dcl40B6ZHUcCknScuQ
+LnvYNwX0lkYVHM8pVVRDdhhrEIkdORcWIEghHKuTDWQlk5JVQqfS1d1a/s5E7gx6cT11fySjwaa
Gk68Nh4mrM/JNAP0fjseK/UgzEhiR4L+/yH1iQbGCROWT+CCGfK1iRODki8JRpHQX5wTF522+mmq
ICdiXvgk6GEdNk/Y2hdomgahJ0pJx2895pUGe51rTh8x81KK8I9fKFjOqJVs20DtsXaLOVLZ0JvL
N5BEOz81WEVFQk8y2nqfDDkUYQlcu5bvrXAU0gezhAaUzoLL/+r7/Y9MAvcZxpEaLM4J7iPMbS35
nmL9NQAx+uuoHxQZDNGcj/dCyHd3yLtJeCX2FeiHerL7e6+Y9PvRvIbOuHh4fKwr0EQm+sc5jnFr
3howtDaEQOur3SGGwMkcZazqwWVCnAUJlM/IrwU6+B6tvQIO4yAeM+H+Qk8RmQX8GXda2KicEjX6
iCtaowVtUnqV0Zr8VopPOhOYZWxAkU4ydmrj8XlHFzTK5EKyy+eG+ZgKvva3wZ+6aNpJ4eo/SlWf
6BU+D6ayTj5AGmrIXmRR6qzt4QZgNB87FePbJVIbo4AZ/OnExAoS8Vvw/gPSmWgDB8sNmZfIfyOG
v/FsJNjUbuazvbwB2LEAtpXldszOIu4MQVBOFzXL7AVG6BR4HE2RUfhhAq5vyGnyuSiQmvEkap51
pB9DWhMBqzzhPFcp/MftSTTZviZkRxRsdTvIqnMN2J0KieM/3waUvLg4G6jFOLDj5Ag2H+Q+EtJt
1oSGxw0tw0ICelAypnZ+krLt5aVnqQNTzFn6tKxD5gMiVzC3T/b0FX5tWMcMASxBziyOUVnD0F7v
JpWq4Qy5Em8D83O476sORp1neuT/UQEExb9cFqKI7erP8jy5Y47zXxomakqxOw8B1Mu/OXl4RNGB
qhOth5E/A8XVrM1YX+Y3diwKmDtFQZSupG5RaQzXuER9NE5enmXutothupDZU3Zf5nJMqKG59+h7
jUwnFH1wvP4Cyk74teOsP0/ZWV4p8RcjIrd+UP9pWoaajVJaeXTWhryBLJdWQx/fjOA7isaQK2KJ
yGvau3t0jaqsTZM7HqRiUSNatnrXFCs/biVQSFpf/AbsevFnChkYym/9yXnFb1WOfU7dBj61mhp1
fmUfLbd+SkJEovoHQWWlkBvL2i3wRRVJ1VLE+7GMhFpK1EGJCQFNRtBjEwtLnNMtHi9M8+HNkFpE
QHaTYR20Ut7ykPIEyu5IOd2w659Oz65M4B0ZO4+TTu1ri2l3EUI0ruCekf+EonbxxMgssT0Y46Et
giXqnZ5LXNEfqSbhPnJWnUcW/4MRRXKSclHK4pkm9f9Kgzi8LLtKGJWPHZrn/X7MA47Dl0veoyel
D79EJvnRDapqqdfW4llb/oXX7nxv2gUatdR4G7IZOdwSUUqH1F6RdZl0t/S4Uagvz+ToDXe6jw6s
te5NpRk6raRz4AFQgRabYftdoiN9rZ+IgjleTUvoQV99Z3nmP6WUNbxEHDPUsLaDMPxfrak58LY3
L2KzlGPFMWTn0DeXrUDofD9fHgoLrsXaZ5TLZs2cAiG5kWMuMXL0RlRtd3PylbS3Su7UM7OKVJbi
MLwYYEsnZKRLNc64qClRpaVIM/EXvoDiXebFZiEpIWQ/bKOZFFO9ksRepNcwtqLVco0YOO4/8YPx
eEfR9PlM2kW5abnXHLeIDMtH6hVmNme15V7k+y+06oFPWmvdclTMx78kXrQeeeANOWOTYTwBabuy
GE/OSbi6HIo8/y6aEzpLSz9Q8MOPytBqR6PWtbS0ape5ZqPDSfBpiCJ6+j9VSH1E3FAyirBkKiua
Z9+IJoikSlHId1B+uD19wD8DX39AxVyZ3bEga59nqcB0ijdAtrxdSoW/SYWh6GXokS23VMb2GHBm
sPBbjkgwbxM+HpSQem/P+UrijqJIrfmTWP0ytP61jvdqUVHBWhzW/U/uf1gbQ9agacaeneUn64YK
5Ipub/7c6UnZVgQ2mDIfyuiOLzgjM4Fs8GtzowXA9N1Hi7oPVbEFUc0OV5w3qBs7uQWssfRB+Uak
hJgROtXckT0fUlM+mJUiZC4iSsb8RzNvQNGBFABnpT6+cjs5dFRGXnh5Z8jN4gH5RbQN7snTc0MS
nVwd8NkaGFnubdJhHBAuMThKXOibkVWo7PNUWKJMvVovWofJRfzFtYjvU98YeAMg0twY2IsrKpu+
xSuWHghDwvjRXTnvV1wbiW2nU7dS3DY+Da9GBxWznpwexzYIRdQQUVlO6jzp6Dt7waVhm4bGDnOJ
5r05D/fsIGwGWBTeiNFCoe4AIJxTsNtMROF5n2GGgEx1qgp+dUvJLIxgCMuivEQZBitdOsXiI9Cp
TqOuCIrBKa2Z+ZsTJM/Uhgnt/wdkMtFHzoHhmelhf+f/1PUh8e33azNZ+WlDE37P1iXf7n9Pmh4b
1hUUuTI03ld7id7eAik+eWEJrk3cZLQ+IylWmy/3oMRfh5ZtBrc9diPEybpZkGltjjkdfJvLd5ib
o0emoHfvSGn46X3A0ZoP5TvMFpEcRwAr2MIx72NysF14qVnQyKHjOxhnDmN3+u96cboaKdH6JDZ1
HxQXxmksUdu/53FlRs6SzTuG+jsqgvZxinp/RdtawVoc85O28gT1TgW293thk7LgKUgtEzH/hwBy
vb2MKupkGF+Rjk6DI0tcA8z+4zifsifihjdDGb6dl6uZRYEbGgQ/6d47yQfiDL6Xd5tOpZ68ZRSz
e7KU0ZrHcltTWFrP0Y2Uqty4+0jhlw6rwYV+pHatq/EbUMEdETwn3dN7bdA2l3Cc+XCIhLlNTQlg
8AltlClwaPUsY1iWcdUywVAlYKPXDWWDCD2QCEnyyGEpmYNdobbS8mgcAGCsgOa+qOlxeNsheRFK
wmaalR8StffnzHxJr+S34RzX2iyQM1qz2/etyHIZkHzBWFla6iOYGxnq0mXZ+4xxe90D7UBIdwg7
2ZtNgrQVJO84dbEVkwl+CdlTvELMOMYh+eVKnlbxQC/hIMvyV6dUKQgHgcO0ZOuujaPlHqIrmg7I
K6CgE3VXkVR5Kk3eQSSLu3My0QOw8tsSbaZEm4Bjy+8DLUJLeQtO9TipxRDRZdK3slayGW8+tmVM
7UJcYHWXWJX1r+4HLdmZu8KK6mTRpK/AoKYfmSbvBTrwEyK0Pw1CU44bamAFMealFNTHsvSnMdPQ
RSfoAwjEMFV8rItzNgOsRtctRUFs4mzLA/tqzgpPIc3U2nyiqSVsK+dv9dRCuDMqpBXxDFNMShK4
1q1eK7AcHADmBC27Y0r38NlpI6wrDxQ1PrL7uABUIPg29YAdBxQsEi6QBnEC7t4CDc4xULUi1MFb
GE/9xcpl05icsjgzZgc9++dNm/ePhclntVRoLKSLL5tM/3vFVf8nBEBMLU6ya9LCYSpGh9U1F/1Y
/Dazww+Ojjz9ZMGOjWqQ54Cey5hvOyJowxtbotn2N1L3F0dqrPYKBgXMGm4u4OtzIcsB3WOqa58Y
CXU/TicYQ9crBPQWXPXitYGWL7e3iuvzcbhxXinUSBHaB+WE2tMfRQGBHj77rqZZRb88JS0yyCrj
ZbWGA+jksuqjA90r6QewU7ND+Fl2c37T6RAqpk5wy5bri0zGpv0MdkjeDETasEqS9WonKGgJrzQ+
/PbHMMQHIzsDEktP7Azhw4fTcD76hUs8mrK1wYlg/zxo0uGs38dL5C9vJcORsemTn9FUhdszQEIg
rs4NBoEa+rXi+Yeiuz4CtRcJAUGfWqyacPqz5BZc3WNHWt9FMo+jAPZdk7CAPFMwFFKWOnBC9kRO
e4Mbihb+VMMBTW01yfdTCW28/HBsoeFWo6AX0EK18DolB/Kw/pAmXpNX5QP36vw+KAezUZqpxjhA
3/dtLg7r7/g/OgLqNs4AwVIVK34TOwXfOpIXKdKC8PQEkrjbGD1K6p43IjIFAqzPYpZqi6rvEQeN
SIopcigJKV0NND9SpUwfdbbVjzhsOFI1PxjMc6SgQ70vIHSgI3qvvFOHuFgIVXVQvzA/oEVyPtIz
C1egUiNlwQEizJkNNKUmp61ItMC+UNkdu8467hBCVDRXnlUI4hcf5HeE3MswvRi2azujkBLP/56p
jr9HjArM/f3v76mGlI1yO2/KoEMpAAL3n1GE8k1km6Xa51GDe6mSgEm5mXZ617a7wDcyw6b3oWzA
OoJmfF3KtRpW0u5mRBYYMkhjYPbGzos10Ob4RYqmEriuM9w68ie5Oa4c6J6/xb1BLTzMcpbDIQj2
h3aIi/WSpv5ynjplce0876CJLmgy8tW0fHrF/orPAN4zAYuDNB5IaIM1TKxchgwIsgMvupiRBh2T
OThitTw621K8D9icRpUHVpvR58sUmybgGOWe1Eg89pGXOdxeA+9bzJYBvYhOmUw0UZO7x8ooznPQ
moaTj4u+pHBq0Z/gN16Ft02nTIhYX78mh0WeRNuLPqy0t8KHGGwKLzvlbavemSbwk1gLaijTjSr3
zQrbr156PmoL0QMgL1IcRamUsBufPDSLzgiVYgQETO/f0U1N2b9MkZVZ6fW5wxROz6X4ljthx0Cf
d7P74Bq8o67b6a8z6rokA4/fvrpYrENIZ7sbPudKm8yVLMUsuOPy0Rfu66QTx/elCsYc8iRZXFc/
v2YN5c5hQvcBWKvuEYKiiTnlSwocC4CLNHp/boyH+ScWBsQu154PGceK3Gny0ylkQzVwUlQzv3kf
8ZmU6bslow3rLw3cQgVSvJ1JaIQZNGzIDQgMskdAcukQLsLMxn0KUmTT1xiv2SPM5VpgZMPEz+AH
BV+B5ql44mDnCfIYSVyhufGqQUbaI8LgqH/hEGJmQiu/7xOkyVWYmV6vds1C4TsLfUco1dLjvV9V
YgBknEOtpvzq38S6p6UE2TeWAO3kUWy29UvZfaUX3GDJbZhnUxQhgl5D81E7Xxd+zRCZpk638QGI
AXk5JZjheNj0NcIEdODI4tO+qlM1g0BGmR2aAcHJDRs2Ziig7Sknrn/IA+RTRQw6kiM+UYJWbA3l
xA7M8TVCVlcDUnPryBw4CDeuOzccVxmPNyOOUprqu2by+o/G8nPs+RVj/8A2G2AtHJDR6cpPZxC8
viIXVT6XyHesicfECRQO9GH+0fRUrOiteMHNyYYdhrB2UeKUAGnMJ12UBJbeP6oNXg0uMimgra/O
LT7O5svC1tsgUE64EzcD4Q1X/0nQo5eZAYDAnvcRyg96TjKIfzH8utG8izSAWIlFaCA9QTd+oUhx
16xfJe0IQuPapSl1GjjtU8smlRVD8osFXdMio+z8/4QS6joMIgE/8yh1MJ4lKgnFLcggp9oocr6E
Uo41zEWrln8qhGJ2Te5bs1ZpNGltRJEAM5pzZJI5jM8sErkVW8tEe9kzgoC2bJLhWvzWKb132ACf
fVPHjqDT3pOUgUvYW2k3qtbpHLjqPnsl9nKVPQax1eo/56VVuNSf9Ml3UztcYtCGCy8OdiPbVDku
yJzepxQ5fC/3lUCdHA4sXtZMIBpV9ARZMfjQMuswgKJuJ/2TjGUaCZojqpGW2n788Cl/SQN1so2d
OpTz3JyeGmWOLWasEnapP5XLvIghKSjcMcgShaJvwMrItdNSDPA1Q6vtEkokWTm5UzYUaV+f2zt5
GC5Rg6bdtXX3WoyYnWCjwuQqvycqLTz4uVsw3QoZ4ijcB0ciqNTUfiVJXeS5e7NtGpfIxjGGRwRb
dhotpf1OFTNvtZKU15EcR5cwknkYAP1siX6K4QXMfQMeNQXaDcvq2WgBrHsEODz5Lh7zPHaRzQPW
dqn3CTWQn6jd1z9rfTHJXl52SHDqJqK1i1ujt/4Bb49udX1ObL6GClNybl6aJKemj8GSKDjGvlh1
bPAKmv3DJk+1GiyPg1V9dc62vIlu8iYjMat72m/rACJy5EyALvyMw/1ryOlK6TU99nfbEkE2KUB6
BD3x3CYcx+vX33FJwTwzqPJt7D/SUOb8C/LjKFrjqrASciR4gL8uQkB8qTYCw4DGzUd1adIaSSlR
lgkf6cBXDnySv2RPPWq0VsSnKsXpKm/GBAloCglbDxhBHmS6cnHMQjkYbIiXnfM8PxlZdyOcAyum
6foOCP6DaUq9iR6JGVSCExrRHS0yIlVH5hC5jenZYwesP9i5ClSmF+E29ryi+JkNi3bYfL0mbh7k
4v8/90tTSTO3STKnLZTL8Wk3dvvQhHhFdE5rGAM9oAEjRG6b+zpRY+nkG/o4n9DkNb6813eMK8P9
WNFNYeX58hzwDg0F3pdCGrtmCLwiWiCaCnYlbMH4++E6Vk77LwowgMsTFhVZcmHzVtozhD8UUfsb
S0Iu4TR8E+jw2/hc8YPtsiHnz47vCLtAthuGl3ioJwDZj811Hoib+24QxLmE2cs86myKFPA2PdIC
zUdsNrHHUGTjxIjvAzriV2qRbLym/GMLuD33hHXyEjZ8wbfCCHdah8RlY+j4cPmcWQg+plkCbaLT
zsQdwETQVISdYDjJXeHBYhI4hOG+5zNjnT1qI0h2CDEUGX5x4sBFrmHYLVWoR9st1HUYFr2iOaCp
HBvCvzKGey7QkpxKHpfHznJ7BkXUhORopGbyTWrrInfKZ7xzmH/XundJK2ttjQbqlj58CA5v3zJr
687u1OR8kFcI2GnHfcDJS7soF5/dg1+Q/kowqhnxCidvSuYy8RrWyKhxWC0BatqRmhMKb21S9SlA
kZM5tfc5T0foQyfDAndcM0QDyoN7v0SdM0wnNz7sWBMKCqW2V0dnFiMek2DYKL4ufP73Gmkdep2B
U96vt8tcUBKKyEDmX6jgNUK/8qO56y4T+AG06JTWmSs6LspdIKfyEhNh3yQ7U7geE71IoQT7nx4B
14xeEskqQS3AfRWBF7tyF6Uh5Av9BkNBE/m05PEQmbD3Xc2NiTuJIrSrNpvfSio7meeKED8rbIaZ
5m3dAgW+U3Uc343xdmVNm9bG2yTuM15e6TI1AdAwBKu6OTuCR/RHEd0BdoWOZtU+0eS6x7BqwEM3
cvpD8lXgs+D2Q6tXhYicv2lwpUFvV4mf7kUfilaCs5g4SKGGS6rVglHHMKv6LQNu3HQJPfeIAKgT
hvVH4D0JJ/RTxS9L62P3osv8WLp4qqoyMwGVXkntVMho5p6VGxYyK/OUDkuY7lNYhwui8kslcCN4
VBM+wirbayITlaYjrb9weaCKRpK0Iz6uKkaI+3AQeOU54mdGi5CJfOOavXPei2pZ08av56nKVBio
YAP7M8FuC+TErXPRwHE2ASQKgyotX+qR+6TRHPRo3humiOMlcpf2q6X+4NePRCAVTY2QGvcT0Q/5
vz9heDw8wY7N4ZUMKevO4ZWQvVLvEMqpgQJMM0KlI0XDbEbna1h/CGGMwM0wL+3sIGjqakktWlG6
RQVsAwZFZsaacvRDHRhReD0+HKKqSTPhFDIN8rUiEm4gwW6EOEW9HT5ysqo9jNPvhvpM73mJcd82
m0S12zX5ReX1X2d3zjs9Ol3oKY5FcuVymg/7tTgfteozoB2TgiAfNNjoWAYBsJuPqdJkh23mzpRn
BP0aZ69bAcO9qlBOfgPzkhNvCj4g2LcTVRNkd0VNLHjVU4aLuOj8rgi9k8gYz5NsZaxRkZbbEmM/
K4WUZcgHmBVd+0oskpqeBEmS+XPtI0Unoq1upxaChD+A/icyd1RiobuM4BpOc/oxpqfLIoPocpxr
wrmosiBH3pbbyGWoj3ywT6NXUpUS7Y0FQuK/FMu9/BO0tiGeKROla74rqdTrbCC0khHy9b8G5UT3
c336YKUrTjocU/OdUzx7tXdIgCZaRnknYc3AmLPDZW4FRGErhjeejQdxXdkLZCuyazrEOk8eaw7K
9ig/L78puyzAxutnsbdJmE+AG0+qxTu3dkNxZkzlUZf2oBJ7RtFb5ZUwITGBkNXfmuPJNCWQEF/h
FBUBhPtOGyniwS5N9I/T7DYhqNI0nSJTGj8oLFQIWViipGY02pLBhpmeX3TK8VmDe15CbfrP0Ni4
tmxEyLrEzOt5wC6Kh7DmZPHw3yol8jiWi4Gei8B3b3VetrdiUS5XA/gcG80WKh3l7YAy6DcQn5O5
2YuKktSYtISVQJCoL8POsD77NELx5QWoN5XzOG7bUGGoJx94OQHUPqhP3/ChxGP3cwUjP6/Mgoxe
xRS8dpsXWDO8Ln/tBY+J07de+niVwXE/j35GLuZUHeFVc/WirHEILpY7KFmsOpN2XLqWpZ7ejADS
oJQZALx0fS2u78kFA6OWuYOPqOi5nFIw6Y8iwczmA0neA9aT0REeIkKu4w2jCdY932O6C9418MYQ
RQOE/h+xdKgxEzwajXQ6q1naMuqygpbSmLjAbp366vC7xewmoUdxTNJAL4PBzME7VehjMFYTd5UP
BowW7RdusqrnchB0JsvcDJ3Kg+p92uu4OQaoymx/mSqNEnJmkdKtzGLJy/2q6PyYOVR4gdmyDAB4
aTduqMdaEhaHHGpYqO8j5V4IMXQWBy0fC09qQIFvzGMecs4EhMOBQuZ9jnCTlWlnR5O3IPkloGx1
ujEL7jMjkrtofwI9ryOuLkYW0rPDSB6j18qAmAt5hZIpNlX255EgvICHqZD3MOkTxBh3zoJtkED1
f9rNS5Vbv9vQHLRL2adAltjCFv1g1E4E8iyCAQg9lk4yjZnBqohvXU1I5tcKkE5z4A+KmE2VwmHj
3oIpMD4Y5nmdyiPUwVCbkTf9mdgTHD5H1/YTmxjerU8vB7pqS7CDgW0drMFGuC6/j4bvu0DLGZuE
ZC+4YBPyuSpCr6Vcy7dSEWnlHwgux8t2OPUnVYB6YFqTwOduPMCNSYXdnTzm1QQNC3/6yl7IDP8K
TvJx+X9+Wlpnc1qtzvBlUjdPyHkGiu650pmdnDYYK7ado3qiuMues8UXvGF6wjfGAJi+/m8qUTFs
6O3HTS9v54vhbD7pobam+gHe6xrGZuWHbMly8aHnVAnBHsSJL/U92+Zb+aG4pNCJ56ThsO+pbYKQ
LZmZSIYmgzaB02GKaz2g1wFuuVVJ70GZGD9fC81OnmNvnNuMxxnRIJCdllFQZlwagmyTOLcWW2LT
I5/zR5iDpslZIFoXNf6oVwmHcCnO+tQpTk5U247b8vylxuSx85TQgN/ZoexIZBps7l50eY6iCsYs
hdZ9sxVu/KctlKWSy5xWg/8+HqwliTsuoOBIwvaUBcKiNj3LhKGf2Hl0UUtMZb+6RC6lLmc90l72
CCuVFoBgzRSjdfjz4Wc7dh4sPEzV4vfVQJn52TTEjLbuSpuh9G5iB7qr9pftAplhkxitSyt2JmJJ
q6MruF0kvDmgZpRpOPosurATfXejLYyf854xx5wWSAvmXnjC1YEnT3sMFYy1bH3BIzlv4/4qKAQe
0Np27ctM7WXc7oEw4TDbZL1rNuqar8LVjss4QyGV18mEUcbHFBTrm+1M616lkBgzJosyFg6KWtWA
AJXJW+Wi8BdDfSQQyWkWH+aCY07hUIiHg53ubWFEUFSGI64q4IP+6cSdUfqKstbAE0q1dIgJAxZ6
T3fkRHXrt0MBoUm738IzLEr80RH2L/BYwybD41AFGSqyku0SKsLQDaK7b85nl5wa1eec+yL78m8C
GCER+x6TpZQfC8Yns9Kjf6awm7WH+jpyT6q4R23WVAUJQEF9DMkh+oX2PkKk/3MftT/+qhbjqmV5
ncXsIlHXJymQDl3B/l8dS0+BATsq5epfZFq5wwnVjj21sRnexHTVS/6o+eUrNdRa8G/nzoUfOhw5
sDMT4N9ITfO3M33rd8ZnngxMr00VFE5S7EBigVMvHmxrPmJ2W+8OvHrgITcsk/O0Yae5G0nwMDj5
237gu1Vci/GaKzWbiR3Gg6K2deQzq0XEXc6WSIf1rGDa8x4MFtAMQOdZl2cixWjmnld+cmXNTp1+
lHmlBtILzN580yLBlenAUPeQRRqSEQ7Oxw0UNcIFf/gXVY39+sY/EYTO3rtIlg28JwozrrpQWKjO
nBCCkg/6eJvU5QyYhdz8bdLd2Ffk6jVYFnLweYux4Qvg84cYT81KhuymBerQRtKfDR1Wy+MjCtru
DkUKfRdkAFWKANtj5ClAqJm9Yfiu//NG6fThsyIhV6+mIKTYDvF9Fb9CaS2HkalehjfRkT+TPWs3
wNJllNUBRnAfyrtlq7PS2mn2marvzeAs9ydIlaSh4ri2qYG3zOMKsAb8gb9XWYj+VsvCnSBhfSK6
jIdUONMGxBNvBkPePHrmSGmiC/tfWlYEo11s+beN6bwJ9zCChjx+ulJNFXS2OsN3IJYkQhUjVygs
XZJ4mBeSX6fVkl6o7qhk3wuNge8LHhfxsPm9o+TIujn7+cLHXT3Cty9VjsyVp8ad35cUC2+VgeHl
TfRp+Tk6V5kHXZuJrGpqSUemmN7yHvFp+9bkSqGpM5XZ3krAVCsXW4mruKNna/mhPsP1Wb3Cu5LO
vjqRAgJapsF8xRLhP+ax/NM5cPnULbOntyVCiUcBicrHk7bVvgDV1smPlovNuomAdrYUo2khxu98
m+vHiV7puPoDyE/Oh79ykAUh2f86zQaWQ5CPfeSBZMQRHIAyEWbjDCydfZVKH6ozRoJOYUzsPhUL
yewDgyzOc4QO7d3RFtBs7H2nVSgVrc8Z3kMVEOTSTW9gXQzIu3XwwvQTLHuNoeF2E/ku42LTf6b7
AzsT11iWrHoB5VS0dm4/3BIMdovr6oVx2BwFa7vcIdPPwteX8wbaMiA1ZO48hWRldS3by5wTh+xW
i4XUyEG8m9l0KJHCfzh47Te9NEy5ilsJPVFlF0WhzDT+v3tImd0RwWa1WAbIjB0cKtcX9UhGkHP8
GRbJfhUulBIKeLajH8S3H1iCR+FQtLFenr1ppPOQrjsVA56pm8DG+PaQ4UseayNeqGuA7Pa8j4Hi
/+9C0ObSwX3aFI7iTCcUpxQ/Xk1bY9dyoxlY/CSkgXRaYIkL7cAkUwLTw/2+9UxP6ZcyiddrUzTD
5oMdCb5rYThF27HA0TBq6l3fXyR6mAki0iPytDiyK8gq73hZm/WUlTyiMj2k+d25hsWY9Rdr+gkm
Gvmb6L9OkGG8P+gUhTF7HwUv3QB+PmetWZSPIOezJ6i7KV6k1gt/Xd1nLaHkKJfTV+ts0k0ouQ8G
hotUoOAonabgIuoVslklsJKvIHqkMiL/hA/58cdSC6PXrGjbbB7lpkBwYjFMmp3tPapUN2B+y+MB
DayIn6dBr69xvfaxsNbhERUF7JQ/ioPy5jp+a5kIMO4TXbNByFmcyR8B7nfWfBPdiZT8xWlBgckW
E1LZ3yFV3YmcSZ6r1SU0ZfsqZotScU8CwiRaHh7OOyDQs3qCoUDctsO4yYShoKN5VrR7cXCeqSmT
WV4mM/xOz4HJh4LAX1mNTX5gCIjnoZIXm3IGozFLUNnu/goyDogwU4bNJo5xRu6vaa/SM3VI0ZwC
fxQ20YeDx8l5Hmh/lpSIDHX4p032+GPqtasmtV7qUj8Zz+an+OPIQy2OhQMVB9LCotDIR/SzqT5M
orUAauNtaV5bqTuTZi33Lr8CGKe7MJybFPrqghxnw2JvGmL0JTyYPabE0KKZJJsKv7d5YNnu5LF2
grQ1Lfxzl4FNNqnTTMkrveGIIQfV+Kg03sWVDjQ1QyuvU5NwDDEmPrFkptKjDHEXJ/9urVk42ufh
+cUcVj+7PwsFeJCPmMt7buFuoWWUmJ42bCZ0BqrBg25SzuEzenopcyq7wutRSwau75h0M0FVuDt9
rPA9Gs10QuKYRnAnoqQxhSNYIxNrlXy2Ex2/aKhxEPGE2g9q7vIHyDHoZij8FHVVrfJU+k989o3v
RsaEkDfGyfDq+/tE7So6h0x8z8+H7BA+sCceRTn9fElvt3Ow1oY60jEVvkkViZeWSb+QbwnR1Vfz
6ZviM+AD4AGlnqd+maiI0N2XIoPvu3oUF/GKyPv5Qulf4j0cdYDboLHgXxabXH7NjzqRoWNmqxLB
J7238kwe+H7sNvCD6czse8OPFcAzLUMu0EHEBhDBpWxlGruCl241k0d1gmDaaOIB8jOEmF6LQ5ak
lUSSa8M53KtCqUYyhRp1SALxUSkd0UJ8LE1L2EmmVBndZPHgZj8aJaI9BZK+lCPnn3Xa/aBTDkYB
NbBC3Pl/CYZE4mMRRS8tQirXd2P+6Pf5xyNyrgyUQEBWP2ZgUAq9AN1wPBee4YNbJEtFR8GvKr8Y
WFcp+zkSXp7aHt8I6Hz0IHLcGOA4BPEuAY8f/BeqyHJHglmWZvibRnE5mO7VY1wlvUD1rI4+n1j6
QL16DyjSkFON2SXoPUtd7Y8qHuzif7h9kFe0Rlhj5Zx7Ggvc3Js67rp6IXh1dzZK506vGgL4Yw59
ksCdGPmcW2XiHZPuLG1QO6LNE1CBqWvHkMvQQFc+MPDxFUeqa19PltRB8k+NfXAtDvg1gMzin3i4
r8qaC8398I+uFwCg0Ot2iwfb8g0PPd2XmUZMzruymX1yUl6ZFXhh+/kBtdjTPmDDHkCxTi+DzSzq
NvTFItNM8ljhae7uuGh354VGSHD4UiOU5ikQttPFsm6gMrBa5fdt2j9LcoFWDA/pAIJE/a0iMyUd
Jq6EkX7ZgCmh9y5ytwrFii7YY19+WGQLKtFCWlVNIhc5p0o1VnJdJFfxmX8gEJY9tanwewbGwBll
J/iX9qDaf+mAN6aToelhcHFho36HUHx0gbjZlVYNZoqmyaosJJD/U0wb4RIFQX/tGWagRXeOSmtN
BOxiI2+xjLNHosLl4xkEUUiNXk1JpR0qmJjDeO7XttlQ2jB+GOHNbVJPgWhgf4fMs9MZp34o8dFR
MamQoDVcAe6HAl++q4tAYZ13BGx1m+DZAQX5WgqoIzesCkYUN4XS3J+qtBtro9SGwlo+/rS8lBcX
wqzR7ixRd0QfSQtTOiTaQKLBGrRVBM7CxUh10zqXaGwEc329R5EPjCZoTHTM+ai7QJazmpQAFavc
U5z+JERPGcYKetumwfzu/mR4bCjAkjir+APHrEhDNRpKi4vriU51pOcgkSNang8Xl6edu3XjdumF
BfzZd2UosgF/2A4H04holmzWW+rr2nJT/9P+PJODeyRfvxkuFOxI5aEjqtGhavyBbvUgA3/FEgTS
11leDjgkGu2nAVTqQ8IhhbE6Uv7NClLVKjhugmT7YZ83HQ1iIDpcdnVhUDz9wRegsmTxT/BfWMVC
aRby6mBEhLfXyOtZj8WfsLZkRIXnmr4zf4Ia9mTLd2NTo7K6QjJLho5dl+vnV7IC4pjXEVT8hpxE
gNxY/JtRNvLB2aNjHmaBpuBH3+zmGwGm/F+EvUYWGSoW9i1l5f0LtVwoK9YZuwwWVhvg2Ix8K6WO
i9Tb2jb2wmVhYYXKHf8Hap8o5ZN6+fQQjZ1WYIUIrRdm8387J6Xd55iw5zOvSXrALO7714RnsDp3
/GuGQexgHp1WXo0pYUnxkVpHOPQm0Yr8kpbAK9P6Q30LNF57klGLz+pGoCyort3Wy4ctAYR/xWFU
v1BNssoFpOVxz9yZaOKEHE+w3285dO4gfN9hw20obXNWQ/dcaamWRkRQssoeLWueFtU/k+RxxQjg
MAng6+eBVm5NpmlHAklgPNwmbBGAaAlWCF2Xz9NXIJYkBtioEAloUXGeKCBp9nwL9NpdBbcC4AVV
iemZtTEMXbFpZavqtuGwmV9aCOjlxlKj9wkbBK7H+jTpjEGmiaLhavYR8j59T/ZHFIB/xJf4XRNN
VOOPXVPscJTfTIy4zUUlLX6cjSw4Dqt0u3mq6oRiw/bSUcZmqrh5jE5NO6m6qjQRXr6NWbQXrhSk
DtlO7bk+E48V9jUHFZMJxFKHwkJsssGUTxivvKBYjV/Fe1+iVWwVETb3wVAcSoTqBv9m009Rky3J
N0d3oNYxmumti85Pa481VCPZyT64y5qpJu1a9s+oIWP2OeyQ0PX8CYhjUe8rxCBZZixxZGSaaGwu
6r7I6JxRrqTW4WrkYPD+TK3fBpu3alzog0tuu7qYNcgeRcrlUBiA3THtkdl6xtm672vv0C+Zw+Fi
JPZQ3+ABTkn+5KZUGHPgEuivdY7/gHTAmLwurqUhX6ZOhVetkxgLy4Q4AahvMHB3+4F9aigSh1c4
HBDJKrl79G3LdgxIVhHuAqS9zAQ+nk3tq7lz3sHyNysEoQjbq+xREhxTXXhugOHYT3ZLaoP2k3DV
BgKpp7gWIY0XJnlV2bjnNaEkXEthoc0cVikwB85yPHZHwGhl9Jb9uVx71jc1OIwnvl6BmlfYLbgN
xAcd4XuVWd8DvB0RbSKil7Tb5cgxBDFzbGxpCpm+mq3lmO2r+V6xn7K5ASQOEs42E0wBCo9t9f73
WZWrfNwTzxG9MQR4TSCmYDG6PjOgJGBsu/lAEQ2Ir6jZqILZka79X1QkNsfFc5rxV3FgzuwJ7MGM
mNgZYyPNCliy3o3rkKtSYDjcy7HB+e9hCahdJLz+eQ1cdBj9XyNRbc9nQmSbB0dCvqgchPuwDmyS
QboH/r2CJw6aoEg8GWbhyAG2bxmDDxBkknIPFcbaZXwbeapoLJOqUpFb4HAPnHv9VitqJ15gaGyp
7E/IYEWgZWTy2o/PwLEfIdbtZQQMu5c7VJEFDlWC07FxIQOQ3I1XHEjGoHpFGmshY4oFdf8RKPvv
LxK5SokZvXuJ6jGRZTp0Lu6pttiO0vjI7RtRi1ATTmIGK9Dm1Lr8o0Bu4DSXNuOXbMYf0E1snHgV
erdNsF34UHsb67jSiUN+BWNHlZgi94I+bAXhB4s8D/qr1sWsv2ofJgkKW4CS9TzEI7hIUZTTMnXD
iDI2b9Z+Ko9c7odvjoY5NOhUDiDrPfm991JumoSjHIN4UFVaFe94Lo5kZdfmOvErTdrdNjfvVEgz
ORAwgoOPvqHdCAY9AFh09Rt+2XaYYR+ALy8kvfX6tlkQ5WAXKC6+RrPgOMOF+BqEKCZ7AZsDhBOV
El5nh4hxbsl7uAK6dnE0ZNHT6/Ro/BhuOKNkpCmK8M4X1hAksLJDcGOeFVFFTZL5VbqnW3R4ij2f
ziSk5461ovZIsO/eXPvzxdXr/8s1yrewxo/91z3JSbW31BWjK5oymNlaNgnDPwr3J8/7If3rSNdH
/QWbXxf15pch8nwCACjpPQSmOX0vZDewIRXXIYR6b/hQCzbPJLbu7Db7ggOuB40vlcLi3+rqlmnO
ps2R+3h0Rcl/X8znMX2xyCKRA6wFgW8iHkUE+yO5ZmydbUphqy1eWCKXvHW17zsebOorPkwm4k1B
vi1YTtzoIn3X89LTW1cbd4SqA4T3H/W8DTNH9brCsNyuAAY2CQWyfbZZqT2Fgewv8mI6TVEA1Vda
U2ZinOvod47ivOTUxoRmIVSs/S2G35P07j0s6lU4Wa4X3IKeQSuOEVNdJ8OrVHVpW1CvlyM2qyi2
WqZJM8rEpgC+jre6HwT+zvUkWaNrWVI0jKxDcmsvg1/N7IdqxyP2j+Y7uJjS31tZzqRYeg5csDzA
YfPnpwcqnjX9SByr3MmSlhR4WfRzJo0/XWGACOtFMkrBLDudr6mnjxAGFs+Mb4zts5iNvaDQP4dd
wkzcHT8AnA1PCxAcKTkTfqoCKxUq1IcAy9XEgmX+4+j5hV+vzKK6kyyveTwu50a6crpGDuIDPa4q
VeCYn0OKSx0u4n/muC8xvBBxJrFB+0UZF3zjmqX4Vukn6NoLgeBZHuBKwJQo6CapKNSIGiwfzgdx
Vzyua2l9JwGdfwIrLR3q3d/ccEZzsZQ6qvCL+tN991bfycN6KF6KtZJGDiBGjLjMWR47YTp4chX0
B5rrYFyRK5cbiVGgbDTEGuHQGR3bCmMJBBbzyi2SFClTSmYCxlV0GaeiT42xMrs/x1CW1d/HSGcb
tzrP98qZSi9lvPfhUqD+qmXVPx8tb6TbkL1bPH2fnRE0SUFYYXtDYCfFKdIkBI0kM8u5jo7ovt6A
75Idik+e2J9/IYRnF9uJaOyVhQTqq1ATlJct6++pg9/aUwAtZiLcAIRnRwvFNCRvluXWEkGLbhHV
lh7DosEgoksIoclRZiWo8G+EFCEKwZCsM8JOmaHNzdkRxn7OrSrejcgxmVkFPP17YM2l8iqFQQOM
PRkmgN9rFVm3q+ypYYj+483DQwdVepU0CaYmUSvIrZaDVNZhZzIeSkE9CuJTUi4Ue8hlLmCIYD81
4c1nakRHEnfuFObaXbdPvvdWgIohZfBktctczqt03yrdkL22aJSheQMpMTu7QD3GsXj36v+fe+t7
ID9s9+mqHPIfZFgdNRcyCbOUxGERy2jTokCcP09Ut0jLpW7KH4I7VXZqvWGDfNgNQg9mroHJ6qzd
es02JoVk7ILm/db+gyOOkuV2dfEt0S0HOKnoH2s1T+NNBob3AjUDd6yRXJFmcqFoPsHJXdIw+Bnu
s4bCk9IRhm/6woPSYn/96tqkM69eQjqZM83wamS9NbnGVz8RBvm24/Li8lyfhtdGRcohlWv7Pmyw
dZ2F4aIG7yFyJlXAN5UUHwBJmeBHj93HaaXzz39zYAx4GpyCDdIQBn4RFYNSShH9ZgE1nBcT13qN
QQUkf4Up/GTFBroqL7QTG6yp/uzDf+Qeggw0HXsnV/C8R1JWObIHpazZJJ9wGJlWvc/v8gYtw2Qp
Df+Tb1GLT5dt1huJxLK1rYPY1GXSaxBmrQOcJvAeam1ywsNYDbLdRAp2/mzPdR7e6AIsETKbJfUp
grJANfOmQOna03cmAadAY+vWqfF0vK+VjpwCG7rTVvkTfQh9Z44PLoO81RdH3NMwUo/Fjw+k9KA/
WXjN5EovxzIx657zdWuO322YIfV+WvzrAVFgL31yhrtGvn9gMMYTwco586UHKHP6Ox2pNLy3wiNL
2EnZzke3Yn+s5/cdjue+3EtH7vdG04Uw1o7QYmzk5yxle6zZhTeodw/H5OJ/XEOi7TnyMDoBBHSi
FecTyPDF7Av5c1aPZBjyCuYW6uYX5dzvk9zQ3Mjv7apLJPwPJ6zvh4lE/DpHsWVQ/yAqa0+zLqVY
sUaeHoA3Hqpap8avmOfq/yRw6Np/pQQmXyCMamno4sv1WRRlPn5vBtUE3HQY4mZpAIk31tFP7atu
fh1OvjZLXK8ScCmYFAKc6EUeMhG3OD5+6tVV55Ua54IqJsC0sBMZenHr5/4MuWNTvmnxWOcK9Jln
juTEWRjwR/p5q5ejyixfPBwSxv0bjvP+BexY4CuM578TnDvHn/fyvNa6zCbBU5ymN85D+4F5DKQF
BslZ62rzeIaftisHnxLYWLxjbUTJ+EmL0oYD4HUzZujjk//qWNpAW8vMruIdeF+fW1JygsB4D5+I
5mX2GlmP5UCcwqxcgLW5lhwIcHcTeYIbc9QjGHBGy0DzLwfJWAYhpSiaI8oms4rLgn5IYXxMEl9K
O2+MFY2UfDAQ88rW1rc9HBoIqlY2sktkGnvX9Hlwd5xVltsPP6dNJFZ9w82BALJ7UWSkB1UUmuco
Py3MbuKBMTNSXv9dyp1A3UpI5dHKFZtPgemsWASWQWBhdXPljS7/NXLP6ejsSxuijYXABc8oDS3T
yYEGquWPTHXEetKGRL4Z/93Jchq2LpjRwNfGAWAbBuqXT+23wO60+CwhhxkyvBqqJ8sXZ64HJnHJ
uGcjTSxZynH+VGVrbqgFArR+8dJPXUBd/p/8+sBX2D3+Pyzbuw8wE/fNxp3NgzE2bg5l9SQa8Bea
gLQ484j/eZv9slsM8DKNUaRkxTRXIyWQrCRXVg5DkMaTff81yu4jiD9mpYHNQM1W7LG/VH04LgxF
7c/B0EpS3BheCT8kx5GheAeE0LaVx8MeMK9PFXvMlKW6zaWJ/gF5voq2sKSSVbvumjo/cg28ab3M
cNMn+yj701vfhgMy6nFf0LFzshSb2nKeWh8VCc0jAK4NFj638dbwEfpkHd4OPjyRDQZZIhh49ht9
l3W8pYbaTVfidZzzn6lGk04e10YwZeRzyqM28qKGj5od3dFvi6mIvllDysfZ3v2Icq59F5wGja12
s+btstD76YFbRiBrCF4HVmCWgmni9M+Qj8UqsZmYwukSW7HonBNYPGV9vYIo6FR8zC4xTaZwZcb1
Ql3kUyvlelm6t4pHKoH77nAib+JaMzUcySfVqs+ydTQGdImN4dUHjPr0ZHUZ6MWs0vEBsW+vyXh4
ZWy7B9D88Ztbbl2qFBigqRvIJbhTPrysTpfJACJVcMXGYcoHd1b3LvotqizrMDLRkfKtoU7sTs3m
U9KR40ByEneiJJGDMQfJTiWp2nRots68l9pSV8FHfnxDabyuXdDtk7vQGdjyVt1rBgVGQjTaf65v
QlJLrBfvun2Th/4NfprO8hCRtMKC5QQY3s2+3PHCkf64PM56lNS3Xv1+zju0FZF4n6RJPbgOobKS
l495fGYuxnHMkTypZbY0+GAwMarQqc7Nzbktv9qF0YOIPWD2XjZ25X/A5+RwI4E5SLHzkJ6+KHfr
zjX/aHbTbxtQ7gcxfR+wLSJbPM/tv6au4jEsmVTFMux+0yE1VeTrTu0h9T7wYyifAVJNNGhz+ZUF
ku6gC+qbuVBMKMXSoq1HKmSgytwrs1KcoCU6mfJ/Az5apf+Rq0S0Aqu5bmQejla2nF+eVhRL9ubo
EcdPs6J+W8oA/Vq5ImV6ioNlQVe9h5la4tISZpw1M6xoWQmXpyhpMqFwHnXB0cjbk8kRmgODzW1T
5A2Iy1wIWPvLmd48dDe4wqCF9MX0JyHHpUx3yG/wvUF8cNkMpt81M0j39Dohnrhk0XcrxLAlH6EO
oRAi3uKvaM57Tn1kfeJaqCEfUAu8POH4T7ZnzF3zf6QVTMexggyjiTIIETO04WbZlKIHK35M1ZzM
1FC+Qb6hiiN1PUq54Hxvw9uwFgU9tyPTZCCCiRr9i99eFfqqEMglTa5IZo4/VCvC1ucP/6AFaXkO
CeKwdmRCOqs787TaD5AfyLyPztYEvVbxURSVQg8hOp3rIl6iVWIwZGdF2I2SV1+UbLV+n0UsCQQy
xXccPRI7dv873LqoUB54GrZqwRxVc1RvEFsMt47N9r56vMew1GvOzlP27yD6vxgk8+kE4/SOYMZ5
nd5ZCBexdKW1funfcWGfQ9V3dqBjQwMON/3mmMAchqH42CJ2ooLK4WIJYZjB8I0yYRCrDfFs/Y9Y
VOkmUXdDjmRGPojTTuP7xe4WMDWCXZSAFo6wA6ryqGRbAMemJyAkl/09TfylnidUuKkCgirrbcO1
KncYOQtm+0o7yfdumXsYXG5gsqV8X1e1jkcB6H5G9oh9qr2fiNiDULZ9HKRVrq2YFRT2Wcj2RZpV
CBr6daTub0gDR7XoEC/UCdFhTWV21kLUTsIcblJpMNovzLGAX6l0S5ag0jpkIXKOHxKaCHtXn/Qj
qOOOZ2PipchN1rxOambHp8/rrn5soIDaXiVb7Mv9jDb0J0rRF/M5xQtiMtTvuYsF12pVUyQaFc19
88Y/jri/12V4k6kQ8HDqnZvisJElTSzNAdoBVvoAtPj/7HFz0Gmvk3gP5M22CxZ7wk5o0QUoxpLR
c1h+x8wZ+bRpCU9NhKPPhy3W5GaioIsP0euOZHYn7FxXOGhGRCKObl/RoDzlTN4G+9GJ0e21w3Wp
hSOswKmshMIGC8M2oZLfntoIWPvPxwL2z0k2JPyYMn/l2+inzCDgSZ0ZQDqbc9Mfz3LfUsEdL1FB
ObN4mTCAluHmIGXWUTdp0jNkxDlTzVVzoJzCxd81R+aHO1WBE3W0Z9zKSJxFTJKd1qAK2ekWCE5F
sGiVK9oG3qh7uhy5Y5hP3nLfzeXNt//hcevnUNs1SncXERI++ejqCnLlhaZK62A7NVadTm0wMfnc
me8m3Gj/2/wUB21GF3ntrTtjaavC2BCJkruwNQnHbOfUb2vT+24zixWCzpB5lwZmgyG6h3oLa5RK
Md1n5kd5tFk8kf324bMeL3S9yjWTDcv5lBqWkxqT+ScN6ZjwDtHUHuvjVVcaLfHczeFpzc9GC9Kd
22lQlduDmEt07WEXMypkUic3/akHDffFbuR6JptcADsacAdDBph/33uDCGMnOn/ylfdLdzXWwncO
LupL9voKpHQB5UbZxl04HQrT34klBHwlwm5YTaoXD350N/Agd9HYkhX4zOvbRioKkIuyhtzpp/lx
OI8SCoRBpn2XDRyg0VpEO7STm5czeBW7N8ACBkGLbomNXbgASHB3Ti45bdoiwT+acJTWlraYvPBH
EjEHBmvONs/Ut9B4c+TWqCN6A059fVoGgxq7RRgUSQynIBVLcprxKM3MFRgaAY086JB06JgB+2hi
Ywsc4cpIYYEzR6xDXJR73hIvKNaR7S5ESHXcF6XLDdRJdoL/ZT4C6B1gjUk9eNWHoFgGO/QXN1Gz
I0dkRXNJ5heE0Jjh15nP9p090XjbSZExbFPzIDeFcDC/bR2JC6D8dzWJooe5xriERKI9cyxplyYV
fiw/1q4xJfunzULm29UnCskMmQrDGwVPX093PnB/rkZDJEKdV496St4krYVk4DyLxmrS4CqNJxAD
9m3M5yajGy9tdXmII9gtlaXdVITny8Sq6kECm76ln7ouMgGf0QKbD+D0GSJfE3iRmXCkqYOtbcjJ
2ZQ3agLY8/NKojam08lJi5kPu5KJiXqFrdYkWaFBklbmmSFHLcL0Yr7eAKChuzuAAeJ9NeL0Q5aK
VADsYoOVCt7xyXy1udFWo31RGKQSqnUkmvjLMVsFLdmMciux0Hnge8cd/2MnHL2s+hJ4eDfl/N8c
KcQvehuL+yAvtFDJ05dJVUD+DOJuGhmAuHRo8MjGr3/gJMBwN8+ochEhfi3yMED0rrKgLttKCstQ
VLAiZY26NCai+EnzVp+FxvPboeuihgitJPgZGTReaUs9w6g6Szixmmtx07kOyjh1RRSLAFaFUhAk
82T7GnMTY76/UQO2OvcfLTEQwmxDc8+SHSIRRsCAJjh0Yqbbxhry0S4vKaYXh894Tv+3i7ZWGrFO
k58FvMzBZxZoWPklJxPzjWMleeqmjCfTfjKztqO1+OdRtpHoD1Cg8oRzq6qexObUyPdOuT8ENLuP
jWdmmCOu/BOvv1IIlMhTQ6jg45r+zRYCAme4g/WD/iXbWkVwaJlsLJ6e0dXv7QmwoJRGju93oEjo
8ViqFQ+5yv0jwRafflEVo9SC7bmBXuXn3McydI+q44XjbCKGkR1BUbGmL/e96TMbWHmfev+857C4
oT4bzW6xSjQBgEN18NYEu9a4Oe+bt+cfGEw4I69gqDN6BFQkHl46nfV3jHzdb26ojD4dci9riEpw
/vTIkZGFygru1HGM17jBW771H8DWWlJ4Hr5K4y3q5aRZfVdOu8hZB06yMNuwQaTgbI0TrU24mOAF
GYsssZ+gpSMToMXdsmgvSKb1w2qmjhssAQ1OHdsxIHMcio07y0JWnkAC6uJhDuEN01QqhgG3Am9c
DFZ9OvcB3XGxPKRRmOONJuFlonylfWfs+U0EB5mNgZGtbQTRL9YGrrzmKn1u7Ss1+3g53gwWGS7s
ztyzgNkYWIBzJsQ7S9v/hUOyvd01eeLkYpV51sqDJRM8UH7B1uI2xnNWZ+b5KYEtVNmoAFZYV0E2
oWK63D2PGS6Ig0DrCusdUQZI4TZMWFlgrJRZUL+dWBBcxxopd7Af+bowkV++UnW2XYRWBt3OUZDY
jSlKDn3ZrcOWDt3k7XnnM24of40qdb+6qeWNaOPdffMF4eQy0zqj/3W/bTCdYSwqU2uKly7WKzNE
Dt91qeJ/eQ2ViWzsDca8+W8PSDFT0nM1wzrnDFmjaWzQQnE1BpmsyuDTBdrZOmUz4fkDDQnE+5dG
Rj7+2vIj2JmHlw8N/hT4yglUTrK5Z9rNeWPHrdOErqtYNpj1Ww5bQf6MvhbSJ8Ub2sJrt2m7+4JU
YAlEBkL1jh4XjkOz+33+pYotBNs8I9vs4jebOBUYlDt8T+VlnRQMmLeLHd2ZpdVBY+QqV4qBeeDU
zwFO13z4+Z7tmYfKASPesMItbwHOP9oe/1khUjoP1qZC94n0kLv/zgaJsTt+d5XznOsLolgBHFQV
WMmEoVPbxktecUYuyOuSwHA1xcUloDv9lIVmvw3xvHoyIt3TlLrIzdnGSPF7HWZaC49RpYgTHQaj
T+QIup1oHVI689OBReQCcQ8uqR7pWaMI6l1bmfF1WaBK96M4NDpzEnLTQEC6B2euEigeXmUMbIps
OLbM//lDn7TRgwy6muabuCo9DDQhm1T0HdRkvzaCEF96L2NaCe/ivfLyTQW2JKEEddXgAaz3PlU4
jMfYFFWLgwTBT6KzFX2J8H0zVJNL6g54BKLPjWiDH218fo03fe6XxJ+F5/zyTOzSmoJEdil8+pEh
6ddVWN4PHDyMtS6OiwZynuTtfi0zWK2JZvzpsPU+KUFelOjxtDg5OJO7iUSpBebN92nV/hKo+8lg
wVzXPLyCTOie49qaXc1eMAn4px1dPg9AXre/L8zfAIxx92rSlNXGNdpxBi8B7JplUSaezzCgzCJt
ADye5JJLdTMFU/ZlIN2eBBKlpFthZddbHFRBlCxN68LtJKzxlpAHB1jrFW6TjsMUtCZiHYKcdZh0
RISTSx6x6f3Io0URF2CLI1bEOiB+osYfuzL3UJ54lw1lQ8Sy+VfV4uoep2JJQr8sVPcmu1MCMcFw
bHbnZeMq2Uo/wDr8cOt9tTdzpI2kQapLAIiHig/ifxE5YXsdyZ1mbBfrzcyYgifNh4u/DyDLVhbr
E5v2oajMlN1VJuiUWBxB6blqcCmG3LPZ1DnMUmlsRVtPP+PDveZWLXAZJxmm45M+XQG4e5dgoup/
OagvSNd6PqRTNW/dpxp9SHh8juNnQmIahVPVQG+6rWLZ2OW3W4Wt9s37IpaHjXuQrxnXu+miodvl
dFaUXgErEqyzb/aMPmZbfIaPiz6qTllW1byfZLhFXAz797SJ320i5U4egTp13wFW+pMq3qKUL6Pn
MchQqsiXwkVqvhd29rIjMHIdhIahw0FLV6Oj61BJDVFHvI8GLoAMxjpWbDim+5TMkJ9DUly4+s9N
G7uZnbF8jrd7LZ2y9w0fOi9QxDA/A7bji/yVHxQX0r5Imbe9X3lcsDJrPIx4ZMMBR6mGs0ce9EVI
3+WT+BIeOVBVbYeKgLBDucQlqKaeN3tl5qhwEp2sbkO7/0m+SFCuULWNXUATyN8gkYXZpjBQ2cJa
M/4FQ/zttueQsHX4W2zjkCOChfMKzpcsWEPhXYsVIfy0eKhb3zdfBUdKxZMMeTQKvlu0vZ8x6GHq
i0uAdLY1u+1vmQ15KHj9oEWOQ9Kb5PieYr4UEtOcSS2TV366i2SeH6FJm6gV9mXuWfniwGJyqpYi
MD5MUq41BZgY+yG0RHxSXQP/trtiAMcWowy+HkcDDXUx2rseKnD1jvcWvmAFCF3v4cqxx8gF4B2q
yMsJr+b2n/NTODrpCO7IDzaFaNFmKoPbrZpHWbBzecSc+d6Lhas4O1wVopsiG39OK7bbr5cDNxmU
3WAJSQC4DWy3ntU/efiUHwMIglMUiGwOu4N8+itVvz7ZDJ1u1vmUpeYL7Rgot7PPJEEK3YLFqeJs
xtwaQ0mt9LueN7BHxkou8HIbvd3jCoqyVan28RR/Ug02poukWZ0k/oKgWTLNIUU7c7hgwb7wt9wu
0gwsqzMVPsq/DNUoH71pB2v3DibTcPwUbwzDYQScEoRDmsFo/c5zVcdVRK1C6il4jWNmtIc6DSMM
laXkLsPVenH/ccrOfEB0sHkavh1ibcFc75+NKuyFGThcDfZYuQkdD8dUCDxF6ZpId7XqJoU0rHbI
y9UlNRe3351l2Sea5zOEOk4J5Ur193m1oE6N1Vu4T2Ly+36J7bOmm2nI8toON/Dil6YjNTKLR4S3
Rd/ZJTZZ5nvTtjv21uOT9w8EcufdrJJkp8iO1+vt4vOpg6iY5J7HRLAjnbNI+N6pInuPrNwqPxbf
Zcr0ix7AiXJ6CF9gl3TgNab6B6DM+4rtuWac87VVIWwlSCqbSHE2ZCQ4UEO2eZ/G4fqMklYE9l9M
QIZMUxHQZOvTgzqhtzM57Pu50+iiFFqyzKkI4SsTkUucb9nZbTg/sA8jqtSATVVKdlXPSpYzUu2b
/g8yDUtzJfgFLGBjeUvWz86pjPUVSxe8ebPAhuOHsL0AvrZuY3pzC2G6noJye+p4oOuSCy+K+iEw
pkfesqQ/HswLawl6zaLMXUikduIvZw8LNCrsPYuyWBe/xyP7boKN783kypLuEEZGGoOc1GFIBn+V
PoIbtLWBCFk0xYQjuaCDjAnCKBWFGKsAcYhGMYEdvmjAXG4QrDl0Nud/G5zR4Ceq+0xgbNRMPGyT
eOIz/zAdngiCuXb/b4P4acArC47OzSfMn9Gh4DXqcgyb8DHJd6LpAD6WjeD+JLCWGzDpspukN5eg
phhJ1I6v2uPllKPvPqbcOn2hhyLWte1tKdHUQosnGYsLSgA6ELF6LEGy+VlOJgIiKR1r7ON27a33
iuZPBfyniSLgXEq2I1DK7V6R/GOEbCdEabmdKcvv7rkkuhZjmSVaQeBg2JS/fCNDwa1MoTYsTa5y
GDruVSEErKIuPITe/AkogflJMADtStpXCLd+mBSyVEd2JJRVYBb+rsCEnzVtoSxLNl/BoHHXaoXN
uZpc9fGbDuhrle1NsqfbMAcWqRlSVR5f9b6d6jePncO924W4h2P4/vZXIHe7WWMoigAYeEsTyXr3
ZkBGtYOwk08Pfz6HaD+3hqtD4cLc4hCp8PO2BEsjOmgVEbnBbO0XbzuTv+QFVIt5lOm9F7m2yFQF
gGF3zJYwp5vVGuJSb0kmnat4QbrOHAdpCR3NQANrfzNiUG5v0YOvOpPKc7AMYKkL7NjIPcWhXe41
5yuzPFROVsmSQgmBXLh0ZpBQTNpSkGTgIbTMi6udQNpjHHZo0fjc7I+Y/dqMgSkhVBDHSqL1RNz+
Kew4JK7Kpnqzabw93nA0Ap1+u/8kmx36b+OvWD1grEzXkyZtMyoTB06utRDBrkGBVQSuiPy5HkAm
YDzZY1AnNA8wCnDM3FXr6ZZmKZsOz7LDwlP84FjljF15uq8gZu1QTvSXIt/NinELjEjz1mgNHxzt
cX8TtKsTN79VVdg/wRbkBGEN649D8hduzvxlhU7TsPrF5i2Yxxgzu/ZTvhFvQPD3bmGUVnctM1+O
WJVJM84t5sy+wNcJjf5O/4+IcRpxd1oAIBDl6YYxoeYZKB0U/7EmVeYGO9a5urkGegXi7ypqAf2A
ohuMbHuFsDWhptvTy3uCx5OhEOzDZKC+Np1xJnUGBL2nawclZp/XRfA8XByImSYQKsJ1xHlqPuE3
c9QLquLvjG+POS6jzwcFicBCRlyDO59cLpXZyqWlL5RcRXy+Om1ojs1fE5lKOZoxHst+I9xHYK20
FY2t+9GjaxipTAEREhcrZbcCg+GoksRUxlVqWS1SpSZUHx+wywpxW/JOdWlASfWAmEiqEuDwKWTP
OtSSKCXvUo7r3UGGEHIWxUNsRbkL2fa9i5Z1VDEfjJuM4sK/HS4gi8rOQJVqc9eC7oh8AZX+YHIT
zPY/sR8uNMBOIbH6MgeqRjKtvhpNgksJWbtLg7qazqLwWnmMYcorEHXqkV28k5ZgDlwfUdDpnHqI
pVvz+oeNzF+6/eJf7qkYOtppBNK2ARyTAe6R+43c8lWv/rsYZ27odqd4v7ww/ug5jJELmNeuuy4N
PepM+cvmh7B2FNBtFnJNSWhEsNDlz1PNkByTdyS+NklhMXdXNJjuJJnHlry0AA7RH0aScnyAL/Sq
MhGfC8IQhf17OiluBVk85aWHJlRYRuoT2oGiy1Y8lzHxqPNsvqC8Q5tUkbqvIV+aEiaI3LAowggK
sevDoyN/86Ah7pJtmy8J5spX0tDMn03uERYimIdnAB6GvZS253oHtpFczAtkppPBaiuHIH0qaZ2j
3MTXem7aa+kISXUcIskFEphNeovXNGojlTLLWF0kjgXoYTlE0W8+fYxBIQ+NEuSGjIWgTZcIA7Sk
ZkoYdc7ViJbO/o/p2gD7aR/BQ+bDFOuLFHMHqTDvA1vE46CNXtSpxJh1lNuRPagusEmCUuh4OSY1
V5XMGuHB6EGGw4NX1TsNM2BPOFv7IdJC1iH1LLzIrO6Z3CKtdtL/uiy9Mrfo0DUcIYjb0VyDW/Pn
z/GlMhwfcAkkXpsJ8Fb3i4OfxLCGr+xLHGpto9+kiE6phHzHN3eHrYTiCFbAUMn49Ui/3ZwyElGM
Jm5FiI0baV8q3X+Rg7fSVIT848tpaZq2UxgtIirleHfqc1tSegh3aKEXlRAvt3PFTrxO3vMjBXaD
G8N6PsAgZgGGWYf84HCj83oGTUTUKWWq2sz2FQ7fxzZs2jdemFF5ItF3O+Fkqvn3dQf3v7J6RGzZ
TEwvZuqQ/xQlDUTNyLlt+1D0mMS63z5kMnASKSsNFF8pZGWRWqjmdMGDQBWaoYb+naV4woCZuVgL
jk8uaj5iNSJPEM7/5ySkuR9F8RWnD2ub/4e5dQyET2RbBGidlvf+7UlIwpLuzsDvI2kn/+R7ZgvY
Ced8VKNqKSf+Eea+pqF/gbyJWbpxE13nVqM4V1mtW/vQkKIQS1PIAb4X3Bd9f1DO7sdso8aGyI0q
0vh4hZGDWQ4Ari6i0sghs0Y0V6f0KO0VTMKHcU+zB8ux82NfNK4R7PcGlPtC6uiS+o/3QTbCBuaG
vATTj0P/5qbN5u4FBYdYJVSH3dXyrvCE5ScGz3wT43lzXGBky9hLpsimSDR/XCqArbYEL6KyqUj9
9tzSqg3WjKM6sErpNCjfYJuipTc+OyQ3BXqp35KsqB6752WIcMoCZRoQb6haexosTF6ILcOQccY+
zoMiVXuik8VcgeAX8Ra4zOFAEK/8FHpNDQplkfsSJ53xQDfjp2o2vZjiOCRZtTT86O7N3wUBQqSJ
yFBQlBNpUsxkb/dWwzn3HRXYfZfFIxBuZEQIAFM213TaQQas8zh3VbKseIo/JazV8yJ1x2hTWzx1
KblyiKPDlsUsoGiMGYhHnCfiADKOs7PXQ1MGtL73Z19h7oODTjT6kYNuStzMYAHIiJaYEfNUIEo+
ZKKHH+Nsiw5nOSUEOw5Fn8IHZINUzX5IMYYj5FxOddgtipAhbzuyaohxzxkz9NMfeVLeYEKsxPZE
lv6T1HVlZUxSSKMTYyU3LLBOPUxZGJZTPYNz100i6NTiwNGuz/CXVulgQj8i0ftCsJ3LuOSNz9hT
mKvm6U68jkVWujcAwg9ozN4rkg9tP1JTWoRFpal8IL1dM5/1nwGZ/Wv98XSeDe1ST7zbaIoBwrq/
IlTLtupdrH+idEpLJYpKm/N7NX7wuyH+u9+1vFpUKsbMOWgi9ekAW4/YCCz/1190fLxXbHL7ahLU
S6NHEpnV1NejELdOA9JgrFemxggV0JsG2dKLtZheQDZ92Tk2mVeIhloR/HChDlpR1/3kSiTayWFe
HL5RI5Pe4MHAS3wUorcIhEajCACd43rIZR89R/aA858kD1aNcGOydhCADaTXC7wpOosMNf+cQpqb
E+5+U3+DtQIWym9Bw6RNgYXWxCByKc5DUAC+2zHXS9QVJnX2FLTz/Xi9fSkOQ6rdpTSBkrhQUMik
lTHSkekzpPXWe7oMdSnxVtlFArqqv8hZ/QPIOEQe9SJ2NLomc+5tqShw4n6x84CaUFnpL9o9FD94
NCe/tXpcAJTKSyizSiuN7xbb6PWOXS2RA8hAsWGo+utWPdcPMHySqo+IS30fVBd3vgySRj/+HK4t
r/EwOFC1Ytem6df18oAMf5LJND5/c/aSc1dg9GpEymfs7BEWS5+VH7lIti8oSy+Ianqw/ShA12Ro
JrNLqq+ERUxS1zlkVktdPJpomsK2LzH7SKcMMuDVYC0TP1V8TFMsuflaTH6CdVZk2Q+JyCOOcmU9
HAJOxzhQ97tYPR4q5JabPx2rguTDM9i2K30d/3DNws7aSFfEI5irGaMu0ftz5xbrHX3Z+3WTeedU
bsOWrZBFUl2xLcGwWZhBzlFJJ9ZiXor9GQG2XijMs+Vabv8EBwTpa0u+P5whhPEre4HuGxuCG1RE
7IGsO7jSZlMsLTRsGMpJ4ZJIO0FxqRamI4nBQeqkNrShYdveDfh6e/AyOQcXcyxO4MiTcbAKhyOn
83uIYYFUhpSdFtEXhb70cFhl+PVDnTga20lKO8gHuxgbxnqETyD0mRL/vMNAay6YnbKgYk+HDpmt
E+j1hSje7sDg6LVIt9zV8FwsuhWAbp2UedH7iZnFJFAQJHkFzc4XZqBBfq+tvHYo+JHV0FNehkEO
tiGSeEtQkAxBIODiiyvqr1A5R5wNwnElZWrSGgZzyyefmOOLWf64dOoqzkSWIfjRiuNewhpS0bi9
IjdPzcAbIiYTxoL5V/ZFiPoJuEqnr6XzNCQDDiYHYw7utuqAYZHW06zABpDXVdICAAb6xlXg/0P7
WsO7rd4HApQa48KXp0aPChuJscwYtAHVUSRJutOBqFJjxsZyjvi08J9sQXrNaNRnmUAHbqZh7vHc
/ZtOsCjqnBi0o6FvCCRlnm9ikYZLZwA2bv8kAm/UcyGm3DgQtxtDPtFTuKB9wUiVegJVWq5Wftvl
UaV4OoZCm9DyqJ7agSIx1CMnlGoQYj/LyX8vf4BYARCY2yIgohjKrTlBH7v40JMVxKICf5HMnRum
XZS3QbaJxjWvw866ung32gK825K9UDvXJOzkMA7HMU6cHX0jsXWlnLmc6+k+fARfkdilDNzqlZkY
ZDo7jIExQNPP1qI2v+b+aYl6wJkkSNjK1hK3VktCTIx5f5XsCfBjBsrZor0F/JEJTzTbc/wXx7iF
55SucG24cN437UM4eKkiZzUAKaVoxN7wCwzqde8Xtf3E9iYY8GJC+AF1oubnhszmTnjs0eGMOMSW
+pkkJ+idc/ztmYUMl3Bail9W1k4Dl28B201tmnR2ChtwNykkd16NRIYURPQ5mhbgNN7aJJO7W2Cf
UhtW0JCKPrboR9serIi4m6VllD6iJIo24majgGQ7axLHL6EBFNO0RIsdvMy5JFg8MFNrCD2ctZ7c
GCjYoqFMEUWQoMEtRvigQWS+q7M1Jm/J4bh5/+pZ67n+GmpmcrF+FnTkBNFAxTIfIKlzES2OChfl
xRwJieeiZ0FSzvQe2lsmY4T13Jp81wYtXNMW2fbbBQLIHC5FswSo6ZnKb4IOI717Eq93mIKTmA3P
sYGKd96/RMcxXcSE0dOfPkeTAukVgfXUBwIFVpAz5/fZFAXDNeWVcBX4pmgkyj/6QUSb5L6ljlhU
7wgM0nnDIR8bJGq84zDbYRJJfRgXKZ3H624WWuEWYiuyocGdMJlmwUHsuZ6896oFRfncUenTSsFR
s1zLFfe4EV9Ugi31yE5ztREvBjndczJO8hAZ4ghTJ6YEo6yh3UaiTHIA5X31CgAwzldVyXB4GSRK
jt1uslFtfAPyWMi3x7P65G3upD5P9RgziZJ8lSd0XlCn+Wp9q3BTHsgTCCO9Jm2ESVo/lppsh6FZ
xz6Jp05e5DLtdqWs+WZw24kU8cQGOZHLEJ472fybwtxuWSNIVR/8nQDcdOw4ERir8LrLXdaUWcxc
f8k0QCvhd6ZMQWasBqSdN/CZKuR4ug5Yeq37dkPG0w9+FcjJEi/As81EpAGe+nnudPkyySEkpRFs
vtU8zJMZ6EkBcuSgCFHnC1ACWLf17J/0eUkAkZwuB6ppIZBqVckiFzP3AIQ5Q9oqHEOpHT+DVnhU
0EJiTXJPZVwYy8NDKDwFc/+uZ+eiR9uBSq5aWcQpimx+ZnjungS0ulUhaOXSLVU3sTFOjl9LKV9P
Nzz5JlnfCcauCtwZeWrVSnqn/sjrg9S1UEXddHVNVh86Lk6qqXi5QUNH5bwsg9J3BcY55XRa1uqu
+LAi3tfeZRGcIsiFmw98+b/DK4PvLA9S+W1lakiHJ0Jgdp93qd0NObtkjND8Z0gbtrn6+YUwbVBV
VrIDTwwW0jgPTIZx+FStOjtDXfly4KV1Vs/kIKlk6rP8LbsDy+5fPYqRcu70KkR78U1Puh9VW9En
CfAqx3D8QEfeoUPCXfXlfblKuQ8UVNnEKK8VOdik9MLuF0CT5KTayWyEqw8s2YPeqFN4EXb9oYDV
hp099KvCtQzg+VGbhLPP3ngGckamqzqTygekzViX/YzOMqOhtTM+CqBuOTv8rIanZHO/XrSbZp+W
8oHkdU/Kf7LlYSAFttsHAoHvRH8uVxh7VHPnnY0ihJwu2Y8U2TLR8134VjbPAp9onXUBPWg/tmdQ
fxpGzDtZb0haGI2VArGS4ngpivBDW052dXAE1ID+CldVVtBtKHxnPlEpLPCernq7D+ahe1cc41qN
DyBaZOXP8xEU92KErzS1uzxryElPccFd/Gh47+qf9P3++wUNLym2fd35RL0JsUhp60dh7JyMHaEA
a7eNvDrj27+lmYMMLnhg2cCr7QntBloEoQ9bKKWBeX/D81KDLbJc+hIRJMoRCbp1V8pw+gVSIboa
lGDN7W4c+C+DWXk0w77g/bfq5k5n982IzYbJsGiwcamxmLiOBGizdG9h4loBvuw2gB8Z0CKqW8x/
nJM/FsEtKGL5OIc64h8PRPy/6PZQ4wnxvomUSkykI1jsAsKkEQLb1wBuiO6ZuaHiQS6TEJgup3E6
6ntf06nG1uiRK2RZnTbHnsPC8BiMFQVXccvyAAVFpUGSriN2YUc1ZgCaVuRA+GqKfipyOPhbuWdR
k6RQJukZ1LBTbEY/kguZ5XeMMZXVUfH0kpkW4Mev1S3vPjsN+A6l6MVDWSZ5rYY9LPUKENzaR1TP
/zMbD8NJHkGzThKZKfXNgYqiSKyrAjnd0Cbkp1io9bKw70qcAzCCQ3y9yGBDRM+3saBb3begX9B7
Iwh8bVbWtGs6q/dXA6xiUihZ4dpc0v6vE9RkAP1lw2e4ceFuxx/l9NJcRt/gVo0ExJSUWcBzliE8
epLD2ynW1LyJgEAmGQSr6P+nD5urdLxpTxnG5umfa0nkJIG3PqCcsYXLgwFKdgAeoWFeQerOwKy7
b0bKm11mzhyvRH+Vyjq4gN1UZatOlpnhVIfA2Mgc9ygwl3NE1IaS/JxWFOrMLFDPkKgsCmbAxBoJ
9qy5CFZjZgcVYIqROYH9xw+YgzSuivrS4HdlrnMss35ZOee+T8Tdis9zEn8J07rUJwv7OpEXld2o
ntpfBa1WL5EwuN0YVIpebyM9BZq7Xq7qU3t2LFW+AxMnwIT3cqm1IPQbXwKXCCDU3EDQxRtnfwhs
EE5B1tjr21CxJMXDMfs2dL8CRv23XPHYJlsbxVRyzx5o2QFDtpQiISO317I7Uy7VAgX6hqMlo5f0
WpPgJprG/Ay/Gf0pKSw6s02a5WaF/Z/aC7f+hnhN7n3dvHAARP0tYJmZ5Obk+aWQVFBevr/5WMNX
NvRzUIN83h3H4PXzJZFe7LCpmc/65Gq4ngbTps2h4t+wmhegleeeSo+PXtAhL4ODP6Ze8LSz1uV/
xo0AN9j7/ca+rFcNjFaibUy/9dAQvDd05K8Z7A40645Z9EP6VFZVnNScog3m7VNQWMGHKUTstoud
KDIUdZPmiWIrr3NipBP1a98VKJ0bl41ap3C7CeDAZWHt6S/onFRThppBWWEOeo/V9TcgwW/wamYs
NVYdV1OpfLA/nGGqgs+4w+PmzN3jJMLhplUX9nqQhl0x9JfsHYPy++17mZOUO1hEJXDAxdBC7mhQ
vPKzhr/zplr39Fscx+epvGovyhbWcD8DK2Krfv+D8B7QF/HResodYGG+aTmDlhewkyDIRN80OgVk
2a+hugGKDKXJf3dT5OvvkI61eGz4L1zLHJq7DiIATF9tmLn866cYyfcPITQ4Y07n1cEO6zXjEcKZ
TIGqO5eOdpindQN4rnq8gS+Qk4l1I5FZknTi+qGXEQVJWAdmAEzQOZy43DKx33XQOPOtM6Y+hJfA
FNvxZMQWEnPZzm+fFfJlayz2zb6cH5npxa412U+gikudcWMMzoyp9EniuSSQgtnNgNq8AYSDusgN
ywh8apR36mCjh1+VmrW3o8UTaVBhcv73+XLsTaQZ61EhVqLXLZjG0pLzjUSPJ7y7rRtIE4NDURTn
n7k+BOOfcxRW40GCpiiYtgp0ku3RwgsYmkLOTW5wCrQSWjhRKOEFdmkGSFte31iorZLwjHma2ZEs
ZdGHrsNT2+Ejta/8MI0Nv0mesCGy4SQvl1wSeWFDzg7zePpdTAbtWFu39xSv9Is6CfEtiS241lDf
oHj8xTPgAGX820RiJL1fp49CW8GFDgYq3pzlp9qjL4t101lp4t5FPCYqa8zTV7nHPvaI70MYAlfb
cWEPndgkir4s5qmfAZLQcSSsf154uWl+1vahGektZAsAIOW4BoE2SE5oJ26L6lGbPkLGsyWZHZd1
BjR4dFVkr3dAD/sGTzS9gA53+aR1uuvYUIpLwZreMAErmbhNu4JjQhyWyxRHhUkCck58iez+POon
T2d0B1WqLkHOmZtbH+eKpNHHqyJfoTbc+82LW9/eKunpQrqeJtamxry8zO8ilrO2P320XSBB25/G
9L014t8PYmE2iNa4rbgL+2bpcfVMpjf5B5d2dr9nnzmQAa6jKcSbg0fHnSNi1vo1zmiEaqLRpv3E
2KmorpIGInHjATNQNl2UXxlvJo283L/5yPqodJxyn+aANLdta+bMkDaFRNwZbFX5RrgbVkE3s0uS
ZVp8cbk5KXLZPn6Id44PkcKNpZr/zivDP+t3SIdFdXs5G3UoAw8dCQgrLydjuqWZd45RqA2kF4uv
4Rl1/lPyRufdMt+AoNHziux+o6NoiJt3ekrcfK+PZBqjSSLz6TzvWO2ZJ1DETMJu7rJF14TrH02S
5EyudSexW3iahg4+mpx34CCP+zGuymBpn0mmqEAGii2QqWzOQhwiFreHYB1lTo+EWywQvXCOK9vW
jCYbiSII04AC4oP3aHsbhbaSE9FfePyW11gzE+dDWSBQvPFVyGAZoPGUz2rBSiEOQFkPUEzISl/6
/Z6iJ77w4ESoh3M89mi/deiHJVugIRFILM55mZFWofh9IkO2jS9ojQdGnFlDRTA9K30az165T6gU
hAwB/sAaqrPIoHl2ZQr84WbzkhnpzifqM8Te1eWhMMix+L3zccNz6e75Y/1+0eEzn98w0xqOtUag
Dv4Ef7Ugphb3Afx4Zu8s7WE4QlgTOGPBz8bysH28mhRq5KCwKnR0iCg5sCtOmEZSzSuftRLY59Vr
kjPGtFtYIP8O6RrckzOgWuOIK2ZrYmlGI6jB6R5X+GPRMi6sZPUf3PI+8E2oVdseBG/fnE9bBCKP
IwHDEWdeyuu/fzeUzIOzVPyT4Qm9uIL/xbuWhyW95Mf2YfSSsOfefRJE0GePK1WJLCpqL/jpMjyy
sHO93mf0EMYMEg4vLcn5Op/f7ytxAHTFPP/3du59etRePGKOtcdUVnY0EMNyDFKZNQ7K0yL+WzB9
NI0TcpKSrcV1jFDBwYhBEyCiZlTfIkeKr3N/wLicOSULRBqd819DjEcjso04jpygRwz6p5X5R6dk
6V2AOKXOgjU8VGX5T+0yXvMsirS4ZZWI0p6SiVXwmNHGDoWKHwSr7NmuAS9yVv3KdmOElTpOpUPy
h9utVDvjm4ZveWzCPV2WhwTkEzQ/xc+KXNCwT1dTvu9CWKiKiDnoLCwf/eEBKh2NQoidn8aBvnEC
RRkbkrT/+FEsV7+CzksfEF8l2gaDzp+OMt7QdRqHq0rvZ91c51LsixgWGr6GgXJj5G4EXAg0BB2C
7jRm8Z25OdZBSJO9QB6i5WPzJ00p3SYmOECVmttQjPfKQlClVTxxiptYoobrSzgkNKIBMHS2mcJE
KUXtTxf9dXPTSk0GmMwz6LRKfOaRK7OMqxM9xqPdNE0+T3Tyy/vwtFcA6JhTJYvXOQ4mpXyZ+/wO
13x1zGocdGldHBkIoghG1ZVWykZ29C0M++z01cw3PLvAF0b+6poKASp4cyXElcE2KY4760Z6bX+9
xvd+zCbQmIBkiSVuMYQ8slkDtAp5LENE20CAFvBvKvbmLaSwCmyWYPdmT/Iycqi/KKqD8FgUtCW8
tAW3+EuMq+lB3S47AMsIF79RuUdyAaUe6+3fhrw4f5pkA//U+T4S6fY7vGxy5upuqGKn35X4YK3I
GXjmqyFxUFzwIDvxXb3HJSJkVAqgt78Rklsybj77QYZ+qHjU78+EvwBlPkU4uT20O2QDJipTOgXr
YFEQl1xdTQZ2UvK52QEub4Wu9aCqbfzCafpkpSBaZXRbuumJlk/CBHk6lWNolHoFhQbKRkZp6Lwv
eFB+S2rJ7X3nbjFrbKOVr/Xg7ggyrmJMH1hJWaNSQdnSfMnmdNOXLD+h940CO349BD0qY71IxhGj
QejhVC/0Dp5SAWXUFlsnWu18vjv/pt+Tvgzo9tfGLnp6W1mUFZhWbUqjWzx8m8XIH6pCG0eqASm/
stlOX2PDJaGLacYFsEJIJi0DCV3uaJWftS1X5z/JfrCltd1K2K8LXDzo61vj2ohGDAJaR9JNkcOY
9AmasZn79WrusP/lr1yIIM/78HZu40ge1wKS7eFTXdLvW0Dy5vH2hGBmT2Y9KbWYTq/ppagUVy2E
tgiFbTv6hj32EZXBjWlgDNfK8cNxsPp7Y1Ug37Z8TrgSC+iyF6/uaVOngPAPLgRupWEl/BkgmarG
nrKq0UVlXLkrv4nA6HLxeu+Hym4pSdlZYirGHLiH+C9CXzIwShrkHqWRISQTdFAI3QRG/ApxRHvB
IrVBBJqQAUqkVpag/4IMkg8d3OKQjSUyxGWDOzvmhLMGR2eC0olFxks16EPQXzIuCAMTNNIr7pvi
X+vKWzx3VGn3IEOnSB8HehWlRwuAGjVtBX+Ke63COmvGeMCH1fgPGkLVhQ34dID0RTaFXSeIjrta
PosWNLJNPu0tkNIVuykn08iDOs70uUOY+q9lwQC9sj83XZQp3mhFdf5D5v9ZNc9TZ2+KgHvOXrBQ
1LbYOz0CH2rw2Lmv9SB1FvbnEkJV14xln1tNWeIscARxw5hwBezwnmNZXs1nOMeFrq6gJNlMRfTP
oiUKG/Trvqke2bRTdJ+1/M8pU8RGeKKfuDsJ7HRaCM/z40Z6b8uZ1VsDV38NWqK3ssKWeuOFb957
+EdqyQqrptk72w/6v3GoqUruayML1sBzCs5aM1EPs0ZYyIIjNlGDUTCE0BqSZgxsvAboN/LfgH5F
tdKEVKEQAwFpdxQ4KsyXDsQhrcN2R2cCK33yTFO9lpT2GBG2zhdzNG94cAQqCLt/yC/7DAjNsHlq
gYAVLKA+v/XMfcLEvF1TOfIFfACqhJiu4NnPSav2L1lKghgroyzvZ7sN+sU/tfmVNj3n0JX1/Qq1
QDRmxo79EYeahcoXcC+j3hYG/JZv3yZrjUf6JZ9E5itYapX5wTHi/nAzigtiWLF+qwFnhpuKAg9O
+Ez7THTwQa/ITlK1ZUXfFTgOkxDYzwAJcV4HuwSHmzYqQstzFK6p3kTRKIy6h07l7BPMGGCnCxsL
+SsrYk32CvoHfqlRBvERKwiJgNZBSK6pcBe9Jw+q/QR6OxxqWkzCi33e5JDs/1gXQmgeeYWc6PsY
uaHtgmJZSunwJt6YoYn3fxGj2I1E3l+YNWWpp60sIo2BE/FP/8bLfvOKmJt6YBvsHOfLdH9Dpvma
7uzhO5vHBLetjdd8cpcKBwZMYk5kiGaHMa3ogVKFwqaK+RtbOXJmXpuR4g5rjE+vNVHl8slTBCaX
C/zQCGGZofZfYGmdQ9KI+E2oUDodG0IkscSxzINt9yE9FemvCFq+X5Ijj1PRyq1pc8twlA8LQvNh
MVfihW85WxlVXZdrEXmaPs3WFIUMNhIzEQvKWbqRGyYlF6JmfNd3JlijvP9JdV2LUOttxuBnz1+7
1vfhbXIOrMcQZO7aJ8ylxUR4SewoKIr5OXypovkw1beTurfgx7hBjYLOZk+MVCyxr0ojqvv8QCZb
ne5di0zbljw/jxPZYiOOg/nUsJvZQDMSIfW8DuNhpV8jsqLsQlo4l5fj6mrhQy3R0i9WH5Cu7nLs
ee3PnMK5P7feS0IZ7D9iMqTYx6V302JiCAgX912YUIibXMtuKI8m6G5zkTG+ms8JgW4t+ezVlHZ6
TxCdTlQOiiyOuxPagiKqXuS/2Lgyj9Q7jtw+mJMHaTrGg0E4qKUoTC9NyOD0BSCykfpPdYQk/17O
1yJJOWgXU40SdLZ59SjyELbbvdn6T8kkciNB7umkm6autlc5yysTucDVM3rkGX2+OfOkHP2e/2a8
PHWxceHRIV8F5yv2rzgNTHeiAGn8b+InrabE+qJwID1RG2O2Ch/stSmhk7J0YXsdvn2FFi4mtXvf
0IFMlUXWhFaC3PMibVGpctA/eOAEOSIUS4ssNe5/jSTzFFa6DzYKFtwbTCNxeHavff5PBPS1/st4
qRhOTZbvAvxHbFxbMDnqgFnMhOedLx10rsGHQQk+9UNmYOq22HiVaE6JQze6tZ3pJPgLcRAkeuY/
v8whENdZOHd0gwwphgNYl7iSO5DyRIXCNOgceXwxEAuNSOPMjkIuQl/AL3zMf4Z8I91N3ozPwI9Y
cElN0NneZFgoReu8nNRd5b2KZoIk5Vx9b5abMmz4VVItdiIsKJ36euGPHQ0eR6Qxjh/Qnx5ZqEJf
maTFhpGvUfTrAOI5pbwpALvWqkeabJEVL1g3brsMoM+ViquD/2LF0GSvLB5EOkwxtY9OhbRbJZUC
wAv+gx5wdg3VwEWirCoKGGyfOKbhstv6CEHSkrV7iMFKJdXr+VYDZQuuTH5X8+Np2ftTDhi15AJ5
83QYljNR0JNLAZiK4XGhe92rXOZDuf3FNUGjJFFyBGwrLRXkeBfFhvy2c8Kjw/G0zKK+8mHS65QL
nrIkQ0hJctOt3SCS+outSP4iN6m+GnaP9JwgFQwbAJf/HN/sT8KdRoVWovI0bVv+mhnV/X93bRji
1PTQ2wgyFeUvbp2NJOSMQCuWEMgCerPK87AvrOcCEVXcJBGUa5wYa7j6dhcR70kyM9lh+Ihm4/Fq
GLXQCLmsQyv/sOFvUCj+teDzopjPzz/wdmOLbzyBy+bymcgtMI6KTANbCry+ChOoJy9rhIASRZMm
LSb7/PDnvTGTuvJwYUzpoKG7SXgVNQcgZHHJeKi/GYHmxqAkVV+XQRBkwlvkdsHoKnf3VLhWy/RV
ZwKRNMh0/kPDc/pXQzHs8zLngDH9GDVLlXoo/2c83rZuttEjQG6x0BBK8c5BsBmlXXXUDXHz+dZt
jfgNHi01NqnUu8+qZ9UniY07iVG0RFMVDQQ+V3LfDhEZ/h9XlFndfzc/4pn038gi67psxyvc3BZs
HAzoL++Mt0e5FNL02Zb6n/gQlyjtivEaQtLpaBB5do1Sqs46+/2WT9RuNJeHSjlQFmOt8whD9wXf
G1ktghLT+Krqct97Fep5L2U8WSFjqLZRZN3n3sv6qzAzUQ+PKNjdwswHRzHfCC7/KFCuwc6MXunn
+ZzkKmdXwwdn6JJ73tIrSMS6Cw5bmam6Q5n8w4VNrQ9fv6wswa9csHlWopn2YaFMKlQSNRVuGm1K
WJo0bnEkgPhEHR2ytfCKJwh96pKR0F4P3U67OQl/z2Uks4WiMNrK2rO4fPN2USv+gwftf0N1+tZH
IMlbtFtA5/s24gJvynRTtOzuPE8/v1B+0bWDpPqzLiTy2dYaeB9ayTwkfS4clR/Q8cpRwtkva3aK
4xRA7NOlLmlWuXSporKDxyamQBn9EY9+wgmcbpF3Yv2XW/JGzjLrHhQCsQkuabJtXufHvJpnIX4l
AvgWV6IYCo1J+N9ZJdb6mhVesBhDeffiWlgrpTCcAAQdBNZ9MMfpHEIkMXDqrI/sHW7EYld4ZQxh
tTceOYv6s9SoNeK/YVoe7JjaGNO5YvYUNqcB0PaqFrIC9a1ClbaRBnCgVxJ50sCGVKh44KJ+lcjW
b8ayNvIeIfdHyh5BGL1CSPCYEZpLRVf1qxVgq+XRRltEo0XJJmHZJkHRhvzF7DB3I94gjZwJ1DgT
gm2OzE26qv+iYO2zHyIJFLRQmWczoU7S9SeG6TkCoh8BuMfKXgtXuYrv7JJLK+901HOgA7BQEOwR
ib4+X7Dkm7jXySqZHq4sx2TvYReDR8dlGNgdb9rkyjfchVJp2x0ly7rP2+vJ6R55eWGreavXlH/S
kuRDHAAioX9HXaC4YXGOdwvKxu53BoganskQpHOqXaX6gQe+y0GPyVrTV/Dza4QxN+/RIILBMKLH
fSqVDPqS2FCIUbe8c3YRCyYO+C7ED97pS8m26b8mqws7pfPtrm+DZbEhC9+EhJ9PjaGTvHMVHbe5
71ULumjtZ6JqF20/bUaW+61UvDqJlnBzn0GFtbFIGYtktUa2oVCVkzBRqLS1IRB/GsCTbAT1OJsf
h+IDzf7Kc3VTf9oI4uXKB5PbH3zNRIhKxTnrfM0wEZHuwls69B+DdB/rxoMVXxDdVUCdY9WO6yR/
s4ubNd+NzRxUyeYtzEZsXBUC/VG5jVAIZhacWujL1riEXBc/k1tpbhYgeeJZbYHOw5XstjZWlOEI
XC30mwUnOfH7Y2lVKkdF/qADw8Wf9PLNQEU9fdGRAvpSlgLfZ6cYKsSEe5wTEQhSZgdcOTL0RMi4
xw666DUYGdgaSTNgYr2NeAvzvSil7K3Q08QEo1uC8lQejkpdZ9XUQwkpnSPXnCRaRaPoUEHGRvw7
BUvEn9+fUL0vY924hu3s8noBHX4Ea1XVJXUq7CJjT0L0GuPqCx9zq1CaA56KlqnlTMA5E6D4amP0
ix2t2GXpPZOxNyUV7oRBtvogu1EzjWIZ0kXSajZHasFIkdQPGUIleKAT+mROM6fqAbCSIC5mg4NN
UphRlVCHKzbDRPiYAJ9x+E9yudlk7urm+M6xu34oNndvRtM0z6/ZMUl9bb1KMwfRrY3s4bXn6od2
OXBqwvl/XtaKFbTh3yW4dgC6SkVYd/Qp4uWX7pK+BySBKwQx5kvYOGSAvxSPlw0pEtr0uSpBRjEM
Q6s3ccAixSfte9zM7dE+ATTEksw+ddpaWAk48hYUYtQfHg3XmuKpdbiXc6kpurpnYoHrWBl+Jog9
MARkQEo0L3KuJki9oVOo//Fu032JGdXJ0aowt0hdGW6sBwFQasgKMkyH2lHjx85ozdBRuXgHZPwo
mmzOC2D9oywABrV2pw7Pl3ZhCb6oAVyMUR8/BBaV8As78MWuVDd7y6yvmy8DiJbSTcxC2mqd9U9B
Ct1lB5pOPpHRkj4wx0vYFl2uowE++VgCN7X8jQT0XYWTydnVM2WYDhUU8+x9VQapk5MeAdEUflYq
1ajB0HTq2MUz3QquARdFrtppfRoyKsH0cmJsBR/rLCTSJNmsRf9TE80dqjkxwfa8WSkDuXXutpEa
7G9Q6GhDbotDjwR7U1K587joCTE6iVB+bgX0E5FXDiJv41NstX0xjW84dcSvsQCvZ4rDU5KFxS9l
uIIE3mlftU5V1hzu9J+jezukiT0m3foeph4UOw1er9y9TFutIl3JGl1Am75Ecplc4vNh3uPBHO3U
+zt5Wa32VigmqZ/A3XE8ONtjxR/uZcOdPAPEYT9sc1BMl7IHV3yXuKZvcnZ+sWQmSTLK6iu/MOWP
VLM/6DSa12maSsSVBxQ+ExP5VEdfUhSoRXGbHhq8BGI+6imxhELW4+MxOlhEw3yqK0ytRnFpbUYh
By6GXUfpWRa+BCUgswKWWgyK+Z6Pn6lXLLVSdVdcrqVTIYlDYQRP1jaGEWLJWcqYW+hIeB/4o2y4
dIqOfetLermLK4s6S16ZvSWxv/9I5btpDI211B8i6CzeeblY8/jHQ0VK20i7awb2Bpu6UuOqyKTM
CfNKV6yhRKPhkKQcHTXN/1YXXewlfnIjOWsXEh7MgjoOGU6MfeWkDvhydR8tLxA5HK++mu618/AV
pizntKF7lbccm3R8TdRhxZCvis3DoJARzJY0WiVrEZulbScPjLpK5uOY6oGSZaQEgo14uDUdJQNT
wKqreFpRFXlAO6o/IB/QdiiAWrLhajj+pItrkskjPhfXx9GZIa8EC2f4JwG506ilkwf/cN/C/9lk
2XZ+16zPb67wPPs/kIKiIM3WGEuZ8TOmfxrrRTVKEqhiQMpeRe1YXE0zMg0qQlQ1ye0G1Ls2x/Za
96SANVjHQ6Cs42pR35DdlsdhZeoweYjkv4DPMz0EfQGJdweFf/tBTFD9fTCH+ybyiN63brS8qQPV
2qG55qARWUpFKEq+ydp/1wuU/MyNQt+83BzBMdxTyIwn+7UQA7ik5BXOsNoGtpUurjuMfMqMRv6s
Bk9kKfkHi809Dpf+BTGZCRNu12WmIhSCr77SKT6JFuNSU5resAViqFPwVjJLTL+mL9CNFKBS1ANq
5sRVozGhfKfZYlPnySeV56hdkvqrI5Nrck+ZQi5NavX9dCWnFyfkE/MxeyQ0sRR/0L/eridgOTKp
9A3K1ybCdSMIOQwOH0Un410CVlskm/jkANU4j0qg0Z7c8H8PdOqDE9jN7XQjZ2F1P7jPeD+flg/y
vDDIP4ohE337CLm/ixCLSOL59dUDMf3K7XLg2WfWAn8sDNUv+u7Dva6CFnodq/rPfHjwmc4kIDnD
vFyDoXTTTO2cFMI7/BKpWVW69BWJEClW4RKMOmRlDFKl5Mqn+9tl7dbA1gxJptj0NfeUlnbZM32p
kIuZw5AhwiOAS9suzJ76NbYAb0uQ8CrJnvFYDvanlmfIn5ZLxFbnKWry/7FzBdJz1Db7xfX4nsPZ
p45sDB0Kyp/VBFBKA9sef2pdZIucHX7hBYuvDsUKicOTi2UZb8JwTUwh/yj3BRFuDagExjZLH72U
zuf9qYAuz9P3WFjiizrr8ItFk3Iv4VcWkVmZVT4nvYTSVFWbfquKxVFEZIhdfGeJuqUAhYpbt9fY
OEVmGx5k6XlSkPtWgTCKKfkB4Mlu1x+tyPDMLK5dYaMtQdV+kQuW6pmFfp8ov3OxYQu8aJ3dhYIi
PPimmSrUXfeuloHSwNJxf+cZ37J/KaoFkeS2ElJYkH/NsOMOdsd+KsxwjtSD48dOOYubf/ZyJazU
7G6wrFeuQwn1EwhtkAsBOQcPin8CWYnLV0SYppRKeQKEOkUvHQFDN5gaKcpACu3UgctpnWKyAtqN
f302d17WEsfaS5LpKnnj7Mstu4dmJbW3jItQO8Wj4hyX9VmpWLTYyX+T3znPq/g+LJgaO+uj4tB7
8g+sCi/dHVq74AEoDSO0UZExiNoY0kS2q6kktNdcL7SU2gFIqM5qWCl2+6RShTd6+FSBLs/eYIIz
o4ADvmnzGwhXi0s0xyPgSAgInyrsfDfixbe1tj0q/aqSZ6rRjvzVcsrtjBRfcBhXr/prfZyylkO7
KuuvzGiTZg2wOXRHzdt0e4xkchRR4GJaBupPqVFrnx+U9JcuZdEW3QT5kz8Y9aj/iGKiNjsqPqH3
xyHGh4eaQ0sFTBDqe8NQ5ou3RN8uuDQjgKoZMoeFA12wNB7fNV1lnUYmzwShb3b59ylTk6WzH0yb
tLRuUJinWZX+GrbvIQJ8qQVs6L7PpsGzkSwoIYqxuFGbyNEJahwO85dFjDVH5END/f1ui3sU9C0A
2xRfNEX8bsEZ5/ZCGyh6AsLciTTUHT7WHIFvGdNiUPXF1Oz/CLNYrzon9krjQwPHXki4suPoNm7q
NQOQj2L2t5FPPHs9kiPA8m10pPGJt5lmQQdeYVrEWzqnaukpAYMmuETmrYoWkcd6OvBJImxOsOUP
2YpoTc9+elvPTSlNGnlULqpAjv6QdBr859wt588/pAvcrlmiPiCTJPKkqUmVl0/cXVq/KBOkUMJ9
8fitdz/imORhlDbL7Mp38C6jBrsW2flNlYMVODec0eNIVXzdMzl+vvYNpfpUD0mrD+G+5CWBG0kq
4FeU98PZeH1Z7nL1F2Nhj0e6NzeO37Gxsk599Ob9tJsfjCAeYynKkGQ6ngzTlCbKQDqVYhq+WegW
DWNyjNvDG4NP5JgFyx7DeITuI+oNz7JTSzSx9Ha7yLKZ19fb2GOCR1kJLIvscIqvWu9NqMkb3l4t
7yGOVq2jCkqrfeafUAyC7FsBeSd8P4trV/SrhzbzTnxPPnBL06jfa3YEIfQpfhkXNxS1jOFWtGhp
6Ojw1g8lyDv0EbQEdIyGEymbHjGaz/viok0BC2G89fkKdj1d8fmqp0AFJF7EN3DFwoPE5zcEJnnT
Iv3e9T7wOcxvB7R3Cfp7iaaOkQteWi51K+kkF+OTOlQP2TgckY2twsD5FOjPs0SsV7/OL1ml51uw
/F/nZUk+oGUFRwMSH2TgdccqfE+aJAD3BYO34OjUOuAGmGl3fCYz/+FdmrEhP47pkmSDqY2nCLkU
4DCeZixD8vBBfFOgvDcqphqdVS2L/mmqOBEs+Ur/5cEX2idmKSZOz2nZaxxjsZpFbLOEgcCRGjID
it1iHsTQYjbH79o3etf5Ccpu1yav69392qeM+s1bEwzOcfFKZJz8tqtpuaq7kF4WueOjwqY5nRBR
LPdSVNrysWzbGQfum0P9PSxv5O0LhVNax1zl7XSNFq57faMCTswOeZ/nxRqwZsaohbEEWRzLd6b+
xGFEjTMTbZSq1oX+A4R/eSXH84ZXl33eR+kODjemgB04JDxAFRhyfEmq23g7WvVHjnlcfsQE9pjC
1InrIXmSKn0Hu3Zu128ld1hEtbYLzlm2Hvr8cAvIgCnlrhP3KU7jDPkWUIemJY2G7N5rTTNVF9gk
pIfs90Ckkl4AZqt4iVR9epDZwXR8whHf/WnaRiDuffob4revtcnmmcEku6nJmMJ+nkL1bYmCXv04
IZ9Yb2elblT5T8uAKHXTyRXzqq4/a7mNd/RLOZSWoK2jEBCF/hTheHBqERcUtdra9tbA1cF8CTPR
FMk5SVwZK8b4d2Nknop4QktMXcASywrMvp/0z0s23Z/TC7Ept9e6t9UFYOo/qPpEo8HG3J6EkLhx
eudtwFsu9St1Ib+3PtNxCvbV7r1DbkWYdqEpDCuoy7xUr1H6Fa/4l2r696KleNrUqZU47NaEvIZr
EB9jYdE+QU/ol8DeAi2lEy5jM/7/CWbR3FHl7fAqgc7tFecj6vPffMCoekb+l2l6OWAmdusenumY
hwALwNKRD4Zip6ingkl/MxCy6lHQifGjtd+NfmV6TS39QCqGkmIO3/ZCglcE294BWd8oBp+W10m0
xXG5x5+Rgu+ytdT3MzqHi3Im8u1scChjkRjObe5B6XvywNAo9+J19890oMTLQQyWm8I+6/OlIVKt
N8NeM0Zk5qKoK07+/rDHxaIPhCXJx9iqAFzqoBSRiWFuKQ+6622li4o+R7AMcRVpqTB4RpMazs+b
nB7DOiyaSPbnXOFLlfUweCkoBEyPvSjXBJtzzrfCxkzmwZ1diZ2/5xHgXcaedj19GM3GV1LawZTc
gd3P7haezMOAbw15U033xsoqf06lc2xhCBHyBSL+HGTpCVd9alUI+0ApA/LfsXLAHtYIFZxFHsaU
WYIpjXal8GD4a9ZxJc9RY/IBC1y4AEKaHXvJx/I5ea5hBw0DpvPWq9dqhUjVhKwbNNdeTIZdDBcB
4RPCEVzBY0DOBEVjLeKC9Fm+4QBgRfx0klSksI79HGVv9VaLRoUt86Kr+zDkUqEVN3NjKsIUN6oh
Ix1PA1WeyQb7AFIIGOImnjK4gEx88b747s8usNCbsoE87+YcAaFUcriIoV7WLEUqYiqC7/d4N+mG
ANstJmgDJpF1ayNtAQ1WiWKqs7bQVNe8XdfRBOk3hNwLNyd8TotJkgzDlqePRdZ7PCSnLnzgGLnY
+8C+RXk3Sns4kdmJB8AbOQsm9gUiJ77Y8X0UN9/ZqyOECTN7QggGmYynhrTcsjZnK8Ylkfs2V3GT
T7HBXE2NxcZ3yH1/ZbKZO2yZPVoBq0PURH6Lqb4g32KbSWMyJKqWpag8K+CLlo9hpSGiQlEH8l9Z
EFEHpVXyNeEdFz9wFAxiPJ42Wda4vqdwMy9GCo8wy9h7ySnkHNbPq7dDYbG+L4EG8+7Sq8ACx58H
QhGj9sHgtFt4d7dn/3F18BvucpNJJQZMjzwjC6C5hSrC9b5OX0x6yMb8urXRNv74zxjsy63DVlGS
UpytnzbPZa5DRnLj2j2qnJ1116KgWDVeHsE9+zWVKdslLdU4ilmHYbJYNbZUyaY5Jdzie6GkaalP
3Zpi61GkVGnqJY95SB0GkyjVkscrSZpJD4wi6TyHeukilsWhFDyq5eGYLMbjbM6wGmnl6gurjRyi
Oc5if6on1QVZF+tUuvVLup/JMfTHZ5V8eugNAoc+zLN/GK85bQlP3ltNtJ8IQHetEM4fD2JUiUoy
C0XjHKnFvgjZYoPPNZlBIucDQRrxO+6oLXZ9+Y1Mm2vZPHyeZ5Pe9nFcsPw9wxvqaaH5rIq0DtsA
iMBE17v8k6sJf1Pty++7uVaPe//AgCFDWQxyrjwfVk3Xao/C+3f42qqYcBqCaSv8xdZjIkGKFpjk
mySoyTJrRHvovO1x9rhd7tc/g7pE5oHyvO2gA7YTkcCvp2VLYf6bQgSy1GgsnY1rdw31xtCjpBUS
wFu9FpnvCUXIBw3PoyOCm8VA4XkP4r5H9DtstpVCiVUkkMMUK9QHa31+6BAXa4FXMP/KS4jDpqy8
nmWzjCzyw7qXzJ2sFbx+uGUuOjWmawEX22z2lrqoCE4deF84B3Vf5/5+lHrEgRUfRErlDT/DwCNN
VPbURGI81Ny4aBDtW1dBFyEefrFM5LpZWWsvKkLW1RZDua8J3C8pntRu0PPEg3ESqWfRIDmJZLfA
VZ8A6ay73fnl/XS01GnvDRTfKDyf0DKSFIRnGivYUEXuWV61G/opZMwLXvh8hWz67cz3cigGJsbK
Zl7fjw63aN/EyxmdvpR6kUoiy0tETnZBOM+qbGTl2I9fkH3NSLoRBk8mO3xCj3gfNAwSDi0mFrL1
h+rQ3mj/P3E9nwDH4Afgi3mItr7oMLGwbYFe8/+VmQf8B7RYVYxBSxK6yxEhXHORBB0o7WQ/b47g
GoSqni2mmBLi72mDAZELgw9OtWKLp8Ar8Iy1u+Z36AzYSn31oIhv2Kqjkj2Ax3VfW6ps7o3PmZmO
aQ5EYRGj4hCmm/YD+W3E1ZepLvLMHhgxR7qLliMwO5kv/vafXtGZ5sqFV5HBh1HsMl/Kx1/Oi8wW
5wbA+lbRDwgmGkwmib31QITlN6Vv/O1F18WfxRwQvGwRT+1S/VSEw+GMFKk22BL5anfe4DNvEkvS
LsDDUoj7vbqhUEPb+4gpidKG3E/0uG+lvo6N1jAmmwmiAO2Pm0ucngMDlSkpqa/gZZZfNr17x0bp
muzy+LUAA5XwAXYdvt3Z1EJnc9oaPILpAGzz3EG8dmbbVp68o4sTm2HaGGuiUj8C9qczIy+2Rr54
s9IAQN27pOLRDBnOWr1T0XZIHZ8n1HrbLyTSe9rBZAcBlVPwDYnOgXYiK7gqVh3HGOiJzPlpJkn/
utDuDPLCRSRfq2FxPLlzCJk+4QyMDdmGNyWMHud2y8mrZNueBZD4Sj+VY8Z5jXNF/K1zvSGQzUWB
NjHeqlNZ0XNTd6vM85quHFI3P2w8o8ZSwVtRl5Dah81hS96EYSMpU0V3kBPdJtTe/ObMGPOScIr9
a892HIvJeYwo09xCxxHDVuCnsBn1uOBWK/lgkY/6W/r3AOqlL9mhojWlvWbxUEMQr4YFcGmR/GRA
G6tV7VKcH0HRQXH+vNvUOGbK73Kw3relz5/Ox6cIG4hy1DfUTJNEt/SSD35mpXTPYroYC/YEIPJ4
+1TfjiN8yFbr/Ko91phVQresyeS5RS3DQ8GjJRv1MRBzk9/airXgYWg6swnwLFiazMEdhGJz/uC9
QnZ21jMVnYc5VPI/dtx5iEt/YyPmAky7QhR1ZQoy/s0Mulkonzei3m96+UEMzua2jUCfOe/Mcpfv
dqCXtk6No54RpLbktRLOCvSdZpoiOL9O9M6YLucEA65vSvojNjQojJE5Ter4FYBJQjWD5YMkMxTU
LmvCC18SvUqRFbQydHM7NtQ+0MlY1APfVr8D7Zinvy+AGNGlM6HTDjzWOZkfkik4Vov+OhZSLchh
HRNpIatz2jNqG+iANpfcOPIU13pWM4bn+H07zQEJEkfzV1IHZJ9m70cXc7HXxUWMBzPcVMaENmnL
YAE0OemQqZGhy//A3rM+U+90cISyf/Upfy/UD+1HVCEEjIWrJiwLeTwr+85hBDmHNv9Qv06iBs/O
yQkftU6S4AHhetUUfhJcUQQqE73k3ujqFcBmqNAvCMnCkLMdKktwCqMbbIYxbYN8qDQ7X+p1CNmI
kAjZ8NE6ZIdFBXOHcE5aj9eML4LaTnQbGPVqMT9yTK47jZnuelk/trY17thCxQQYPGof4yvQ1erM
TjFUFYiJkwwP7Pqh7lkm+SjYP2b5KOJITbvossaQmBi0G2MGdrjKef90KnNRWHleh4CsMnfwGnqP
sf5hr7oFi1GpEEK+PBSY3q8rC/Dgh9SM8/fs2cjis0Doonye4JweQ6pNuvcjVJ2x7x8PobmawIWL
tnuafiQ41nFrfx16jy8X2N6p8PyMpnUM5yRqjxmi0ZpK/n9RbzfvV9m8TyO0G9nfCVhB6MSBljX3
JqISeYBAg4/dgmSwusSIHEcoTLKRttXs2+yG7RQJ2MfM6DSSKxXaHl4uwYolEi1GA4NfgIuD414I
4ZuB+bJGr/FKc4CHIKY9Z82PEH/IaaUk8y2AXDlSo6YWahclCfFz44nYA3dwZ4VhdBBy1bqDTOBb
pO5zo+bLxmDtHvKWmpqjEMk7vFeoikUk1ScP38r/XyWwOTutnF+gWAQM3qBhijP5XltuIvQJ0mq8
XrnrzZiFEo1MBq3ZRdF4iws9X0kPzdWkqiKEmVXOPx9p7z6O7inhOh3OBJT1cM5ijYH6Tluh+/FT
qQKWcDriwPDrE/FauSODJw+mvDrkcD6YLTe2ytIZbozAoEnH+2bxZJYyy4MxWjFp8p+wpg7LV+Vj
g8h5FGxvRdJ1Cv6jS9UeJktmw6uX6E8cmLB2AV7NGigKsr5rb4ksWuV2B5+avJ2O9qu8clpPIXHO
IMuGAuCHrAlyOL6NOvAKQsyp81AAjkThICPxIae6H5TfITSMYUhpIxoZoIlM6Smbp1rFywOq3gu1
IAH9K9049hyg+m3JnBNwgDCZ+Ft1Q5NbmCRyIWf3ldxvMFm1OhjWVm0kc64FscEj+Ucnveaxg94G
XeR3TCvUo3yowAmhfRmcUGmpRv848ahhCpQcsJHcHTdbWI94WGaX1kR6VchDo81a0suD5u+lv09m
4aDV+C9cCGMahaxTVmnHjADlh8z1tbEEb3QXAwJtVho9U56qCJEftI/HhUMgFhIC+33UCWVd2a+r
T/akamR15KaB3X4Tlbj/IcI0eUb3/IVNFMyOki5eaH8qW4/O40Ggm9650uAYbCmtw88bh2U0L+va
ItuoVgubWLwA3MRKCR6DfT329rPYU3GWx/NWkRxEeW72BpwkasNfyIcMh18O++WobX0zAe8Lu61R
/PFVNzz967giBMCJy4+8DJoc2u0USyvCHEW81M9j+iBcEXUnyRbhbNf1RE5vTxoFt3u3NtCcsHbX
VWV4XokgoUll1yrOTwAFz+R96eMb8aOGkW0OAXCtc/dmaB17LR63cUhUXOWaf/eLEqkUm8di7jqJ
OHQEN7y8IkMZpVz0MgVaxFSTzN8t2bl4GeMf5a5NoJYE8IwgDoKoW4XuafXuNDY4ZiRfEpGmCcx4
RYR+Fmr66RvDkqBey7oenhLV/LusPpfhD35IeOFjXqXTu9Xz6D0l03L4xu0ik4YC5fJFvASppE0o
0zk9AUWUyk3HhOH1VMWf0CNdhhdpF4O+N9XUJyt0IJ2zdr2nSgbvuMuiTVPI3TGGk94D0EsO0Fmp
w5iEBEduWrOth30FxE1HfCgaZHkCc7Dwy1hPkxxkbxrztPmFiQ83wuXcuNpYK/TRTwOc/uxviQiV
mnl2kgzeu4sBvDzYwh5zOBNtuPY5xIsgJ7exD/Q3nZqJqJ4t69djdI7MCJpO/8HFYED/792dbM0M
XNHW+xcOWZkWUIcaQGbwlJuKYTlKGS7cgW3dhXJKzEGr64RIX2qVLUIilSl6V/CZLQMyYuA0Q0oT
TWjOLLLxR7/SJtMoCrIOeqzwp/uE+dLS7Wnwg1VAWF8DoaZsbM4SbqPi33fAIPF704P/1sR2yohx
AGugwAN0IPrFZaqyfWKJF93ygwa0wqpYdO+XSszsYIFfiq7DxeP1OQxNX9ALQp+/8p8teBYTvmQQ
qEkQUAbL1fNmhfEc/riy6Q+UZbP99jfNOU3MrZk7Daa2wqvaRn8HmvatlOnbTRrPRj/9YGrgOD5o
xsWpDDa0JTfxvLzJZqd+gDGvQnBRxxVN7Yl3CmSn5WkRZF9avvwz6MLBEBTCdTqO7WbARXJF4cqD
AjkDj4wJtyMEDeWB3iOUZit2vk5RTONu6FuAuLrsQr7Dc2oNtZu+fLNwXO7D5Ib+mISPveX34e8s
Y7PA4MysY3Lb2WVg5c9geCIp6hXX5/PP5j/pKNNZ/mCjMuXXB1a8Z6VZ0ejN02/0OdA/jtQ61RdQ
kEuGwHh/tKxQ9C82IOf5LT9yrvWxMs4GaXbfgqSxXLbdejBOyYlnXNkXB+PjqhZstdT7FTWfKU6y
x/jm1qgm+/tbuJiRxmh6iDJ3yvZB7C9eG0+g2g0nfjVOJAmTXXZRmgJAEVo5VBOnJdU2h05fHJFz
UkobX5WR1qkhNOQHEQWUf9xmMp76u5NPxzayEYmyc87a/zeUlhw+gSWEsflQfpnowxnSUXgftr+q
2YMDcG+R2PHWdMx3+1+WLAb4pP3+FBdneD+ZA7v3YunWg6w08GycJjWgP2mX7TR30gi8LWGy0HTU
g4QDPLyZfrV7ibN3sTMVkHUYeGAc7qvedZxNJN9tnpJmHGEc3IbeWQK5V9PK3JFNyTZPbx2V/v0H
Q5DLdIoFISaNZmsaC5r2b46W8IUShMO1qKhyyfsECxvrZRnw3pbe7THexb1XIEN2mPizPNl7tkYG
7tNR+OFrYkkVXyJNfTr5Zi0jZMXM/8wcKpsZlDl4F77P274muKpt0Hkmu6cFqaG0gwWD0pvZaK7j
yswM7ZE6NeLF1fFPRbrkyU2oeMWBtEmyP5QmUWYLzFIwXeWq+cfhGsUED3rGYyTChTIyqDYgll/T
yWTXbpsPbg+OF+0as+NNrebJh1HkidlgeeiDKuvzYsOHCPaiVJQTxYqZ21HVJQiIjtaGZa/2C1fG
HaoGnWDNXpxXjsPKzE5FjHFA8YSaZPbKIXnNBp5F5Tx4cMs7XfSqFD3//7PXgwLFPtfthlSV8u8i
0PHqI7nZiC6MXHRw9WNbD/u4CEsSuVvsCN1wS08uUnGTA5ji0K7OnufYnRikOdK8virSSzbzAb/a
ojQGO7XNjp9gUMibajy+iTOELkPs/6uZHHyBfD72axmB/KYoeTu60Vim0Q8eZL4ppzVvGH99UG8I
aQ4NoxXYaE9ZPM7tqndo81PW9SD2doZG10m/upY+z6wZzXJzyw7vOIsN6ZMvqIoO6Q1VuR+TgCHe
nRwyUZI/Nn3zUS3DWjvNPF4K3x+mvghXvfkO3SJOn3gtpWRV9ZRDSboGjKZ2WgdHk62bKFFExhoG
2FSUYrXE79mTPEokAC6wEkh4mzmTK9n4+/YLzlqOmJRESZoKoKoeAa6BIT17vtq+cUz+iiMwnVfI
jYPXCeth9b55oyty9tXgrHOR+AZ/1dA0qYFt8WHdP7YMLhixFaA6g7fGFuT1nNXA1tX8UzZS2OJO
3/QzF+YYR3SDTgEF8vj1qDfR4+WbPwciEGVe7u+8TnlqyZxzOJM3nbCPVvcfOkQmukTBSgNKduOu
Wi8X7az0U4sbPrSoq6+rf/XKG/nPNy9/1M3CC5vFAhxK7G55Op/hUXqc8zIMYUTsZ/e0QVQDz+Eq
mCLOJq4Y4CmYumkPW9wBFLnfEkB/+WbqEPBgFAglg4zykHfBhZf+3lXscIqAXAqcs0V8V25k6JGL
a+fd7yCqQmvX+pAjS/0TYl+/cPA+E+1wyIjF0ueJyJhAHtmaN4oYRapxxH9jonqMoOR3lvpzv3Hp
BIOmgCRUhN9Y6o1PNTOATioe7NGtkUKR6QNT20vHI/usMnRBKYyoQLhasFPdEkRVOapbXReEwHwH
0DczW/HSWuyl2ntIuGYDfvTGhJbKtHoShXclbQR340JBlgP1SbBKCGixzzzulMVgpA+u7o8d5fwz
oWHZYgTOV4yPDvsW3T6oVvRijwp3eht7TzHiHt48j28c/tOBRkxGuEjQDolVS06z3at74BdXYKmY
Ux8hO2u+BNRs+O9D1zdBmpHqPrSSYSG8a05P0LOmPT25QQc/PpfFUIMh2N1lUB7Sx1n/AQEduHuh
/ZYgMouBloQV4mlqK0vayaztdqI33uWWTa12W4U5RvGWotwMnzzby+6kYYDbyv5/lA/7nGXM8tpp
QolFQGM66iqajCalL78dFyPdUksL6Nu3fYz8PZVS64Rj3KiulW+EoFSBEzKGwSiJ/++JhtxA6LBJ
nZ/87MY8Y460KKG59QHpN5bXehJfNjp8C3u96ZU1d8G8hmhaApitYr316B0OwjuoWwxz97Z5SnFQ
woCgam1AhIajGfF0L9lGpTgV3uwApFobQA4VaS3W64b+sx/jqwQf/tBUT5p5yX8+bpDlgLkEVvCO
FS0ALFQtDqa2NofBS9fmDksOlycbUiMnOzsiMwUcoWRJd/68+YlfO9V8HSN6+2mOL6qBT/E30A4Y
M0Lo9otGoi4SrPdl/zLEMA3pK8yYrnWBSAAQXyiIVrQz8XASkhbn90RRNovvtis4u/fziEathIFy
cX+9SFiQjctxs3YEzD333qUIfdB/jzDGO+mxhTvBVuUmp2WqrZqNE9hlpkXc2qAc5P68T73s5lNy
gJCJPapwCDaOvsLwMjq0ZdG+jU+8FnEPzSr3afuybh6pjpN1HsSqYqJP0ZzNTUHaz/h1QLAIWRa6
0b/0r+3LiJis0tXMKRdt5ObgKckhd2L2G+kdmI2daHehajWfHg62QjAbX+z4hFa/3YF8iuX0FH1N
eV3e9+OOpBLb0/KSuBJxjWZ+qSuQ7Awm0HdD6UZ6Gza4w8vELV7cxKy5tLv06I4jhbljsOMTuSue
w+icdAgR+EWQCwKjlYTO+gBCxeRioIIlR0Hb5SQPXY1wkJnFgp+a7yZ6wZzF6P2vVOScjQgWrOAR
BSDt5h0r30JpCTuwt7AP+39FZ08nNAHDROZvRoiCakAXnbOqZc8OhGT6tXqpA35QRbM2AJMSEZWo
7U/N/kvJ92EqreMNFO7Ok5ME8kajrEx6FERE/FO7NLt+tsJ6LbLDmpIBDaJAYiE3Enxj7o63Zvsl
wzZ7V9pCjndoGUkeukBA4w1b6D1nWWpm5aRWRswsRBNy0v3UXNKvHND9tYWOIUXqVKtHa/l8UQc9
8TppYB8IV/tbDbXlde8be//f80B5DVlk5vuUdeYBLzO2qJGOriclIuZbBSVfn00wPgY+TQK8Vnjr
WnvyFho5lDDVJilUQavP0swACQrw1p8ntcT9SBCsrrwI/+wzWaBIe3bowLeqvkckcYPNfzDsq6B+
G9m6fCqlohunr7H4AutF/a4zdmP52SWC9L7Uc84YMzt7ZAa6kWt1kbDytP4LM/+T1PbiupNly3rW
87XfOJ/5dACdi//74sgoiD03yv/cg8X6rwsfOUoA8bQDwQ7uSb6K20LBO2wxFsPiF8ycicvv2Ofw
kWBZ561/UOCdtmoU+rcdQh1cETdlrzm8iutg/U67rWXuHBK3xaGWKOUB+nvc66KjjHXKCuLog/uu
9JrJ+qI1GkOPW7j0f3/Re2+qNchntmitjE3lN2x9dQeQdTncxMBKCpm3L1kGfJy0XZ2NMjNK0pjE
5kppGZOjsk9ar1+vSGdUH+z+y4L2mYs4gkGbT7AJDxJtbEzbzFi+yiVGtQMYD4jsGuuxBsxhl2Wh
fdpREWvRRwO9KJmo5zA/u2v/asqfcd7+LQuaKoyrXgB0BIV5YHkG1utQItNXHzaQN/QyssixTR+m
ckP9hRVmsYEWkQ4rzXEVbSfEJm8/zMXw4gw12XovvzVwB+MAU2cwotRz80xgl/R/fY38dtBaTXjA
9fGuRf5prvjuuK7YfyQn/KXUce7a+wDlxHguu5JC2jWY7CLyu9fwHiCeKSYorwg41+vNJ+joHU1j
Fi5ANTmaQHvmmbGlk96lhbRTat8K2kSvua97hkxsqXadcGDJ6aRsB77zwFDDaZb0ySLTHvwruaA8
SPtfWQu+Ue84/w0uTPEOqyoQ4eM8Svpy8yGzoQuXZXLUXKLTri3WG4Ym2vWFvrmj+EGg+wArVI28
6RqPRHN9mBNCA1EE/qie2QJEbtYEGQwarBVwcdzU0Kmp5MkEbKxmw7Oy3t4ejjsDgy8nm6a7izH9
Ov+68TaCTQzzeNUGpCd9t30Cjq3sjjjkA6P67WFOLKU5MoDQONgIk8amOy4cWd05Xsj/URb3PJKA
EUbilKWE1TYfNh3Py19kE6LvEEclBHZ/glda2pgKwp61c669MbikZliQStK4jnMOvNiq/4/cqhp4
T5VE6XPgxFxmdWlQngWF4a/zU1a+pSQhnhJzzUSVQdFA+eP/4zcbgW5XvW92gZcX+zFyAyWUi7vh
EkRflpRbYsGWm0k+aCreV5sl97GdHluFRwL3q+m3htC8Hs8iEUFT7ydEM7JCQdeJcNjlKBykCbd5
RySOYYOJ2YM3CJUhTHtlXhRBNCuyFgz0VYeRZLBhFZ6E4VvD85mTOl4+d4cWJstYbIY99sp0qniY
tYikwnB+pxTZRebbwNfPrRsHiB8PVCFVMXDkVBtsPZ0BglUJSaRl+qNY15n3dvwH2w9BAIaVKybP
NVuWiaZzzhSJXBwv7Byd51nRzbbLxXGMVgeyxK0yx8p7hKH4DeNbPv7R7Kp7jM4GceSBe+DQe60G
5lNdMOif+FbrdMuSsI6msDR2f2v4nQEEqNtY5RaHoxWZ+X/q44SDrZb5syYF5ph56R90Wow7iJAT
iwz65938oBOAGEGDK7HVAhJUGOMIuu1knv74Xi7GgS320wTIPdjB00ksx1JfQZra4fO0kNtxpWaZ
jjnBFYxX1rpOm+e8ZSCp0MuEavud3rp3pCyTBPrZNwk9RTY3IKUlf/T17I3+UKPe8L/mTRkYiUGu
Nr+Cr1cCBEGm17FQflgjZczWbV4QKuZZaMla8aFYTQ1rxWg3nnTVIXTtsn7Sf1GVqk0w/OjUiEoh
DSu4DLEKPGoaZjKcWzzr2h76yXdMA5d4ZJcVbeFLbva5R4TPR22NH4viC3v/2nBdkv7vh/mGg1xB
NTWOzSTNh6FDPYLDVvlnp6UeURMsuKR9ejUtF/6RckLE/a0PUJdMno49VVXIJUPqsb7YBlcIQwUf
yy1arJhTaVSN+7ZoRzFVOathoZcsyEmqXA2yWhSZI5Yek7Tf2uholDoEj/WDizOhm4v3thaZUxIx
CxB28ZWs2L1VCOitsVXDnKiTUds74AqgMA/KiqDCeaDK5R2kKRRvi7k+j5GrNHHnoQWS4y8ULEvU
IWc+rosMNNRC30wrbe7psD283wVosd2EtsCsYGZ3VYanCvipu5Q+sqfjUYbGvO7wlpYDGLXpRLAo
RUMnJU9KpKVCv4brPzoIhiyagyW5GZiGxdgKwht7EWMgK8j9joAj4XhaIWPK8O1K5SaGeTvOrGsY
2vv3PXHnPd0/p0zhG6e0B44IqPMUSmVJtqA5zX5g0crHx5YxL7sw9xku3n1BfEn4kphhCQKuRycV
gz7079v35ISTEXMxBWxZgoGF8d+yJtNN+Zwm0MM6kmhgAg2gas4TYcR+U1oDaolyYdopsyXLzhZp
dxfK9GU+jsudajXOtbf3sUqkv5rGN46lVdf7almap6cDRbn5UUIy0ya9MElGB4AxaWMx1nptpvi6
tXj0E7dIYFyg8KXlqYMlhTRC9y6QXxNPwDIYOGX98sHldKQ+ZV6b+UtMJu9MOldZnDcQug6dugH2
Z7BRwYn9VAF2zdogvYHKov5seBXpgjbaseuKrZLy90P9BABh+C1dZ32XR/7A5XXdvFNW/LkHlAwi
nG7Lwb/dI52QQNGue5VlVjQ8wNBP/glUbVEi44lYzqS/WDAK/gkBDhR4rjfJdk5HyyQVuSDcWaNN
jl6PCDjuRviDNws9wXDZjrji4NE4/tEMOjWWo1NrKck9Z3EXtXr4DUnBFRZRK5Qgr8yPFPjrXksv
xp6SAdDg5B2wO/BYjv0HlpvvlB8YSJvZ/vzlTgagB0O8JlsGvChAOVr7VJwTXpnjrBQ+1qqkAYmM
A+N6sEdtZcHYTFkCpYeGgiOUI/w9PMCx363KJ4hkqqf+sGqmSCU19mMg/v+TeqMlMcVYTjUiPjL+
dnYlLOYc2y88EI4Ti83Vq8IF/uu2GywTxDK/YVx72Qu8EYCsXxwfJ8wyGliSvwaPB269PjqCidlH
rN9B96wxF0t07cyzT2ite2pJPE8sIv9K+t+5QfHxkcd4gYSsVKEqoWlHngEUWnQXLJp6K8wI/61s
mzQ5VaNjWyLKXxHL6ZJFiys6sMyFYJ5WW9q1CQ++22oADeQquGxzYwHucm5qkpJfwipSz6Dcb5Cd
9trIyW1dvcjr1cRLjz/xzi/RPw2ZmuyCWSAQLljM+7WnlcSK9NnTkCKHjGsjw7k/nAYD4zs0Hh/V
U78pPYr2qSBJMjRmfnRw2x6nx2bGiHPNwV9OhupD9B//J3wz6gvlg8rVi4u6Zj/BU3/sehGYjo9T
5B7QCUmUI1p+cl3zvCtoZx+xoxRnE0YRNZnHpyohQquTsCNHBfDgtU2zS2LZ8M2IQRL+pnLc3hLE
w0MGnoIazumwbhqFrD8D1YyC2JFHi01K0Oxf+4VGDcQojT1rl0/XlP2ukTzygnyguFyFu7wo91WO
x2N0Q0zsqLwxLDnf18Dn/VG9yXtE10TGUURX3eO0G19EuYSfhQGbKJ+VLPdXZyfHPLawHKnP6mGf
FQVUDK4dBXrIxtXT4e2/AcbYOiv6O6tXIvTar1w+6P9Q0sRubSNyU89quO7+ysdHP+c9ri53/MXs
Zj7YM4L3LNLp4F1GDvIQROmRN4D2/Ex53jMRe1HZtsPWZxySUgD6PZZ38edCdgQiAamR8BEpfaRa
6rqEJUXECt97V0Y1NXH36AyU9n9Pk1tIS1kUi4g+6RHoBT4bFYgSrkh282doF2g9jF8I7qshjiUe
Gx8wzaR3/cerl0uvGSxnCza+m/Jiz9/ou0SUl45m0Xk+U0BrYB2iUO/VRIgY8SuOkdhpKPDHI16k
A8fk78GRBk0LCsXdg7hk4E/j2OxRewwjieOjdKKqleRRKptkygBGqwJ1qKXfEw8rxTHsZoQkhI1q
0X3iNLYf5DVLm5KPc1lt6mu7PqHQXT6JsYYPC9WOS3KQ97OGaMGlEQo3YWBF/s80FezY2riciTa9
oN3ljY5z5XNRZSgaetGu/zkiFEVVQLWLuxr2E9rEd4XjnbK18lOiE5HyvNI/QLzrq96LOfgXsU1q
dY/RSFSECLnBgSQYhJiIZIKULiow9eXxcPRsaykEQycwxXRjGCimhLkc3FdK8wn2QjsuMN9qGPJi
VHtkn3xle3aUWg6nvjR42lhMzp05WDs/o9HDk/RKjp3FxtHqW53SK3xuuUvPWiuWSlYyQQy0mMM7
TRg+rUh+yfAvXAy5r5gRObfaamsZjX46pthAWTevLgnLr5Ri4nqFG0lwytzlg7RecPKdBG5+hVWW
yzni3zwtuaTiCPqAE4hjTWIgRy7VPp2F9gbkpm5NA+enaIdlhwIKd/ACkuBhYmrO/nnSB2MnMGlX
aIrRVl+cr8SKkQcpOBubARKJ5eojKOmJW+A9UOqx0H8KZs1KfeulMIlqoFcvZmYCFAxwBmS10+LI
iiigi6ThMbtFeGJsj32WwMZuCiGNX3/Yozh/CTy/8qVT1nmxd3OjvVZXPQQHX/g4LVeFC6IU7jox
lXQyXb5vnxysVRB1wEF6ABOQCBYz/tNFej8mEJ5vW/E11ABGEyKbdJZy/rkAZGIf6ULtbC9UZk3H
ojEia6DDvSyxTzFOVqJrKZNu6xOgXw/2WVzuSbiGCxJznbGg0ZpI7MARRz4rABC9thcfA4D838rY
oz3DeKNSVfazZbIVOOAbExyLOlNoStgWsxjcBiNQfcWD4N9RzujOGmuoa+7FYuSlMUL2iG0iBXMr
H4jl7IsYIii/T1wnVVaaKNdtrXm3ZvPy9Ir2L6LOZHnW8KxVIrJ2GDKUVANzZazeu9P9QF7ASbP0
d8sLW3ajsHgNNoEPjWvEF/oMt/HZxJnVzipjbpWBn4L8RrEOfTWXobcA2qhQlWFzxWdIZ4cc+VSb
g42Oew6hfjAz4v1zabY0HXO36PjCb3W778IhiUAVzjsQ0kwohydX5Ylq286YrZPNjl30KohGAVIJ
+26jZmNl3m0kWIMHh+e/874OTCsCN8VhhnyuoVhXgHUreKH4DtSt2VyPoWLLHhqjHyGJoT+91qRG
TKHwFKVgYB0umN7cHdQwyxQ+cE04L15K02lPxt9AtqUNaZaYEPntaManWANKKMbRc2DIg5Pc1CYq
2xImOuejTrnme7VyR8MQkWykZ/IFOJYgNI1t1GLlNfIUiRyi5qpkw6fEIx0eXg12mLXVtjztMX3v
ehTptZHx/+ollXwQE+AnAsX+q5teKEYlIKgHP2hnihzHFfGhSABENFTS/ESKC8KFG9aim5yHmHlc
8vUpfefBs/ZW7QqjQjsuk3vVauj4OZKvR2g1FIPXB3zKwK/qJnWZdtzM/XeckqfGKsfCTsKP81GJ
GqO1srnVMY4HNqlcQJe+tUJsKntMdhvUEH8ghZ/mBbq5tGymxf8/t6aHk8dt1tavN8bS6EBBTy0c
jdK/qUI+KlfNvyWf80t2ZsAD6owvBEx0fAiJwDwKd2f8hIklzfdq4DdQQjauTCNO8aubvxIwv1ow
WMqOuJYyhe/utanXVIF3iVB8LOW588+4mug6GUr+HJZ4KZXi89QtP5Daq5isYia/KGnEsUeCtidp
WgG68VjLe8MjrZjamFy5GM5lU6YbDu91be7l1Jl1YHIw8cFpUThne8GCjFWkVQDHhisMSwpj6z9g
R73aeHCCiJbLQBJ9oiry9az9OOcqasgcxZedAfPS3djqBsoHN8OFgbOxGa2InLh7ZauXCvync6el
sZCrAGXEnzWWQx+6/6JNK8iQNoV95zo5DzGX7HtkdeXgS/22+kuiUjvxLvZcJz5jhivPkeT9J+L0
glA+gpqsVquOZbqlB3NYaUpk0or1hK8mWv7dRUJ0HBD1yjEPNgzTV4A+hI4XPEC8m8xXlwzgdVwc
+8ul7cBkU58woWsaEGRi6+2vuQD7b/SI7+PBo9ANVZJ4m+5sss8KaBBdlSUJ6KBShrgjdUkK2zyG
m/zQuqT1blUa31xr6M2VTjCi6oFkEbPbnEMrnDpV7sOzGIfBXtQ/ozdDQNqnNSxlTbonpz9ORPUH
8pMCJdrJ7q35AtS/LiBhdUPgudLlbUbdIpfSk6pgFyPAwp5dt8gyjS4EWbGSQYDCY76hUPGTkvQb
8u/gnnljyaMmFxb2eOQSr1+oSWxFQJCVKJeUQ/J3PxC/570zdNei8GTKEeMrtbLAsO/UlFrL9vCH
U+L6ePMUO3IaHTkbDNJcgJVw+gzBvjOQQUJtIUu6Ugb+HuimmLJHTlX5cvdel4hM7QWxvCsCQP8l
Xh+scZt6jolkg8NGgZ6KW9GqTB1KK1ZzRGk3+DqVoIvWY0otMsFuLkEnyE5ia4p4q0NM5WjFdoot
RUhMbY7o+E6ANu6MJB68g6pf6U/n/D4PF19Tl+rDTNzE91ZHLYePIAmOf2Z6B3voYu18vJEwdz/p
h7nPmKrBwVd0Gs5uUZCPsOsh3JdMlyoOAamMt+QHj2BA+YZHKqLLSCGi0YaWmUVH7ddd2nYyt8ni
gIyMfbvr4e1X4GVEp9I9zeLm8aFgbMrBjIM/X5u+7Wq0q3w0DxLJ9uWJNEzwnQ56GjTPkLRWuQZS
1t34sVov2aKbfarmBQkhls18/EAHYziag/OaaRepuRF/0WOm0zUPBG7G6r/ZXW+BnEoIzfREjjJ8
yaCqToPvmq8k/VisIPnbgOMgieV+osPPpx/FwK0Dx87Akkojy2Y2ffv32OBIDPvy4G8SXcB8jQ3h
Imsiw4kCE0JAxsmAS9uWKjDESWhnL+DD/HGUncpedR7LaZVVXKaKFf+Nh/T0aB3N8yequJSenFTE
d5wVm+9yO+1Eg/oFThucoVZMds0KB0Iz7JDXOB9TMMt9UXHYaY4Fvaagl00j1cKQ0DMYZo1HyNw1
iORDbA8fILneh4GMJym1RWpce0DAK1cZ9O47pY8VGZ9HGhvv2idrTts/LJyKhcTHvL3MLXQOm6pL
81oEahYgCBq5l087JHf4E/4l4YckAUqMOMjix0sNZvPOlbzurRFSaJT9/2GQPOAFlzanAWT71kye
D+pmMIZbZEwG6n7aJtbc0yQ2SbqxEHH80EUY6dcx8524FTkz0bd1WeAIzUG/TqWJQZAsXaLXIWvn
91XsFR+8i9af9sTiGwVBnR7AxHOXqWwF+nhzTE4P8BxFZCpK7QY3rkWj0A/J2hMsW3X7j+qL0Fsc
GOYdwlWBmixp/FbMQLu0853r9lDxu+zHMMNDjtmKWj59eavbDPN6pz3azHpx78IUdTYxOSEwIvL6
mH5V61tm2bHM1/6bKazSc/xvDOBI5Recclj/4Y6IqVWn2Sb8K8LIiuih3v2lXtq/1fZJXBhST2w8
u3gmtZSw+B7iurjX7riW357vwVTGs+q3VxrbD2fR7awPD+0Gs8TGwJClCvACVRYttUSC1bFqSVuA
edrTIxs9hcTrLHHdFX7Os3wpfqBisH3dQxCf+R26YRVBps908XrCxrh85uJSosG3ezNHM6jAsdyN
Bn2NEUTfwfsd4fzAwrWEGEyce+x/jqFX1BA8dsm3Cnng1kq3xb8tDOskNcanNNqTSKI7nQS7WXUp
IGAHu52fLOlvhSI40Tv8Xc8/g3geiT4T+hC3ATwOWOAf6YkUn707+c8iCof8mPKJtn2gUW4hj/XX
G8P6w5wKoKp0AzKRmPpKi1PR7A7OATOoejZFhw9pe0UIpKVQrKvbSPULW3fQ8wcxlPxS7rfve2/K
2dbYc7KrPAEKFFDlf+yFK2UJeibNvm7TMACK2CYicu39IdDloVLQpdKvOTJuJMPGi4kc+3OzJhSF
kXZ+k1GxgHneGNkusXllYQ2MWzXInLg+CdSA+ZRnc7f3db/0HDOMhlQ6AsIjLoxHtCwkmfCuVNiO
1UzuBHrbSTuXEH+HGtLGR/dK3GF3AQwaosDto0BdMmTvFbUSHCUdrKZc3oxw3cyeZV7sgJtF2ILi
K8sR8mpluH83/aSZWIvQwjtw3QwRE5D4X/55PtpOs3H8njYMzdkf820H9Ayenp3s0kIaP7dSOYdv
p/Rlo0AfjmbXEcZYGCiHSGcv2RKelxJ8JyrpliwbWiRYCEMclJK9/1RwdZbJ9HFhvoJuDGxpZ0z4
xpsyWKWd1V2T2ZCJRGNYSn8U2+C3XwzzB9mmR/I4O75/CZQ/e/2z1YvT3Twzn0xM5YCSwhVpjNLG
nv8TFX9HNUMvxZrkb696jDAChU02JvbHi8E7UFmZGKP093fUWtJYfVKCMdss6JZoKfvENKd3rlZN
7PfxyoQahnr+UiK3RG5caNDc6nI6tyeM8VyqQoztI3TB7YmK/VNjDerSe6c/GhxAX0GMpKnKHqmY
mKjCyjXYl2LhdBZJ934u5kWqfQy7Z7s7wcME5IUZTqhS8ZUVpKe2oYC51AuUF0O2OMw4Y7mq3iuM
28VyGUy176BdBVBV71ayt80kRJnitz0YkjRz6uN0kR2wUv5pwu+s4KBwGqwBIAdSdZYw5vxWpQDY
BBj6qFLf77sXfnpmJL+IwBhspEjmPQfwPSil7dwvf2fklaPOAOkTcKirhQ3NCek+yhLSgidJiGx0
YC9UsIxhWwJ94PDU2msAb9YrLtZbRuBebufVf9yvXx7WDo0A8T88WFU23N9baeo54aq+ovO2ny/Y
fqkVwfm6SLW8NB+7T6DkHhYbXnAwQEzQ4GlMU2n790Znl7YuqYDroBGiz+qnqhEKwzY2xKDtOuDJ
1NEse7emcS0uqqCTcqD4xpcSA9D8X9yq363q/82ZfKpLdSDAqb5Gwd8ElqNKG+tSIYB7DGZEAjkQ
9J4o8EPXmRo1PUzrvh5vh3did+e3UpmwoevB2RBlrLWfkaEyjH6L6YHEXvtoFdUUPDpoFvo7A/At
xNNLLvqf7RHdVE5EkNMmvsfjyYvEXDluTLamo811tFNQcM4Bb3ZM2oSsasU8xEJu177NqHkr4bhw
K537zHU7+f34ub0YK/jWEiw9eOzzmDGAlYZaoyQtw6YK/LZBYr8AegmEQ62ZOOrfQtE4QpX/MAFE
1S3Raq0n7vRp5zzwH897hz+DY1+pNQgGnNDWyfjqnz1i07FNw5EhbRHsoa/8XBYi7VE/vTs/Z6wx
/AU6x/SvdxOVkCUptPgyZyiG6D4T3jUgzbiE4cYTWBQDMUK/DSaA/mLRy1YgbJ4U45/7GOGNsYV2
rRNkLoEVN1RHy7QFwGgpKlJ/9IeNohAxRjKUzr5IUdMJgzmaiVKftNiCq8XsCxzheI63YYya3bMc
oACJ6VqKohkRYeugqWsq725M7Y0iPGmWZRaFF5VFG0hvNZZNxig50ksWOyg6Znw9cTJ4M6p6J47U
079Vu9ArIfYGGTmtixvSVhS/1ed1Aqlg3GkKKCbMN6k1WdoWzpyfZWz5dus+e1D8cqoZinMrwe7X
jJ0tLz4XgBXDTfXoMTmAEbNL+8q07DaWhFgeFiSS+h4tWkqCpszTUc7+EgFAiC2//gQSC8AR4E6W
auOaz5CVWudhH9t955OFmVVZ2xTcJ1tdSpuP4YXPKsWpbCFTHKnytaF38PaX2IyFDAlt6jfmkh8B
k/kBY6p/BhjZ6f/UWXTxD0LmSv7zuy3H+en+fGtup79SB0RnJTPqvMH2/e+WlCV1cHRWZC8r6IDT
SyC8vp2MMCykWS/M6NxdaUMsIdwhm5BGrvE45B+uOSOwy/RBMxPoHNZAmjSYGyAptx6M8Kzd3XFF
l9SKzkgVmKSfGTXzk42qKTGtmItp1UlBIR0bQlC8d1Wke1KhdoE8eudxwuyzQGq7lOiZTUVrQifj
eZejhpS14gB794JzTDAsLnLQGqosjxRte8cm7JnCD1PSfFOzjawWg6UKam+nP3PSnsr2qX+jkUVI
6rAmcdtJ9izEgX8UurqpKYUXHjXASCaTPd6ygPpxw/Aoa8B/QlAf9H80Qx6Y01o3u+9mksLtz5oB
RmQ1QZxUWvD4U7svdktjYPAU/h/uGCvZJ+hBqwD1VgkEWj3Z4kIeFvFKryccjXHPfVq7RhllhkER
HHrcR6pnWLkzwITriJSRblcKABPVBEjc3cNQg06ZBPJeDQUg5FI8w/PhHynzSVYXb0ecpi7T4k5s
YyOc2BEG3dL7RJVP/uRSrwChx8oPsJbGdPauwBEnDwGL5ed70DbtKW5cLwKmApovOMsLzI0UKurh
FN4mQLEeO8Zctv7fyWgVSvXBBsaWdEhxjaY1o3jj3309tp/n+h0QKSbFdEGKmPywT/glP3cZY5Oj
F4f82fSeR8QilOHosOMRkpii++osc4NiKfwYuTOzgcBxbBoBAjfumAaRlY4+D9fsNWlDOFqLn0e8
oyi8nn44Ifa1vvetCa1V7pnP5seNwIF2Jb3Ab6/yMf+QlnwIoskPrhyA8N3pFlUCr5ZkHcPhH1zE
JRsAOIrYvbQSBWIU6f4jlD8/1LAoNq2mCWd7mWRC2N/elHMIDZYA+LZHwl4gbWvZknIw1pWVXzPx
O+wa/Orcp02PBhU88oI6wpQ62CFUj0Emwcyhu9LsI2mLYGDheZ8tgpEwwTCQI4dsDwIPWjp8P16V
fKsGzH9EHDDChbMWq/Oz0uMmacivBwtjS3Ep6FoYjNJcpooUpfuOx2lw9piSyZ9UtJSBVU/KeRVk
J97+JyGIbza15tfHeuzrf0SHGJ2FByGeGPljAe4K2KBF+5dJ7N5n/puGfX3ut6jE0NNzGu6DX86o
YzVrHfeI6LG3/PILLcnEAb8LEtMOzkwAZSRIt4TSlppWkcsAoQfD0hnNfFjyC0X6dUcdiwZTX203
pQZ8nemGfLTKr7xPFZOn5Z31jruHYdD7PE4tZx825GalOVWD4OIhcwiADPOJ6sNVNg778Kq4cNK7
UmpOPzMw5iPdiG7UqkgZpB4v7P6U9avznihsEShgEUdbMXzpBqj3dySJJL4ilQRreKdbVdv903CW
uQCggrf1dSccABobWkvFcg9HHrI9CxjFpu/HXV89xNRQeengUF4n5eNuMzlvuNnN3e/JCpFil6di
XPCiA//7aWypxmllboo4xYsgkb+XWcgKD6PjAwFJztpBAnBSBz3kTwcCDpYeAHFOhnfkXfGWP79m
6B8WbDhS7ffUOABNxlcZfYPPKCRAgEhWY8XBtPTyniWKCeqjnT0L+CBE/2hzjMnXs/ydXW0mpz9C
AQ+ZnFvsINkR7CvbQN90IKUab2ClmkqAJeqRLSS/FyM4SUdr9Vm/Q9itcq/z3Zz/n4gYxL4bRAjz
8hFNM2YG3lbpoV/10tDJnPSnAIutLIiZcNFDxlLiBoSLRZ3Pa/i3H4xgQIVyvtnKsC9xK2DGNBL7
odawtG1fqRQEy1b+8B7W4ppHIgT8D+JKC3r5tHzxlVfWxh8XvO3trV6x+WmzsP/fE63WCCv+RhGs
RvVhSnI9JKmFscZqHQkeRtJXnqhAndMsb5p+5uz/UEYNcn1LG5U8LVgAVdL7gbH+jNpwcLsmdtiZ
X62m66VxsGAkCNMzRFcOnbrSZwGR0iK30xriDdXDWy/acZssfNXQ0CPaQhkTbwBTP88MBO/MBxoq
NCCsYGFySZuEw/KDtotU6u5nQUZ8Flt24noOAB2pQ+u09JQNTdIhVf9WUke+Ut3KSx6eISS4z8mX
uK9psOr8kfX1VdVOub4SlYoO+9HMpHJ8ZpinX/2B80pEEFP/SKuP4u8j3lNxTli/vdyn2Hw/FpSx
jZLKEmM68mm+Q7UZcKumS0dVZulguai7So5STBEMp3zXfoiKHD4Z1yNQolWaTbrlPe/CWnu8YJ8j
0kWRt5gRvGe0MP+OIb7s6pS9zwqmKDnM92HUF3odpSZVtYGTLjbGNuxwUwwEoyLF6J0sNtjpehrr
SjJrLAB6cnXB4XUnXNqUDnD5oPfqaUExl7lhs2Y0h2139Kp8OdUBIKQsbHvCGPS/McvZGWNrpXXu
FZ1iZsFZRPAfqRuz5YkeA9v+/Iv8L7WLsqfCJm/zCjCIb5+Xnvk8AAqjlfvQlWcq8HrUppq+R4xJ
ucyllvYKe6mKTk96UJQrRlnBcy53/EO/Fz/5Ul1pJnZoCynSuc/z12BAiUvXPhrp9ZFTDboQCCuW
ZfWfiCYyiqj939Oq08AO8RxaRBUSnm+VB/KOC8DSpQmabHDmtC2ORJ9kuLQ6X56Z0sxyfTl9PvGW
5aYrmNpO4Ol/hmFx8LSf4yXSg7115kS+CIZ9d+P8u6tVWDqo1OGaQNweSOF15rtUA7Wm8fCANFF+
pqdXDatKPWDkgjtErfAqnw8muoV12nI2wb2Q5XoNDCuQ41knPbhn2m7FBgI0/BZZlP4UuSHjO2e3
DCdZkYFQtwfpRphcjC/FmH3OuyQD8ajcakM6WJhHlI6ka1a2jNo+b3dzyA42V/Oxo4fXbIUEcskR
CSRvfwGpRujEkotAOpaVgjaWqzVeO9q7NA2EgFFwetQfVdLRTaFaBpjahAZ8vng+Fvi1lAH7bQED
klN3XjHTudvozvwEpqvMzF+EjtiGrOrr/h6dGsw1/HYI5g7N2jxT0KyAwdeYurLA63b13RlWmauC
y8CIpkdfAelhMXLH9UNhMHu5hfK/dKXE6tF6ub5mH9SKpU/dzolS0NikVSG6Yp1CGMv0flNV084w
2EUnFTgdMC8ERVgi15sRkxvSx3I8ITvigDWLi7eP620ackntPYMobWXhayz5OGlcqjBe0732Apcz
PejvSZKv7XkbGt2r6ZXERNzQCJm3IlwxOwiZJu0tcph4lt24w9ghUB2zp6RH1hwmKpaUzxzKXK5e
3sZithyL7KQbMYTMyVij5MS0x8pYlV2OKFRdL6+m5iX2fMZ3QfetXR0o+DLltCvYm9e8eT6uWDyn
/TOml0F9lwaGi0lxGz/JGQUkG6fqgBfFliB6iiDNSSKSh0Hc506lgFV4nFkdilaqx/WVc0NB4JXl
DPGnH0AUbAA2b2LWRXuuWtt+JUhnGxxShRTaglNQDBWF42uBYI1HakPOnVTSABjqdpJNeY/fcAXp
RveiPyG89XX+3++VA7xk8kgZrq7wPZX8FKSecNzote6JMRso+UOTkZip7oUhpNRxE6Xp37f60AK7
dmxyR2RzbNExdufI8a/XWBoyyb84gcN8I+3KkD/DcQWx6oHzEJ8AM5bsaFweW9X5siJ6X+AGZ8F3
T/U8K+qoJE+EHf0T6eTaBj9FPqDTfdKM0BzmKC0C7WKEa6dA+5jGS6UKETH8NEjNs+zWFbBZKFPO
tv+ILlJO9PX8eA5pvma52JI3iErfa97AjLfscvG0zICvvsf91q9GA+q3up494jzXugdSHPWVoIPW
g6+/mkODFbmwN6PHDo8fI//AsL9fVbd3ghPR+HOpQ5rSxV1EdeFnLsjaDsz+hwihmuLjgXH+LWrb
NbO8CG4W09PpoAPTNnVh7B9z7FyoWe90awZ6i9BJLkwWFDfeNPn9ZcgeN1uG1FN8lVzXKNw3/cUG
4Oraupj2SbSG7MHktRb6NZmUMJ0VElHzsoSamDdGFgqhyl7fZ8jzfTMGDXH81qSCd7zgfCElopPA
gXIr2ajpttPuEnVsC25IX8qOCd9XI/Of1KLe2Q7c43Munfvj+ZP0pGhPMn+uD4mQE1S4neqjD2kf
RfdaPfbGnb/HsNzTxAc6hKmEfAdgdizJtJanC2OZxmAAsylM+3dBBNvXeEWUNzBO14QegKIsGCuI
YyMotfrGWeUkrGqxLEigwEUA3jbP7ZRC+1RojODe/AH1wtT+ISEXkCQCDxO17ypn5hmC8f+CeRcO
fdBt+ZXPyQxIUbOY+17doVxJbvYsxVg3QV/ZW4HSXi4xZy2jrT96br5k3Rw1pESvFPb/rF3Iw5Ep
K1dbLKUHo0AK347ID9/mVhbhPfXSHUCLynYc52rjnJ+WBoRwbPUoW3aWQV2Foaz9uOdIifM1kXxB
PwhD8qYmWIcCxNUwV5UTd8YAnPySZhSI2rnZS1fWdi6GcmnmGQYQMrUsMNBik2zlNst0JV49IsQp
U4rOARm6TB1hgED43n2Mx6AFNrhEYDJmBKTig1Vi4QGnVBwTSBKO65WARo9CX4c7n0L4oLVUPB9I
BSUhALeQ3Q8W/NleaozNtLF0WPY36ZfmOkl6q5nRX4D35NDnYkF4ZZ2O/3Ipt+gBIIagbVSJ0xet
9YwmPWaSPJH5Kat7iQ43RKqcqtMBNszcFfoVRBR9gxXEllS3JC/RhsjNbghkxhHhBFfqYjqJekrU
4Oc/0ND9likJ4HARdQNWNshGD9dkOJy+Gi2BRUMDDD2DyhEhiUYRkHHpMNhMOUt6jRx0J5l/+6b1
ee5Ok0QSF8P16pY4EVvGVjvRypa/YDEGOd3+FfVQ7ofEZFC+w3FEaSLlOHh3oBHd4VvtfB+s1nO4
U3xkd4BCin4kM2BpeF8mr4yCA6OTGjQy0n0cjgZ8LrelNg2puWm9iRkCTLJ5q49L2cLTxBbAAyCR
qenLindi+stR3gCmgH0UWHm9jtxncWm6XKZE526B9yoF1dUAXcWFRDaSnzwx5xC4dM6oJ/9uvJUW
HtTofpUf1HqrI4NB+njKBPHzxWecsWWWUF17n35Kju+v3BR713OW0mAWM/ON8BbPojp5xhyQ4eKV
A4iskDxAWm7maKB6glSCfJeWwJVN9XluZobJcFx1+5t666dmnghWDshLNst8D2RZ6Yi539UpIw3h
K/dzah5bPKwyGq07hqkQs8Qp1Mid2fvjFw/TF5LAyixP9RlkLp0uJfVLwTku88ePWlEww7AcQj3U
AGSaRyUiF22Hn6VPzlzoJE6syEGaFmm/erY7VF5LjF1KmmzEFP2IzUp3OFE4FHzGbmH6XFdmSj69
0CfRNGbR0Fn4IZ88rf2boBqu24ej+lEG8q1NQTuKh1zT/RsTJcGkBHz7cRES/p7wIRHwGk/X0wBy
OvgnOtoH9BFtisP3nAAGeZbdo8FGGzstnDbGVwJcvLJMUne5NFQrcmPAV0rJDW/0PyTnRBNwLQRB
NlQfVvY/Jc2+ZTfUnISSWx0urwGoveoPYiQSD8z4zSC0WGC4SpC9CkADHLHHU3VsO1Fj4PtwdyP4
DRTxZaKzJGXXMpoqZHo+3jLD/kX+qUY0IdlYTAuibAehXAy6pVkLmIn6MPuLXi/sF7PVb0lqYhX8
M6MHNoE6ZzTUYuG3ULsUe+wcKDakFjbWGAn06uii0Ce5WlvTZFd/MWEIMHRkk4rGZbwlgeDvhvPN
lcQdqjHMzWryV4k0n1yvkzLTF5jaPKgsiSQ8UFgP6q54hT/24NuNwcoOQ1xmE57dPt33qRp1njQq
w7pcl/ANpOjBSafJ1FSX3UDLBZy2rQ6zV7jOp3vAgd8xCnJWN8kjL/a8xUXMlOkM1w+2y8oZLU0C
MoU3I2wYFGjPeeGoadjUUfOqlGMWhtnF4krLFJUkHjVzNjWEKd/JwdzHUQCvZk2F7odhn5P3/rZx
lsMq2v4DO58Ubm5Ihn2vmkcJXZ9smmuOdmZm44FztHIX93YO8/zaznNpISkY7xBuUNcQQvcl75XC
j7NVVWAjap+2E7VYQmiUtJDw8QdGZRDMAiUoNqhmExIKrGs0PveTHcDrO597rkOHzL+FyGJBXKw9
95l7z3+P03awtEdL+seqvtzRKeuAYOPEsZLsX9Cq3ZQWbgppOaYLIEloCd6mjizlxognZsgoY2px
ItD9cWvyXRDd2EZvAxj2gp7/EjmsyKp3DsZhWpteFql/bqvKx5v5X/SNqRzYeHwyD0py+vFUlsP4
uBaxo/vDANoKyhW/2J9Ox+LgsvN0klhuWr0DOzaqYoo5iUtaX6E2H41nKLbdziDSxiAyrxAntf6f
ck7B4Kpv9z+F/0xQERXSV8ZZG/OxQ57YuqeWn8zZt1MQWSIqq2rgdDQL5BK21gK5imS74twGloZ5
MwN1z5N9+RV0N7i06bFXQzQZqQ/BQ+n1Zn2kIMiI0x3SVkjX0Yg6zjF9J8WOmXm1SbF/yRcZJWE8
F/hyrh/sxg6ydrllGuUVGJ8xiOJpfJbqOq0ek6UGwN+9oKl14iSTCt1b7GPLsm5X4oackwHEJs2b
uPvC7bVUHxqL6MEFg/LhBbxH5HyEazhFqTuMdFu2OGGFfISDlqPBqJnwwEnygimJhLrgKxbU+a7P
H6Kn4b2WUEQDqPjN4ssl5zembYcd0b1WYgiho+HCU7EWWF0+P9Bu0nOCoWVssQhZFHaYh9B4uLUj
1q893emKSSLPuB7tDo4qyxSP/19mY/ld4l0xtvP6D72on54aDGfbRJ6g67W2qLqewlT3szvLifd8
Dxs+Z6cSeLwfgyp/niad+DXZWMiFmkdOUP7qEjPFQLGF8FboTVQyGyilf1QjSTcUJu4rWfo1/JOu
QeWkxFKdNYzXpVFeg1qwcBZu++9iMj3d4VwXCxBqVNh4BDbyx8wX0QAo11yzhQafgq2QQfaIVvB9
M0kNXhEtXySf+zJ2UZPPyBlmzRx+WJU6zEHbAjPybLlgv49dpV6CW7TaHiNLh6ILaOmtyK0jsh/N
/MU5iMXqrvPMqzkVwT2+mqw2aR2IFMFjJx7jKbtA8w4kwXSjZiMgAzrWhA+A0WjFbmTqjAGD3f8x
8RrdJdjcUOYHr4ODVrGk1rtdpDuiOVZrCR8gaNtrx+22koaPTrKetJlBB3nRATg201eCy2kpm2v5
vEgxlwOJPnhZ0GZ5HDraKW7Pwi7AaCvHhq9vyE5cO/Dql5NslBSbhvWtd6GPFuQxodXMND9F+bFe
gyMBxbn5qdNXt8QeHMcseVwrJBE5u5LASvxCGaUWSOoULR8hl6sDD1EbDuEQZ3oXDZ7GGdsh9aQ9
6aM3FqffJAyI+4QxDDeByhxE//NPZikUq7NJazf+nizpdb3x2wUHWkbHRPIQDp9OTrmoBoZ5aHvI
Ol1yzCc6sjQhpLGhc2fU86OSgY5uEAqLZeQrE1IJ8wdVQ81nLeQwcnVgcq1pXGBBm0vBvujAgFwF
0ZUsLktvOM81CqBouRAAEACkjJewWAePgCqKPx5b3TDHK7B3LCY3T/Qd93tIzF5AkhqKfy55MwEk
0mp2ST2IfujkIR8OFpWqnxjLslW7u0ZT0jA9rZgG4ehwmpyYtrnQKgMKa1dMqnmu98VVOY5LtcV0
x5/Q0QQr97mWEUeG2SUBF/tUfNRIiCcG3eSUFc3hx5geFwPryATv+hGuoZBbmoh6uJEZnzmg06SN
I0RazAggCH9wVl59sAagLOkwLKH/wCADnvH8AJKIhtLDqKLCUqMdZY/Yc3i7YV70r5WZ4Iv2atyn
gQ7nkRM7o7e4KNPrQVnyFn1AfLqbW22SvUkb3WNOADUD3Oht8O0IEM2g9GXuWop1nEluBrIphetd
r4SSNwdAEqG1T1U6U0cUrCFL/6VYoMjkbzAkQLCZRv6SewwuJLlNGFuakSsGLxqi24KH0wx+tUQc
UQwMZ+gcT84EMXi4W4NEdXLnCH467iA2xIatDdJX25DZfhWznxPzb0/Nf19UEPQotMsZ7+vhkfC5
OVu3DjKJoIyha7Aw7COMp/6dxqI6nfcayqoWww+RTUF/3wAujH4ip07Vx//e8VLLus7xq7an+7Za
wgj9CBwpyc6SV229sj1foeBAubOQ1o6GjS3860sPX663ZFiDxP1egcELotp3Iz8Q9RMbO9laLwvg
ix7O5VSXAZnfD7KvuTyA2VfRkGmLLzOUipdFzkFeTIsoXguFoVwra3m0WakC95kx0UWkeimoIKNu
XaxE+pYTzU8DfBLFM6ArqeVBEQ8rn7oLLkesyMvP8PCrc/L/vH8+8Di4aIoJQ7pBBCqU6yrNH84K
SCj8MNoIZGRLUeeHBsrFVB2rTqTw7YqD+Z/hLi896hWxcRlAbWgLcbQ3dgOh6x/q7VCBRVtVq++I
UKOJbiRcaT3DhljCSdg9Juvad+hX83iiejHlRNaW8MgL7n29k63qvbfc+lCsZLKDu5DNkbPXfUjK
B42hmDl3YM1D1QRaugVZzsTw4l2pFdkg2wI4JuVryZM2yaSF7k3uq8I4+aDNshuoLDznsiqARjnC
MFq+Z4JVrPOHRkjLylqeordVhG/qo4Kpjjz/ll8dNfvLu1pDgkskpaY+jPhzFhPJ1tSdkor089gs
rm8+PQg9742/y0bXU3g96Q2cUXfKpUwLCnVNmvHobdPBrInUbbZk6sSixGY7OlaaSB3RqR4FttPn
krfcAy7s27in5fh/Ym2rED8Qqn9xX3KnlIfWrv8dh0fPWVMWz+nJqkFiJJwSYYAxOOLtI1mg8ouB
ceFA9fbFjF/BU0oPWFFqgQ7Os/30QbHt55XHF6xGsZjmcu1p7NtUXrvtstbJH8yunV4JXkZJTWRU
sLhwCDN74MpbiBaqYw+JZHqJ8iFudLGtTA30oZpdk5VplOQqjFnmOQXmvCEaGKZqfbJabtPsAngM
/brb3Fg3bcAI2vFFda5M4ijK4t+otYd2LlToDHNRx/01oy1HJIWHNsEMAoAvYdsZcs+w2i+HzmLi
oxrEKbRdkOCrN6KkRygavN3kA30DvR32YckGtvvb1ULOTmlt99A1cTAT3W4snO5Rd0vmmAerJHkJ
fpLCSyQ9KRv2l6ABlLRh00qH4I3PPs2YLMf8P5Pfvz0dTSJ4w6Vw+Kum3+c6SbcL/IA636Aebys9
4sMTw0raiLPg6WjNsJXYCuCZFROErpaev2k9ZUMhgs+p0ne4Kys8OWDjIKG0U20sO5YJqdGNTT3o
j96Mz77qdOzvUSnHgt10UsTlErkLM3JVWYsbfG2nOA5arcCa2CeG+YRQL5IHod1gQHEivIr8hzjD
/53UXnOZDnlW7bF3AwlQaP68VqmCrVK18Rw0KzlFpKjIxvgf7cki+mtm/S78yRHiyUo+ujo8Mh55
tmvQ31gQv4tMp0QKyb6z+QqZpQqJy7ihUyMxXuLCAqM2mSgEnhbaMQclNjlybShno/RkAD1pKNf/
hrNkW0LYHvupIp1cf7AizZAxQuJd+pmZigcEPzY9GjRx3IkJTFgb75SMwi/KOJ/4Kr00nCTFYJ/g
mB+DCnubzcU+rebbsjzeBXxvRqNf1SdMNsukE3lkH379B5N3tOR8hpt9Pcr/NAwNhGJvPdvlBYPO
GhJxrKEPHLlaO62Hr/+Prh4q0tvkAyiF0r5sUmUFOb0vVnZZJTL3Npoa90bKi2iIR1S+FFFY86ST
Piul9AXiZmlIeXQGxspeZ5DbZy+yeI/lEf4MwB1hSZNYz+NkxgIppyd7oDek8oNLEDLEGT1UdCKG
sbzfGaI/6K7ldT4ITfBsclDWkljSuer+6R7gZ9vM+Uqw+ArtoiOqbZ/2JEMauFj3wTjCFtb9P9A0
osSS1dyrQqm5Lc4nWcUV0nqIQvuJ4y5ZZNx1R4wuALgQ1ZkuYUSt9U3NdL3qluoXk6B8f9RjCgBB
4KUiwsjXwqbQCch5uZGGBBQ6qSF9QfO5vaNiE33G5Q+y2bhZ9/tRszSJq26hbcFAT9F0y8lodYlN
vzfWgyKbl0CikE+QWjz2QOYOin7sFvakGTUKxTg0tV2ZrGGi/RYEOILgA+2G+mQ3CXdXx71aH1aA
suL8t2C/hfUpQ0WojZVBV/cz9vE2WFrMke4XSAa7QFHGBJEpGk2V9iYJ6boA3wnlMuUaZ7pgv+36
0kJXs+3qH6pNCMXkemv7jK0gVElOJewFPFXm0Pn25AZVT5cism6Bk4J1P3ZxZ1IMMIAg7QOlsBcr
F5EH0+6uFUCbUILaMh+ko0aXhrJFeL6idUQSrQHrZXhxaIB4KS/P20UE7kymhJb0/NElkv6CsbnF
9TP9XAtEOG95DEUwWP+3EuxhQ6gjOXDc+mhwabAOkmNynmrOBYgdrIesALYA/aoJuofWwyPQ+ljf
NRGiuhps38tdEieg0CUyH1rgNW/EzHGYznOZnU+1wO+UvYkXKd4Hl2/3qL3NJR5MpkTuS3IW1Ju/
Rq1IgHbxHRIc94fnfInqRCrREVdJD9PfhnPs8xoUp8vw/j0Qsngggyg/ASnBHpcl+08MvYBi6A1c
fwTGUmNZSD4KzEa8ZIMAa+F3XrMnaSSZBz2NxsKts2ixRttrxcKnUJKTUrX8SnL0NwfV3pLVoR0e
bIOL/FnIdMj5byVuJ0MueSnzekWNDoNDwHqhD+jTNVMAuZLgFU7bU2qpCw2AXr9JZTnrOfoSue4V
2ZsPES3+xMcLe4YSdtPjTdSHg9GpVu91RxkovSM1vCRbDpdjeOndTQK7I/2CoF8hXvAhCOfPVdoH
G1kCtgFgwxMYD4HfLvPQ7cjW4blUPffOP+aRkhHtnRgP7yfPe6TsLdt56ruuE9oREXAaOBzyk/H2
1iKmqDdlccH0pAya71JSrO/no99BG/ppgTFU19rSUGiDVF6lyrQTDEGn4+hsDk6Wu1P+lUtU20QR
95gpxCtvNLOu6PMiZnvRmt6ZXK+Kk7lCfMsourBSt2uRzyPTHPtf7Dne1/dqpCYE6WkKm4GEY9jq
q7C+dfe89hrx+u7oWHlvc/6HlECeVslO0dEud/dlOvZa93hROE9zN4wv54d+jx4BH7W8XxURTFx7
Fmwv6jjppRv6MTXn1wcf4crW+3xARhK3N0N1GaL8LmCp6PteX8yzncrvGxN0rv/HoxmWnWr2mnsA
33jdppPo5Nc9vn+dLWGCrmW/m9DIZpRAOzWMDs44OubBjc8JElcAUB+EVwCWyg180bAvOTIHeH+X
o+SFU7odwCRamUB27qhJEBtA5CcpdYk9byIL4Tqdt1AV7h/DFvAiXcssBJ5X5h0sqTWYsrOsdqEe
D472Z8wpp12MmCiFhGDyY/4KKELb3z8JItnEvuzmyFCO+g2bG6F5YrXu5z/ggyAVkwpdr85uw+F8
9cNU+B184BFqvCwNwVJlThJITuIaC68jFxhPg9UT4vKjz5Bi5wmlPeANCHBBXxCblMIcssy/fQS4
d+2NlK5UqHk1cOsOiAzdlxxWInMoKYTri5eTm/reVkePY26U9wczkQ/u7kX+4ajtFG69YB5HLwFc
HjMfBaMxRPLb4PBK3PHMfjcYEs6VKELGAOJPaY5im01G4yKYFXBY+CR/Jz+mOX/E2GC0JSgiaJry
YU97ageODw06L10cgbVVRotd7aoP5fQa4yFzbzg4X8Kv7cJiVPi5EWqFe2h0mQB4AA1U0hjbKWtu
bG6gwd98S54QwEXj+xXVyAYh8nZVxYX3goSj0vyVD21CgyUBgUGQNRhz+9vwxkxTbh24fKWAH41U
M2GmDyGvOlDeWxd8ZceEyPhiVKzQUjy8fUhLfI2/uaWYM4dYTced3LULUmRo6c7VObF0fRrG+qsN
UPMxCg70RzsLScQMhaHLgh+WI87SdkELmrmIW2KPTJSq9YUpoJJWCnT1/BVlJUI7plS0WEQYc7Kc
D9SCinPpbzM8QVMX0jH4HmtT8NyWRrjTtvS503UqvbnPhCEFQ/b3BwvuTywIb468snzMlGeSaUj6
aHakVYfhzwH4GdK1GHKUVxlu5yJiwa56EQ4CWTYosLw7Eo44r7mUsKgSqsdB2KO1kBr6/FyO2VoM
ku7Ec6nQPBk39tu3BMQ/MVVuIBzPR7s37nu6fc1J6TSqnILRDxNH/8D9bt1deJ2BPK1MGRegsgJX
wiHgoRZHjeKAV4urXzLmU2yVk6iXWFCdWEBOeEXcDwJf1KHTwG7zukav/KnmE9fbzIE5hgVBeoDa
wMQpLB4F7zwyUZBiZjbuH1B4fwn5VWS3kXlPX0iIBmMljf3i1wrsdgYChX2VzyUfogfKsvedtaMt
u2hBR3hg4R6OVWYSnIRykGZo8ESSFJgbkCkEodZY13pWRlOSoBLdSY70wU7A68C8HY6krRBVUFKX
jG2O6c5qIM8SxpjGaJ5ZssPiQrKEXWmw9CgVoMAGpUXO++/zroh0hiTz2hiC+U/fUvOA12YL1X7W
zoh2ZUiJfPTKkY5DLDb/cU2aVPYKDUpeRY0/5oQkRhLU1jCPct1ryp2+HLpABwJuIkBa//9RikWb
/+rMUa5C4W5h4nYN1v2NlQLjB+L+1kfDjRDG0y7Qncrx/22sBvD3fHGZ3+HBy9dWaG6WKxcyIFLJ
rVoCoFMUxIAFY03PJ6+2ApARdS1gWFpOdMy+SLR6EYXkPVlJN1rks6ZkMYpWUSk7ssH53+zteyzZ
QS2TnDMqR+4ZV4Ip5fbpb0sMlaePTJPYcwTGlPfehq8THJe6Al++AsxFG5zw5GSUPzpRt+qTJ3pW
OIjYDAoqAYDJYg1GlPvWTSzxJe/TDiKfdj1A2m1+vbuecvzOPG/HrE2EZTiOc2CWBooUup/9GbYs
ywZMHGKiBkeijvfoc4QvHKmpsVUNANc4sX13g1MsdxhOGIxjbcvdPnnp0w5z35fXRM4xPbnpC8Ky
1CUrEZvpmkX2ceJDGq0bF6ik+MQq7wLf90NRq7HiLaNlnuqiNf5FQleV4K681bos3eY+ZTgoxctE
15e2t/v2hTFZWEdSw3AAmydM0Sg1+L2EqxzqQg+09y3/beEBZDjgnfBEIQ8w0Bl9x+f4On1eRhGu
lzdVml/PbGr5Fjb35wqaGkUuFVHCPy34lT6t5m+LGOqBMZwSDeo7ImXgS/Suuj0J6FdJ7y0z2Ho8
/38pxb7CO5UxTR3cMQ6L5z/a+dqGTcZiIxdcpcM2t335YWklVGXyiH1Bi8oQzq1M3RCyhPTDFl5T
8MM5HRNuBVPVl9SJ9gWfq0Cp5SzVaNvtX2Sptl5mXmTABM9+TSFHExRYkiovZA/TCEwM3IEOWloj
kDQRgTVo1HPB+ID4/bGEL/epY8Nrt8Ui879rnBPNPlsgv23AtUW/DVE+wYN7tVZ8HNl2s3On00ky
Gu8ABS2IURh0juJ27LhWJwLgrAzryWXcWEiey8P850Tm54DgfJx/OiOIwkKx1S9/1qaJdIdlk1fz
bRw6/l3Q5uWwr/8TO8uq5u5daXt/NglQ2BKJ/fV3rpbg5tApuHAbPK41+WA2IESJcQk+XlqX2pGV
y3fL3+EZmb2pZ+Nyr8x7olnz+FuwcyIlsoA2PCfu5JrG/+WmYjYRaA/Zz8ni7x9aQhNQwVJ8sf5T
qAzOkE2sUhbYeYYxfBH9vjFUYLOOeAX8zYc6PPA+nqgE5EK1tp7kMj8/Bw//3zpmqJAsnOQbkb+B
+lbALeWhnyIiq6Ry9wZbqrWUXa5SP0Pl+yy59wE8AflBrN4gFf9p2s0EQhdZJQE4N7KynbyY/MBI
28GXKJv/15ATWaZ4plGjgEcaZNDqno9Fm7OLtzewzZMLlIEzZjzRJZ8uOesPekms05iz4tV+52V3
LEb4xMQjm+Ql/ZSvPNNkQL0I1+5ZkIDFf0W3dibUiNz2qlwkfgiePKkk2G0jpFWb3h1JZYOSdXVN
XhuO0UexHQtRvgjCYL6xfEqq2L4YoLNJ608b9GgwSdyBMwiRfjk6GSb+GT417R4N1l6pP07ZYRmC
dQ1gDS3EcIMw/VN5hwulegUXXi67yBN+VvSQQSSjDRqyCXr9FBdUbpqOnn+fJzkYDRK+Ok6026PO
z1nNjO3NU4XaAGjQWF+Gs3gicuNySbcy+OnoamVSMuUu9BnT0zRGeYPzpb/ZshTCEw/0QxYE9NqG
vjY2XS6OYYhnOU+Qjy+CirEFCvDzlAsJROO+tsbgeL4QahGWRst4+EwmH7WGDriWYclk/6ugB8OA
/hP9RRETkG5+KwA5rnWHi0GG9E3Q9LIdl+OxWn4mTNeWeXx3DniaU5RBeud2y9lfpZaUgu51uaN9
BgTIhzFnoBYT3Q/swYbfyfUz0OlTs71Vrjm11F1uHwjkX52+dJEiJ5Yhq4F8/74kHDnESLn8f+Jg
y9xo0E6n8ujiQNhMUxE8bdiu4yGaR/hVl9yJDGS6KL/alh1VzAzoLzS6DqQfpT7Q5y8r+BQf2vTK
Phx7GQJMWVIwI9QpTpBpEaSv/ylODfCo0MVgNwKpOwVjUKJEp9r7X8M1SHHmu3lbtd0Kgmj1zEDh
B0hQCGE4AkM5LrxZzGqNefhnx8ikcv5bN8xrImsdPOc2mIpL43rtkyE+1k7HnMeGrQeXn9yZXznX
SrC7knR5x2D4emQB8019FYaY19cVVNJG4rZiDJdZWrCbDyjD2MwG4rXOZmg9xf14VquhUelTkoVR
thSHe9zjclHlX/JJQc5lKV2P0oM9hE+eXOaOLMyehWLxB3PZrfZ1YOusLJpBf21WDH+tXfDMivME
Vdd3QdZmCsh/UbiEJFECGYTXwJzLE18rm8wYorRZe/StNSkKzHIvUNJ0zB6tA4VLjMmBoiLaDBze
1OyCJvFm0E1FBFoV8fnk6rGsd4k/XC6fJuIsnIfndcXJy2sO1iNRAIH0Je8xk4bii3yfq1QmroNQ
RT7D0zaqDQ0SvcNPNthjCm6XyepmQg8mzGLZwrFJFvk9cT8kFHngl3SPkYbKN9RxPko/YsYCteMr
m0zeWB3zogAMxgjtjtFKiZ/xupOHZ6CEP1d6jsXrYgSRSyELJHERAsJk2rXJDkgDhp9UM6Lpzcg7
RSu/ep5yYCVqF9WHBGFShEH4aELxzzor0NM7SejckrVLaQE87J86RJXNp/pGZuuF1zGsoyh5AfA4
Tr045SigUrppx9M7sECSXh1703ABVKoGYfP3y222Snhc7fRwzpgPjz0shVQ+qS3DeJTHXB8yQmOE
IbGVuEYLfhpoERAJUdBS6nxsaIrSe36v3Fg4sNXgFsj4q1NPHjN2MlLwgzy92DyS8U1Qup3TluLk
Ghx+D72ImuyXS6tagqeaevTkm9S2B7rxh6dhiRQmraaJHKn3zYIksZiCVRvikW4wRViocwTsMj+u
6Q5L+PNFwirUhBQC+qGO24QD7Z9321FUFx8hA+HwQsCSyY3GBjn5RWwcgRfd9fwd34HwIugRx0np
5sRr2rUzA7Vr4ICoP2V5rKQqKLAq2yXHLRZidjZCmmw95evemYFUFUACXWhM5rOx4BQg5d/1TCY4
p1FBrl98txW8gdLyvUvrNftF7UIgp5PlQcJXE8AbuGklITqeRvEL8KMS9F2icnZpk0k5kiGur3vq
nVhPZBrLcwGDUrh6WRAQT2NgcNn5jEfA9BbzaU8EjKLTRbvDhNAT2zUPXc9w5jQGqnWzDBKpK+2W
2MFD2UVeIWMSDbTRWuRvZ+mDmqTeKTrrXCb//kC43BWELZj1R/6MR8WQilLKiTjBbbsjI4uojlIi
eltLRR/HOL4D6ppU6gFSqsCZjOXjOvD4YoBAaaoDDz/ovY1N6xEaIa57xPnDz4SHOUlk1pZ+GMfa
mujmNBPdxFCcGSrW0C2QfZJm64zv9cEQndXiuwCD+KEXYMLEfHCoUCXl6/gblh/4VKw6dyDtwp3Y
SBSm+F2YpjhhhBhcVrA+LPYcHO5iZn4UXo0skas1/JiQ4M4Wu4LYdPLPdhEX3ufNrG757YF05Bfk
IDSEIli9muUuvi/BcjEKJwR0XLSgrZRhPs1UuJbjQV2NJVK1FKPtx7/iGSdcDKcCKtX/KCjJei0n
FnujmLQz5T5uP+dORh/f3UBVPoRKfN0yQNFGIsOYH9o6l98FylwnI3JFkmre6l1EqrK7IenN7mMH
op3YIzy4T9mOeKRVc8Ge3PvMiPOlAslCRh5oRLHxDQZqUiM39WUis0PnvFAz9n3K7aspMjglxzvb
HVP0MDSq4gZIUiXBgIS9o970L5SqwBNGk3uZaw3Q1JbmAChZK47StS++65hsEjukUoAL9fdKwMcT
5322DtkmeP3L8m0OW9Zat5dY2srAJX1/qsaR69wMIUdzbn0YlYjN5K6O8b9ZOFAijxaBOn1pjREx
teF2wVZPg/oJL6zYi9WribfnHCCyO+iiBhcIMH7k/ujWzhnfu9WSVSrOh/ihWoroi+U5WgFcY22c
o1kSrYugOVfUFxtpFrcQ4PRs5QdFHkRtTRiO1ENwzjplaP+0vrk9qiC+EWbXoLMszmCgWMmwWHJh
X5CcpZmVZayJ0DFvDVAibiBCui6DkUkwVDW/zkb1L3CCEN69BdZsXQ0wOQ/kGqopD/8UpC0SOS/w
OM6No+O5/B3Z6OTjSrhq8kJciid3SrTEuxJrH+gB/z+OVxbCAdlyUGdyyT/oYScKIf4wcfTGHFK5
ax6xg/vBVlGbVOUPvhzzxUZPo49dfQ2XJl91+IZXoOBerTSsuFR3A4qs2y9LwkbjtNigJGX4VqEP
yu+jGGtb9fgD7seW/Z0zEALb5rCaOgwQmseRXCRZ7YlbUJ0PlH2dKKa3t6T3TqL9d8/XygihMSN7
fU9WY9pgU33dcaV1kgSPFXgzzRiAFB6iTeYk0HhHupv7LoHlCAl+l4/yyEW51OvIjO7HO5kDCuWA
BranPRzCG805Kvwah/SeINp6RsbBF3+5E/08slbW9CAwZpTzoImSI/Ti/bo9U3aRaQdNqNOertLF
BvIaA1+LgXZ+JYG0Ymy1aBXWhJA6Stkt7BQxHhkqPu2uXoKnQV7O5H/Yj3HLxPQfg7LbWIpod1IT
F75MAcqaNLS2aVVvL/davjPaZPDwBP5860Yue8PrvNdP2cXDHRXDMwub/L4+geCH64KJ23L9jsqm
Bi1HNHiGxksvPEiKNzlSBegPABefiP5Hz8DyGdXLxPVViukGD1CAL6YC7aDy72RtymglMvdGJCjy
LxHQpIF9KbEcabPPfxHxkSSK6MThoPauAsy03XxM3234PVOQFu658R4UNa14zJ1/QfWnMuSQZY+h
O2hDp1IBb0ygB5ScsNIRYWPJKnPWx/Wsv5IzxoTKKQDfTRKpjkr+LcZCYrnqgbpMLYHoEmPpkSlX
Pc6cDVPzK3DK4QuT7srIXxTSgN3rnzy3Kv0JHo1hPpOy0e3Lx99AfULsGDKalgzu9y0/z05rwbWk
F3aNP0dsNUemQfSpumcQskgVoIeUoz0eDbAFpO3Z1UQR0Z2ASJ7ihwmH26bocDnsTc0xXqntIckN
OQIWF8FQIgGZUaeHVX4/VApBvDFd4sTgWRErWodT3MIsgFIXav3buPpwBwJVyq5dLsFkz9OgMSmR
ramdMABV+PWQl7pMMsFfY+KV1S7AdwGo9CrkSbgopoGboVwJF6vbpOwccTcasdbJSFS4e3f7Xd3L
LQ2auRTrz3kjSXsnnmi0srAuqqildc1k5W9m95vyvZwmJjznxiWLEz6+ur8lbThOUVFcc8gmmF+V
xqzi8sBsLLg3Gmmr+A+ssXVvgpJ/ch/rHTy0BRdyJjY47cTGy93/Fx6zBhmTt0GZX7r5VFhetred
mQYIP6+qKOJsgsy5f7be9AfNrjQMAH0UVgIcMThrBWl5A8pYShOfdZLcXa+7cz+Ak2yKsHI5hJCg
EifDNRu8rOJy/l7wbM4LllS8TomEcyTgHS9gItdvBa0cJV/++yZOt+u91Wg1IpLR6T77z3CaMHlY
kP3cRwFcgz+aaH3soRuE1foEKTF/jWP/hITGqCtBNSJCxIaXHUiDhSqXlZ8YH+6iXxoDRrXPamR1
kEuqGm9GZkHBsiHFmpUpyLK71L3f5tugPKr/DxjyrLFb/RZBzZi6G0Zc00oVlbqFlRPD6OeRanhj
DUOrZD96LsKt+qhtT3x7ppw45+mC4fj+PSPM3sLFDr1dc4q/h7beo6Q2RZmfq7ZC/bfROiqLcHhT
I72FK0FDaLDeeMPwG24D9F8rgG4+cF5nXc1p98IyqJb4SMr4IPUk1OZo/PAcIbN7v5WFPyrMNheG
6N2MCi820HOw6ytHWl9eG3gmvp0HOUrYrVIApLqqH2AinTbVRjVOyzFG6O+NO1r06zI7kCm8G0HU
wcD43TplF3XGz3p75+zqSv033GEAYoF8X8co4Vhxu2bLfsY+MvhaJWDqSzv+0+Q8KQoauo1NwzCs
CJ1xh5eHzHkyWX4YPo2VThjAPVX8oZbsvA3Zg4EsYaRs2focn8wciGTKkBTsN6/CW1+KLxAbAxAo
xDB1q1rRiGnrV1uSyYJ1jNhp9vwAZctvKCjf5ZyZDXxaMY72SHy9GRlfAsgyqHT86URGUuPzSiIy
HUlmcub9MsIBKLn4wfkijilw4b/pbtZDpdkJTjF0YLZs6WxLUrtfSlU7ufRvOghJ3LZX79R6OB2j
XaH5s8C9S9iIoQqt7jlDFE2ZEZq2EIXuL85pQxK81MTnk9KTWDUVSziKbeULZIcho/reJ038+5Ae
/QQBjEyEuDW9MyRCNtmP54V/fUHcHUlzR1C/DnPunGioFy2TQ0yPc6lIDgtaaYNEB4uPJFfSTeqQ
WoFB/ieqw34lJzaIOijJ8X20cvoW8ifovu63FG6eiGX0sg9Kw7qJixCIxZnczWzwd3P5wtQpdgRs
ztKtOaxJl/r7op6ta2t44AmgIiSQ+dapsWnaghgIzYa6MZ+CsbCu6Jc36nAUL7CwL0tsvSUYv+hy
9DdlUpI7bsXnzLoBdKgv69W8B4bEk++wDGRpCF9x2iwPBUe49t0y8kUMeC7YhMA18292WyFD14GV
b4OU1jjQEQ0vLofXLK/TdKmfPzS2CBZDlyrM47Bh+/Zq6OlGW+NrL2JsiIkCocxB9ewfwk/xKStG
mukJjyz3UiieqOZLYIEIuk0LABNjUaQG8yxmmKeZPh+sGZzxMrrq3Dq6L+HSzx9GeURFdpmozrhL
HtDcpw6nWdODaUX+zlNgtTNOEBryzDm2ePlMA0GnV8SZr4+p6DA/CcgeFbVHotl8Z6G+ztp/4Cpr
AkdtTVWwKpvEJGmpwfacFHug9TbQu5/Bxe0lHrgbGd5QgiaFwVBqHEmzEACOcSr0FKe2rV0GKSeC
ElSxVYvJMjX20QVkZHjByYqcPLEnqn4usjHXzwrIK/5y4mgjXEgk7mtrvqWV9egbBa9Q1DlTPhou
PdrFIHVajnZ49kBSAbYDmZWaKz+y9o+OlxUrRqzNSjlDZpwEB8rDheGBIKZRkjSSYAf1zHjuQAyE
uGFDUE/KTEacpWaDTxUuWn3qVR4B6twWrd2APrVPThfOuEBC6Cjpn19bEf5B6NI0U5WJJEv5WwPJ
q9UNrRVjEOZ1TJm9J9RsJLBjXl5LoYU8gxT+f9NURzhe+ESNVQRYjikmU0zg5g/OOu562Btfh5IF
obspUdIoSkkmLMJ1JxADYo1IOCEbksCMkhCRRdvNxURwyfN045b95SDpsD+qxrg4A+bOpHrGr+Qk
WRsjunbNNuIcoazZZUUw9elGLH3msE4ig/TMSOUrYo4whwQzChz36rhbf8iWTah6VjevNivn31x0
bmkc/GLETmbkcB2ZXGPLxJfu9WuvNGHCg2dLr/bPJLrgrsAfzaRY/pTuE6EjmcnoNTHe3W7aZ5DG
J4b0zPaEGLMSy6n+AgV3xD7EU2C0S6ry7mUbKFWP/NJ7RK9UuI6QeIDVWKfbqC7L/huTjBtVv29J
oMYktwAe+LdfYSdPSSUAYA97NL08T1BDdkAKxY0vPKnu9om+DmGGF4Uh/vPUcOzilzKdAe0S7ZA6
M9daKPQzkD/wxJdbsjfmLfwJ7VxLs6noYrKdRJmIOgs/K2/iHjHSVKBhlF5vG5iroSjvhhaRyYtM
aXnLQKaBECVu0oGNdE6mBbFX0jBVKMNOsBVl91QbZEdVlC2GYSZsYr01lkN+gw0N1D5xgpy2b1FW
ziR2d5edoVgMdwcF42lDc/lIjohqkiuJ7PHaHl1otOUPiQjrQk51I17c9lIP+Xwyh7ONAgru502G
PO66/+DwtHVKDVxg7REguiYCYew0BkqRUq3HCWVqIgQ5WQP4OiBqjZXGz14AYBbZBS2VxVbgwknI
AYcb/jV/+fpVjVXJyvYFiIWuhr7kHY05uLjIBcuFsU2D8Ps88Er31rdEwHHdKxgfobc3GNMZ+hN0
jOiwwJb4vOpSehD6cbBdKTz1w/sidPueeOVh1Onk/Gf7cSK68cDBJPday+Ca9QXuCo/C1ukAQmFL
Q05U9OJfgeSmnuFqZPrqUMvUE2/F2gghDF9lryEP3RIX2K39oO/qWxjyjPwvs7hnRBeMiGUYm+w3
uDiCTV2JWDDPs1lbv5mMJHo3MfrBOW5coiP0ty0Yq3hxF2hRfMg2UJYAUAKPVxbS68j5XZt5Cokl
YBHjdk2hwz2V+CwP+12EATQa00GMq1pR0YYsspY2jolENabNVA9f4bLpKNEYVsFA7/t3dg89b17+
3Xxy7lK8it0l6/c+NZ9yJ7oCSMi78j7Anwa4712gchAW45qje32yviikij5K1uH4pS9o5kXBSLYU
qou7I313YNx+Npk05DOnDOVEF4WMaqxEsbSvZMIs5YO+Na2MPCpKLg1LRknOYfLvzmpyvox4K6+n
FJe5P/COAnTdmQz8DtvFFB/pJwD+xMU293t4uMxpV/ZPpxXcaaVhAlGAa56/zkSjjeoBxSfQyv/W
btyRK5l7Zu/seyRtCbUBHstossJdZ0bf6jQ15BM/2mHXJ3JuI6P69+KrC6+Fd2MC23UFNMRSFcWr
GC7T9BJHd7RbjcIM1BNUVr9VtCsioD2KbaJs5JLjVJUWXNzRzp1sh1gj9gWyPr7hYSFBLfiO+lnb
EXAWDbUddI82k+a0PaZaBRapnC9j8E0qU/+OIogAOAfwKFHFn/vyxjHvXxqqdIBSDVCJPaohrZhE
p4bUXZ8kiPeos49adGC6DkC6O8XHZ/jsa5HdX652Gfc09vEVMB75liokc/jFESlWtIGuL/htSB++
h4ptxB1GZCVIaBL7TgUxYBIAJ/9RiZQU35xUtrRH2zQ2ui0HleCxaFYAExgGEFt64K4p0ONSS36O
LZJ8jFzvZAn5tMAM8wPG/0iyelF/Rdlzpk/csCx+3pZhz8ATgpCYkqCVy2Zkb5vTYUkftnwO0Sqk
KyW+T0JWjl94tibezRl2xFC3RsL1gFpdKDP2+++lOes7lt2pl05PNpjh9/RGWtzHZmpHW91GgyDw
C8zQI52pCrTAdgJZVX+6iew1qWIEZZKEF22ghENZzo+8FVZzvR3iprwNruDdCyRdGueaqHqahcvN
PKvUINbIBxxHO9pAFdH7Ct+AC4k1W9pLah85hOVNfkEejdWnJgudeMGzcKRWOZFybsZ5lY2OyehV
FJITCdbDChBMOVr/MvlXKOxMO966sj8Ny0+Z2JW/FyyxMmElav3M8VRNlBHQfH6e4E8oNGmylKwu
Kb+Cf0NoSIi8zVOuW3r5IWlvCdqnDaMhgOQ4tvdQPXOFay/8I+OFhw3FMbZHLOXo278FRKa9MYjF
eKm5JXHtWS52qAep3+hjlYGDb3qmUyMI2V4Bw8+MDaR4lBQFrZABpXHVfRVDtU0HTKbgsJ41/EeN
cYfRie4w2Ucy+DkPTAjnOhnXiP5GSqv3JVTRwNpdrr1qiqD0Zd2nLenc7zxGYLjDPuy/mPx7tuyO
cPVpbUOf/rCQbKtd+Gs1Fs0eMbmcug21htjGwE4hCrh4uFXgAw3nRvhLlOGgfzn1BLDrtuppbmOa
Ws9EIH4dgJvDx4Qu2UR+OMWupxhcCAGKNFTCMiSui5xp8oQkyu7R6rp7JPSQNbzP7ipMYn8dWH4W
i9utxZZ0WUuqRF/WjbDUpU06gbGsqkEUlpSDMli5RmdupatHITlg4gFKNtESqf397GOjaunx7DaS
LNyskpaR8+NMglEEjH1+9ZPQhVQb7GgSzb0E+s10Ubr660AC0k71hh0jPNZ92EMEe+U1EPNvyZgj
78tsl+rp6o36tth6XU0RULLkERRn9RnntCHBawyIXA9eQnIF2eNR29o74gEagzzqxdhKtKjSogko
vB6zBEkTL9iGW9/3JTdelfp9FzTSdKJR3f9N24lIAqd8DjGCmiAkIXk4Y3GGvNITvePqZtF6ADau
WdZWGRgxGq6EIhoK7s71oBPZsOSixQ5WgjOHPCxgkJxfSR9ViX+R2bRdlp0bKhLgpvttvoMLyBB/
bmGufS21IS1HexS+q/srkDBHqUrdMbBTawfg8fBi+zLZpPaFIvZsL0+zTThx/ZId5QH0lPu+Jf5m
zZUxc2eh6gA+wfG+EqM7kHbg7UX74Hp7bilrRNTc9Vw171WZMw11TtSh81z3GTvoPtgSUoIfTOju
0XbJB12YKGHnTRIVMxg4Usk7+PhHJdDf6z8OpcpgQaKwLelXOo5zQzdhYNSEqtZiUAJiRhpCSmbB
HDPSF9FyPxdvvI5QrVz1F9PqUNL85nw9Xk8pUtSuN+1dAWOkzZ4Lk+JzQOb6ZvYAdD/l7vnj4Xot
jg8LRT6U4/H0lg9ss2rPpzdRbgFZL8lmegG+1QgttJr8YO68T/A/8HELfeoYpmXD1gVyjBcEHiYe
/1gyxf6kOiWBykcG5hWQaFhlSIgpXfZSBGTA4H0mV+hrsTIDyNiy5dDnrIW0ayIjbrQIUoPOc7vG
7jbHYyFjHPTs1qAuFGM9eyj9Bm785T1W2SlxbILxc+D6fRYcTJTKhaKOjkaM/cGkJDID2A4FahxL
rEFd7Rqm6OxxHlZZdC5q6O/hEtf7V06Kzlg+O6CpT+lINHr7/owF1bB3mERgEnCtu1euaJ2AwRPf
TrUiWP7leLoJx105Hb5fZ01jpXO+Gf9H6Gsb5cFI0xTYxVIlAt/HgzZGt0hnaS4jL53yVrnNYHoj
xMv/T2/lwMbG4V2rtHTbpMsPiIELnBREzDUn2FJqKCTbbYaolqpbRO8zkLfMbAHHPpCnU6iC23vX
u/AKF6GjLriSe5xeL+Khg79LIm7mXSt5CGr18d4amau/Y9/Mqw4qiICaj9SSExPALd7hK1Ha9loj
xR1mRTaqSkyscGTlaCWkxjFcYP7vPS0l20PTXg54TyH5GzkQ8zTSsucdGbdGD0R98vrNDjkOEy+Y
Mu0vHrUSty3HyMq6no332ydpI15k5DYeD1QbsBLbVMLearWLXTXAg4u3ESTZ+zHL8WVPsIME88nC
Ba5gaHkkO0/D0NrATfEIZUCbL36ByDwPZTu4RFz/IGJvzahREU/1qmcmtnwvcd/67wchn2DwDoYw
LTzXIVKeCWo2ZoCfF8Ac608j+p+lok9DFaRakbdOAPsWNkMsfA+OLDXLF7W8cCu+v2OTJJ/2h+rA
rKdnUJ2UInqoWlrrX/sP4cMXMGSJmODQR6w0UL+ojHTYOO1Oqlg9BDYcL6Umm/UHEKxlaOE8k9UG
DpxCWmUM6gC2Mk+hED6WvJLWsrlJ+pE3GmP+OJANfJKcUxQ0yGTcDM3I1HFrO8Rw2a6d0ShGS++V
X659VDJjoGHWkb7h3SCtCntDhSdZuD7qlHbh5vo6UqHRadqIKFHSAOjl4BA0ISMsBeyOVNhYdfTG
ABdU7c+rQtcAaK+2kL5I7rVx12RHhQI9d1ojjsnwMKjO+LAcu3+Eu4YwTkzV7Q0hQBwjb1kLE0fA
yCYkW3GBEc1F7r9hh2E39ZakHQpjK7P7x6+S9FYNd3+LLWmoS/3cyLQA1OFeTzY/J00JrTqvjg7M
fp3ricFFyV0va6ak0GWDZ+7Ffn/Bk3k4dh5xs+8631ojFdoWcOnpv4frnpBsta/9Sfuc9ssVlyBC
zcBRs9M8gHCsTuSji5wilW3J1Ux0Umtd7pvhoMHoutLPOkjM8f8TLbHFVotww4SPMGUICQA6pJtQ
dmdN4fNZcjdDSnt6zmG50KW81y1oqGwAn45rPvyNybBcmCSUz6/+xFlsQnY8af0HzRHIQUeeeLxG
raufpqUFU1zOPkbpQtHVdUj6OIhDu7KC8D1KCmqMxedhV9pX2/fr7Q9PH32k71cr6HCcx9uGPyGD
bRHB44gXUZ6tvPpP3/4xqm9qoG/k1t/ApUJFzRuZhew+74T2F9et3W8xqVMJdjxqz5EFNJeJGyzA
3CpIvAciIRuNoqb3kxo+2FKMMJ5JdkdNrxN/yVnZR5OKxkXgF9BKHvl4/NeykUzkjOXGDdptGFwR
SUYs/bYXxmTaQtr1sSx/54OelVd5iFyTMlOLFoD3RMiYfLKr2n+GZJNwRLtiqPqhczDuVamEFBUJ
P/IUpqwJLFUGoOKyFO2VMa6Idr3aHm6u0ZgcTnCbiWkW5PWGaUQNWLUh8lW0eliZjm9PeAVFGO3s
FQX0O986Rs5L9IqX6oozYhN3IC+N4VQ7VdWnuPd3Ll00Ngek7cjhm3hHAS81qaFV4xz8Y4nanA01
DY4Tlokp3PwARwb98wh8ktyWcC073BGC7BazoHKaBPtNHfmqn2gCX66pOvwoEF/r2zVjpCxAdIJk
35eoWUpYYH+qK549vsPsdjSZXu/q/KDks/gyP5aDztW2JpGPMtDP/t/1RF0xAgVkQW9F0FgeGN9A
ilUw+ziU4Cfz74eRImxIsMuiY2xRJHl7rSzSzkqnTyHoqjp2dLuOxCBpaJTwFvN6uNuStA6Y++V4
Wb3Yx4WQSWv2SmPcgyD0A+OQmmMmD/GXGcXbfXETZftaXDYwfpq58mtOSqKMDgm2sQqBqpBbkk7I
neIDZjvsnQWoQlglJppTQ0jOsr8KUGr4QrPp3sfvUY53qJzgcu4GWyMGvjwip8Ai6+OFOyz94mSJ
F/hSA0N5NbGuLk1h7+eqNZP/MqzF6YIkIGzx3LHCsiXK7E2dC1itvYo6w/falTfS54ojwQJmgrB9
ty3HwLm0K9C3/0gd0T89+h/fEetckd9b9ptU4E7DGUdF+xiXYDffP4qPd+xftZ4gyBglPEaQHxa4
0r0KwUP361qnm4g719WW2MYzxaTbRn3eKYbIIrV95dUlpzU1nmTN/bx0JDfd974yWNPZoP8OtzJk
/HydZwDpGcmIh68ErS5K5cOhcMrmWiBe78PJnodPIfE6F+yo6Nu3zSaZicjw1AzsjEUaTWUSpXyl
tzBPFiFY7oBTBPxptCbh6HPKxEAsQgkzUatyCkhTTTVitegYp7qbds4YJQ6096hFpNcp4HjmBxmZ
cZn5RRwRftP3NkbBJB7A6pSSvXNr90Ue6CBx4Dv5F7C4ny9t/Hh5fBV8vwMuasLka+VK96v2bAIR
DveHM48LvlRg7g1qrMYP7cKYeirmbGFfTw3cFiXjIYawmC9dgzlBTUAyGcxxnNE9sRe0Y2VCkrQ3
2vMx/DhgfcRIRdAn+RcsJC14dJJYz3KO9IjzVx2HvlSTo6w5Wn39/TsRBSs8SV9nSn01gsdRQ98J
oG3Lg0Ahm+MZ9U7TUzdad79yLAf2J4IlYInrTZtVvcCSke/pgv9+sfvh86iJNTsrNaIgycNLneUj
aKDr6M8nh60OMUSsuG+QR+4ijQPROSdJpGS8QcRFcdBFOl9bPlP7nLGC1HExbx558ZCDrCJpqcX5
kmbpjX4OyIIkxcv7hp+ZBDcAneNHwVV3wyQH8rqP8+Gch1wyzT7jxXbfM0dz0pAgjivcJrjwyQcZ
bgS39gHxxNXml5BqlK9yPbD4WiKyJgKDl4c47ZIb4ur9L7t1hXCQAzLABzjaD1FLv+aCyMINJ6OV
ahi+UXV0HksEZAZRKZMco2PlTtbJ+KLWkqPPDKq3OIzSGNY3d4ZGKCOWMmqUqrLfj4Hqmn80RI/s
sVjGEorYfVj3q7m0rShTLQpGTFlojOG/Ge4H7cXVDb/qXYj1TkebElhG+c1EsOg7NTOBxjtIZoAo
MIWQ54CRx7KZnnEWTGA/M0EWudoe7SY3Rdpd9+CI9oXe/IFQjbwTP//T2Moe9xGnNm0ITWuS62VW
bli+oeVZm42sj1toDp+Naqg7kBSg/EwN8ql3tC+3A3q1Ynr8X7zxREQWDrUrYPq4lpez2mVDEGcN
BsWEv/OlGav1oik1gCCApPr9HvhBUNPdyiQSyt/1Kvq8qUs6kNVRgnH4QaQJ8pPPpEspV0q8jJ9F
9EHYYpt2Nh5lAGMQ4WQdvEA5szsslhM/TS49Xlqxps6FWAkHMshcrzEpPnPfiyyfEP7dMEJh97T/
c8bbvfvUx/A+yogsUPq4XVgiXhIUMUBUEacvBHbQo+MBXDBckCdEFaQyP4ffNE/0GODRN3ZHlL/5
lQawCUa8Lwd//v0IVTKQ2p6oK1DiJEVUhnioXaMNIP6aZsTXw/f89riJHHcE5at148VWN1f3UaQs
HjmbjXFK1pQFceBEXnWb81TJJF5qwM9GoG3qnevPPF1Bnj2ijQIaaHZ+EFHvB1VPoTNV+JFuc6uP
3ParQNmxZsGhQalsgbsFEHmmfVGpV97q9pBdKUumnrvvUlcazUeDgo8dgeJFpsdQkbI4N5AUBKeL
+TvznVaheXj2XfCfHa3q6KpHX8ZLG2VUb2sEVaJeRze19WF/daQxNvQI2IpjuUgKzFHFJXTIb0Xp
iXFRYMyviKJ5cYCr73KbYTPuwUAJgW3R27mqMO3jXPvPN1yg0jtYpnvYjKHd12yaZirMiAzfejuY
P+G7L2lfvyqBZMkpVtMBEsYIT3uMqhWhzK5MC0BFRAvfFECpzCBppspTDy8GtLugeWqSGS/MeY8O
10pXrFylugodWng4FxiGhAm7NR/R7DMeSlDOLVU1d1P4qBg4QRsLxUZgxD8+p+tNcnJ4qIoqVvhl
Z5l4pEZDXBWxPgbPRxN2WYDVOPuQo9HjSiBOPyVxt+0tTex2tApmGOa+lEKzloGRfzLJdLUsm31Y
9MQHii2osKgk2Wd6DeQt2PerqF1QC5Gtc7Lq1rWCOCGkYjoSqPfXB6SDVau6gugrAAdYxRhGW73W
G2R/CbSFEwElOhMjcfrEXhAGZCdco1aQnwlu/IHJYCX0PzB9nHzEE/dDhNPiEsrI9cFR40agvlhp
kZCsRLC8TzJwXENH0k5wAQ6GZ4Wn2XOTlrPGvcPOYPW3ozXOWAdlYaklIL/N9oTRiT1pFZwALdTd
AdgIkqDTFHFTna9sOIfGpDzBekrv8qdZ8NdIo4IA7XnUhCa1rLivOHNFKCQ02fppTS06W9iBXg+n
rNHFjRbGoEUiHJJWQy4lVzG6E8qIzYEBfbdGLUGctTwAu/N+CIO5e33JBdvoEzMYG9fnlIUh3rcu
Ndw3MwaFgtf55uCpZ0A5NqN1av5rpUqtdMQSl7nfJQ1YBKJpaNlcxd19keUotRT+3i+rDceJWARv
aODa1VvwAvOT0bd1GSMZJen7mHqrLNM61u8Ro0+5yhy/nxhPj68VLShYIRnl0xG45qGHJPTnaKjP
nSpwqlx2zc+fMo12EevPbAuVvNC+Y4DUjN0Pseru+3Yzt6qS53P4FHkO1Mzb7HEIyTQEj7wGY7R3
FChh6oAquwgpKxOHPKAby7RaXDIHoV0Ezv5jfQMjtWMjJgb4VVlml/ZjWaygeF5badsjhOMb81cf
2nFMeUGI6b9cQaGhmnxHruqJxNjI4XjJ9ewNBZFm8/qtQFsm2KvVWh7TTM9Ka/RKO8tJRPXayyyQ
PNbw1GIC86Of/+x4mtf/0vynEeG4tNJDVJOZqVZqYsNwfvTO5JnHGlix4cTyUNX+wze8J+BiaiBo
mv3YM71YzHwXWVDszShTphe8cUvavvWe21x5MpCnHcXxVyrB2RvLhOlkHwlkYXaDNiXVbQljHFFj
QIPCq+Nagz68mD2VU8CJh9nat0YKaUInfBFEsM3nKDlB/PVHYTdWeIXTnZ4DV3MPAtbnPVUuHQvW
cE5gVUgXWDfB0DVIzOSkLSKjU0TlaykbBeq2Xxywhp14YzwyOM7/O5BiSIXT72g0FSE45PtRecso
2/WYlM+ZfUO3FRqWhYX7xTcHvvlq0EQwQfgx55DgZwxFfjfvV3GkPDGYAmLN35bxQfCbDDphdaSP
jAFQhrHI2cCmWtIZZxHqgfKhxgxwsV/4nPaC5cjie516CbwFo7bU0S7dvuUp7jwLjp3I8lK3OVuQ
90JQfbDFMh6r1dGPi5HV6ma2QFLaQ5dh2rObWHeeyxAmPOW/rQxdiONeGOXUtwkpWWkNyz/YyN5v
AEEQYP5923cnbPdCI5MKvg2j2HBsG8pnQ1taC3uqyrf1TzBU1lhpUgo9pV6+7cwlHzO/vbcW2v/S
nP12R5/NNMZbT9fo80h2vjyQ4dF6Xvyr4uMUtG5f6wgdtNLN/HpuBsz7I48R288TQnuAbOdKj9nU
HypsFuh7DS8IuljcaGGcD+MYC1yNneRcEfOgi2UUcwoFRrgKgZzA/cUB8UOZW+92eMjiOMo4Abwe
q5orbCQqEHw/2UUN5LcQgwGIR5qmulg+5ogQP0y9Sngje3pJEagLYxZaV//4Moxmagaer6wc/qRG
UvOo/CUqul5k9YkxELNVfSKzUBG7rSfW1u3uc2scEUYZeWB/BIfQaYRN4xeiSHRZKDmMznY98Ma/
DcOZDKsJNVgXfAE69YDX5zOR6zEJyl3XEG+AUAg21Jcc95LBHmhZGDjHCb2NpGFqGGE78NRapeZX
IYPmly1Bo9x4KWJ4qbDdKXbwYk9/0IdRWbvcT2R8ItTnMGZwW7tI7S/iWjagirRKcM+j64RNuivm
UYC1aWmgqEMd9FArMpwJqTHCB59kpwvg08XnIqNKAnyElo4TuUBfOQNDCOhb1HJT8sLMxX3pZQWF
QaUKM9ydYBbZv+8jUDxqK1YtAtZaXSVVRPd3Qkz6OBLlY5FZYm1OHcu+4j8izI9lqcjxSF9kQPJ0
wiqWEsLY/VEVKsYSwOg8hbFTevy5QZsVO2T7PFlOEuwWiVNylhsR3pOvujo4EtzTuEV0DWWSPfPm
wUAhZiEk0ae/Tu4t5iSHxhMaSOAQe33gjXxHEqN3VmV4LHthhGxn97ZyPBkASlpBYJlLrMrZhq+c
PrtkhZcZXwOq6VKl5VO23Nb8mIxjNr8JVtIhvyGgSLIH/kvMZM8mBJxluCxRAYkbzUENQAzT8lLQ
LmCt8Gu+0snr1AL5c9nbw+Too9VeNm798FdLfATpjIg7EoRPWbc0fDZ/MeRMhnZ6Es0RtuJL1mLb
J8jrsnc7VqVitRUZMuiRp+njxW6sHszhwtACVNp2kqNgbqxZhqrDfVZ8GoQ+cfPPQvUeDE1R0CDQ
5/qJ/23wxX5EfQg4avi5N0s6EMcmvmSsTNLNGGc5aqvYvb31iSIhpe6RWzgOeQp4IFcNhojcOpeQ
8hm8Pg7ia6muR0YnBgiL9yyUMAG0G3onsnFjNIItOIzdIkYJNzXGobf1BZHkGQmGoIIoafQewNzS
bdx7nyMQqO25bPYxnLVsQ6gs29yYFTYx2J/v3jxmTY7u8Lca3TsNazc8AoSA3v+NgYoC1FKMHcq5
SJLKkL+KRehxTgK1lLkstppMdFq2p0TQ2EdQ2V/Sf6bCDsJqLxzQ1JZNJjDPt7I13n7PT4uU9sm2
hoLpRmkij3z3vw8OYmEybzfJzr7iUDMrNaGXaJHgyAyQ30iT8V+x1AdyU9fZefOMDBME2JdjbOW2
hamC3LRAuDNHuzijCmoPsqMsXdgmqMMgdKH0fI3O6JI7+sxkVqF6K1kZ92ypa1Mcxh49Xeu0ZL2p
lgAtBZ+EklQH0CQ60VEph6P/Tn6ebG0c3LNSFzwHW7ZRS11xdi3tGMFOaHcEkEI2v1AxeqVDdyhQ
+nb3PSYPTft0ItozEfBIru5HEUDiqP7U+29O5mtaxLefcRTghPyikkaJg2jXduBoy84/vu9CPOPg
2GYhQf62vFu1GGEql5/nuQndic9TPXSrCC/YTfA26L17olupVi7V1H0CaqiPclAhYnXr/tw1iqoX
dOrzYyMrM9JiWCcY1jK1WV41JAx+YiPi7UKk1mZOMDmCivQ9kQOGLw3q+JYZgUfVVC/SBoMh/CNA
96Li6X/3LnOYdjsqJI7j98lSPvDFHfqppDt0dZxiqhmRBySz23gEMFJlz22JlsGgYHKhNeBEMJHL
MWs7T0xdUEEY/gSiKFt1wXBR7TUH8QgdGhwxqjSc7xKRyGJT189v0N+B9d0jAR/d6Zg93GXiuxAF
cZL7JeHmoLAg+jYzGAhVCaAeMN/8GMCMsNUqpc70+x6pg7QMWDD6OZwta9EN7XQSic+VFvPf8HAn
qjQJdv7a9BqGSPrGzuUJHE6rbYPn0ejFrQMYsL6qT6rm++2nthayQ6nus88fJCXSrWTquEvzsB3k
ZcX/AFBo0dgIPl3SGF3k39MxSuw1W1FbReE6+9tQ1k/rBnRxKPm5p4QtvsV1vpzY+a1Uiml28Zra
uljIO9DuiQMsYONMto31imYd+KhIAxgk2MFA6RCflMYZwxIYE+IxmzjDqflMZghW/B29GYXl5c98
8byf2cBGB7K0GfVKHZBfFh/8pZTc6a7VsfnqGqFVHMfGnqA/xOxh8A5ARQ76jFeyRfASN649Txb7
v5DTbpkmrFppocxHP/scpGwdFi4b+J+erk6Cbp13sNFmsM6FilyVgzSzjnNWdd7WTf1UmAKCOwTA
tJ9ujiHEonRP22DHxv4wqP5GxYmNFgz5O2poC+2LGIoK3Su7FT8LO+91ZKffMBnBH8gcAAV8tiGX
hbOdlhADGn3N1O9O08Dc4FGceeTbBN6rvGCgMtHpbW2kpXvHelYSIAyBTHJ0aQq9PRRzQmBMeywF
1p2aqa0zuiEBly4/wrqYlQWl29tTjLD/9ZN4gSdbfAP7lNxbizMnvCBX2/VxFJSphoe2bQmMN4Kd
H7Jca0gICGOOCCN/S2sBtYMC5WrSvDIOV2PiKpRYGbcHHaPr1JxcGUsguNxvR8BCMgzp0n0kdvyD
xEHZ7EXqRaKQPjwJIbtcHWWn5n1aVgHYM5U51807iwpgQZdpk8CDIDsOCMBV9X9/Rm0NmZXdi1Ty
HMc2HlAxJacZrBO18wiutGqoGvK/lSVqOrYC//5q+gPihGPwjsaFlK77gJi9aqfGFP1feHGMYdMO
ojtHw9nS+10h7tInDI3lvDCBg1vclov4e5OQcsRC970pKMeUQepln78hxU3uoxs/56sfu16WHbOQ
RjFzNOCIg62xnydL1dWCI+h+UJuPAgiSvnLhgC0AQp03AqqJPx/TK52cmCDRcmPKZ9l+yxQmxTiE
8IyYFd7timZIDGCfJLTtK02PymRFOEiLy0MXMx96/0U4qpGrES9SPMr5D2M+RucgnMhvGBDR7fom
Bnn/vmLJwJ1pEOEmwpaCSM8sFan2DRTQgf3iute2etH/pHqR+LToZcRiuUEL6Nr9i7UeN9Nb+RIf
Rk5K/3okQrbX9STyoqN7dAnEqOg819OKxBGHjdJhbmNGIfbNnAsmbFMNHsKblEOmcgtjVJleix3V
tTze2XvVMUA9DvuUOJ7zB+mO0XAcjZIdgu5SnG8DbCuh4MCV96kra+RHFR377dVKTR2WlgrOuwmZ
9eVnbZ0K6NSohA6jIx/HfejAPGmtp6qYXHsCtIXz8VN/kQQmh7qTM1BIj0WB5mQXtbHiT2g8Birs
ZzzcnUM4mfvJxTd7JuaiMWKzSvtEYywJT/s0deeQdUphfyPbav5UlEtYR8IqgD7sJKURT7Mo1v+u
1IjHQU+fwzEwb6e2XEiEYzeuRGD0XT4vjp/tdQnKWffoLqlwhhirB4d8nYIt3//PjJvuxMSFw1ap
jrw6HLVVUvZN/OTlv76WsqAF700Max5aKXaC7H+7zoXUgsbFujXBuq/mzAHj8Pd6zcIK7WK4gs0S
K6rt7wHJq02vqPP1VggifdqMiFp2UeRsLGGlcKyIDttBLaAkeFOYNe77mvE7p2N4mieKdRTzeew8
xCtDxrzASg1FPt6HwEaiqPiTPwEO5Z+0Wde2o7mxpbf9TMgrKNjr4Jiyctuaca5WmvjeMXDNPtTT
klbUAVrlOETHyZqpmri9yMDhp3NWJad4L7v5/ifSHVsru5TjOgj7YIZ5tNqZgx6IQ/DGpnofWfRw
X5wEJ5i11r/jVDKcnBz2KFitPAbcIlKysekFPtyw8aHvsr/fG/Lu7hWudeeST/YOajjXmJqgqN3n
jmcH9dlJ9vGt++3vlYLL4mQiD3QmhlDwLx7v2YJfr60cCRxfsYQlLqN7SHIyo6eGrHH6BZDReBGp
S+mEL15dEGJ4OEmgLJs/SRmSADeTLk/AHhGKjH9GJXcu9+EPG5Kbx5ElkmA8bWPmrjgmBafVnd1p
cm5WVdm3sX38yMRSKPw7BIU4WXa661WzzAtbnULC2A8qOCwPbiS4A9AehL3BxFRoL9eBomvQUVr8
h9VXIIG9Nj+jcf01PBOiKIq7weCisCmkypeez75/lim+KcpW2GqladSMoisN0aYE45Zhhbi0Z22k
cGj+mWUxuHUAIpXvVZTJAf1/E7hHYGMtEH1skOGONMjTkqylhTGAp+Ba/mCU3HFTxHXnR5Et6g0H
zzSEOWLBxLY0btmWLBhxc142p8EBcAUPqYYGWxFg6ykmRJjEMRA6OwfxetiPEeNI1MjM8BxqcthI
KWHqHx3CeHCxLcJzBls8mPtA/FV/WnMohXyJjERO2fgWyTC6ccRyUPPqTarAvYuAqoECghq2RyEk
s+LGUH+uK66d9BLUZlp+SEZoq53w/ru6HJg3aQcutzoLKhkTU6ZzWXYfkenUvGJ8RMwKMtaKuKPi
XXpujtW2WyJR2q1LrxA5aIOWWXa5vHYeLHsAzz9eMVhaaFl/U8hi+ZXyJdTpLw9k0tF3uBmERekf
oE6CAeEwLdELDMhDlJtvk34eUdWx3x0teWXLjIqZZHNQPV5ggjT9eXguJHofrD7+ea++2H4l4Bv3
oUFfU7DbHPNFasuVBF88tSM7ulCdlHeL79O+MHB7jQv9xgQjONgqnfOCBlmvRQnfjxOI5LFBw4ti
pnf/gklEJuO6mlbi9UPydusj4F/mHDYIgJSwexLOo2iwEaaOzRmTW0OL/WRvt+HLU+Kz8XkNH5G6
D3IE+oYKCi4gtBXi9Dok7/N6+immoXPDxwFv7RoTx+gutqYlA8Q7SQ8Rw00FgNmFDhKEJEd0mrC7
xUlTGZM8P5buIxqKyQtj8IezaIYemvjGzi9jc0BiRJaBKiLz0YmPJYsaD0z0B8eurvuo/b5pPMR4
Hk2Yr/W7oFaey6N0QXFCBcOnitkDC/EW1bWqZiIs7bxEse5xsbbPEHtAZ1XBaI/T5fo1N+BDliqg
9rb4OhNOJr5i3EDOxtfjSafECSMfv8hplWzT0CLBs31fBQXT/xPIKXlVKf0pmjzVCyla6xA2e60Q
83YtRZGWQNqx2RmzIRryk+GGTjeG/4omyKr0wXOIbRP6daeNHgriNne76SkZ7iOFTZA2KYM0YkdL
IVeaLS2qf2kHW0j95AF9+RDPrvTpCDHEaC+cfIdcWolTSlS1EaWCtonGcaFLBJ5aYCTw4DaTu6pP
CPry+GogYwNaFKhCGCJ82mj095iei0cHWx/E2sXh0ZLPEM6QafwqqQfyp0vVYzrwsSlOfx3OwplL
Dvg926bLFrbVA9PU3hV51tWUF6f8rC2GcTRz1Qv8Gl8wfekEG1s09C27ho5R6TRhQe1wDrW9Jm5s
YJEpc/7hc+8LFNrciVbFQ7zOZGxu8uUh1jt2xcm7g+X9xR3GiyfYZovmYKAdUEKKmxCztcwGk4GI
MRA4z00rr16RaiR6fUhMydyLKQluLeQXcf4jiOdp5vD/qkvl+f+WqGOd3twT9Nz5ey2R81EL3M5Y
krdvvCTgvvjkJwHTPB83bd4cstnPv4MS00i55Ai29EQZM3wo2T4GrwWS1fXRC7rPjLDMF3jF/dBe
THUqSv1Wj9XK75/RvQSy4zhDwyMq/6JnIx1HZAWFmYjJ6x30kbVEUHkOrbDAXLURkYq3tlosCKNX
9ysKQeGnz0794B/hhxuRlKuqXQM6Y7cECNmjdNQG/CiF/eGN6sLuyu565ZebQAxZlFFY9C/7cKys
+aBS2nUAnaRdAdPa9613ZZEsU96eU5KLuI3hCmrN6kjNXh8gylgrNvzx/VUUSVmds+i0FQ+uUda5
/ggpyW8Mr8RZgatDXvKIgs+hKrcOQCmvnu/a5yo7kaW2+LUNzkGh30KsjZ9/RKkbkvBncYk0GbJ7
zpSZl5VhTwq433q+t+XPHokZQHqzbkVHU3SSKKPoMYIvU+fOoh7Thqx037xg1xVs32ZPHwr2udiP
m3zUjQA7l0AmiKf9gg25VfJWG3LRtFJpu1rZEHDa9g8CRlzM+c9YBv5iYYLyf5ZRdB+8587rB01N
hPl+l4kyNjrtfqNtOhj32/sAzDKCbHy+tIUeLGEGNh2gRl+OOXWPQJZwpWjMGrpHMhRSXfRrC2Or
Ga7P3iDVRZh0XTAbibD6h4kdT/t9Ribmv1pFDNoNS3BYog+iGPlVeaNr7fgmz0Eja2bYAdbmAhRC
WyHBMIET6bvc83qNyU1v0KURyTaAjDzrBHSeWLClbP+iRmbtZ4NHUsOue92SKhiW9BDex50kX5OC
3STTNE0TbXNQ+l20tZV5C164R4o5xVGHyZDFtjg9CYE9sncCDXpHJIsWk+pQZC5P4brd9i6d6gPQ
qwef3a4wdazx62h6tZnQvEB4TAsS6JuG3wqcOZYxd+D9ClN/NfeTMX9lcgkequ9AYN6dC1SeFb09
kksDhRatKTTjxRnzot0QFn/oqLAQldtTtSypfMUxsO5y+bhZbnpBrWJ2Ct97bKwf7c0bxku1X+25
xvn8bqjKYV2oeKjnAZSDhq99UMfGSCll3iSZnwj+rFwgDN2MaE9jJ76yaAytbZl9j/DYxmM9MnKr
PzFElV1z6n0e5NU4IMlXkvJAHZsRLa3lbTIzQu8xSnrE3a4KT4qjZAHT+/sNmjtboIE8f5x0hQal
C24HnijifnzcGPYZjSUJdlw15Nfz1qJn/SQQFekHN9jyODBlgKIDCAZWaTbBDpoyZfBcBbB8wEPS
hKZE9k6oPrSLgmpAJ9UrbgiGSGhQiJAmr2pGtRhICuN8Y/XT81YRTM3EZwV4MK2TiC35b8Y89g8S
o85EViZ+FL+FEBnDZAIRPxtFaOr9MVbfLvoh59WCNZw3MDwi352aFFtYLLoOc+7PQa4JVVStCZuQ
KKWzdS+Lo/Pk7O6mhPxDIlSpzDsdKAZU38lHWpOk35dcr7lIMtj8FXRjMoB/2VUJd47VBe1JLK61
3rpYNJ11eTP8LC68qXLskRwSH2GwRINQ4AHkZ6znb0RdQzV9L6X1kZSW1q3Hz9uhLKpi9sSlXss0
2oX476fV2dN9AMOtJWiB357pJDkr12CMnCz3PDd8Bsq/QuY5Ncjvdg4EpYNpSSFzW1+gTX/BUglB
eYsnItNr6SJvca0SaoUtQdtwh/IPBjNkf1Srmro2IjqE8mEbXMXNjXR5ppOmHZNsTd7jDj3kGkwr
Q8gOzWTiD0yJTl7RaL/JJXms9uejCkG2M0/+VAOAqkZbR3ZRD+Al6kUWcoobjsqPdMVXjDAftrBU
d4tAL9Mul/HA+ruNr+Up+TMwp5hcxwO4oJ4+4Dn20t2Lo85cu6UFT6LvdTnMBta8Tdby5bx+jEjd
EWrnSvW6ph5S8jCLfUQR31+yIakXGZwtR8wLvSyjIeM6t0psAISmEzODZcXTBL5iqjSBx6v4cTQ1
uaoNVsFpc8Yn0og0lJj4I/CJrGcqFxvoqkeKksOR9ptwUvCjuq6wEZ8sE/YvZAVbl5jyX65oURcQ
pW3sL9zI2qfTiAhDGuHb1ub2tvUv53vtc/5ndK7vCmZHmFlZLIP0/wPscDCqts5AgHNLX06m8ujY
4rBnBcC+MRskTXpYJYiBkiu0Pp8kzZQGeCxX9gWz2Tky/QvcouKFQjktbC3udyQcCtxpjJitcRSb
q+dfXq3oe8u7x4VVEoDWBed0ZcK7ko/zxJChqqonpKoReBGkmRYe4gp6Bp6Y0hxZxey0k48HoDyz
IJn/qPsb709oFgM48E3tplKde6+nqxC+4r7/Yl9tSOopMXGLYYRYnAMvhqwcfATek/X/K16FJiPG
HRiI8tl69Q0UJbT6QmH2onGrjPBHiRYdcEIvDbYjDU2s+/Xurn1a2BCtRgABrMeMlpRLb+8mdDLd
z2XyGaIhHoO8dmLuEgkjWCH6dr//+CyO7zdddlJJikz+eIVOEEZtY3pEtInAzILKeiOA+P+p86xc
YobtNp9xbQHkII64icjbsSgA5IE8D1GV4uXTtjm7zUGWwkLgCz5HLcZExEXZkzKuMazCujSALWpD
aAPuFlyRpe1yjdlBVHnvvRtI5c/6lmwWLoObgeo8tKngajhaWxF2TiUY8UPA7vYSeiQBiRwtt43T
mhwD+kwr25OTUWr499v9HYhrgVIh54PaOdqYD2MrgqoSf2u3ynTfr6BgWtZuap1qAVRfMAS4Ibm7
8JEIlDr7izKOdz1ffHcSdDgNFLCAoNMiFhcJYc+MZZ1jwi1YZm7lX2HiKietmkjCvPcVyZ/PuBMv
ijkN4D3jNXun8lHkkDlxmxyWjuxTMFbYT6wQkh9xQKn4JdqhRga9FW0/9aZsyTqvO+YgRDc+Qn6o
6v5gnJOgEtBb54S7WrcvbqOoXHxy/RjF33zqSCLxp66DxVA9+I2wtidERk+Sw2/wZGEGir3sEI3S
lJEBx/6FMxqW5XjO7c3obyj61o3dpubRnhqYVOMwsglGOe/N0uYcfIaizmmoLAsi5dLmq0LHl+sS
MvUw12UD7CqxGBXTB3ZU2C2ZLPK+0YPIMZAtwnWcFDxOp0MATQ7zPfEp4DbpbYR3grF1H4jjuzzz
gd38OTL0mPF6aEAgAhbXMxAy24U6t1s+6f7B808QIA1Blpk9b2wRweopQxdBommCOk9GC8RkuB9G
l/BiqPlxNLcfrDnlhrq2YE/qWjSu/etWn7cEYsrpJfAK+RQc7T7PVMkCCJ+1gVcaeS/BqsWu4fmM
OEYHUIAV2TtYIXLBYztCzBFmFntwQcb9bvULFSwAFxODNJg3JTh3EE3xbqhTe3kVPSqSL6rpmUv5
WyYOgsjfodYQ5T6QtOthk8J0MaYhMQSvIEhhrDv8P9eoWJxx9JQ9l72e7p/lPQvs70L8Q6fIjgaB
tkq82sFaUnBzdl+o7M5f5G0BoeBggPPAoTVx7+NIeVYP+SLZpUV0J4Q+iPtaX+6LoD6utQPFrUeQ
K1GNOqcNPcy6Cl+i6R8tTlRJ0QHUqxc9dntWRK/EADkP9S/9IWoJgYvqe/DXzDuzRjJylVZBuWhd
MuUeXZtNIYZAEYFGgSg448nohItr8wK7MKmh8vbK/AdeVjmyfm1yHDgA6EZgtWi24/84I41Dtfe9
WwLB06+Qw7ILUrFKYQZVdKeDeG25WHbESVKnPv0J4j95UPSrTUFEqH1aEGqnyvoU0CbEP54A5UhL
ikRUQFVpKuyOrCBi6ULU+2Qq+Qa6b4XfL2GkSYjU2sodjehhFMxeIBSSMu4ooX9Q/ZLD2cFDhrls
pfORRSCE6nOfTG7kzaAcWEmDXQXtxVCv2li/ndyihsH9wENy8CWSOwzT3n6pz0rz8hfiN+FQgRw8
GXykSizZfTh1levosr9aiBF1SdcXCBEAKAK6FmFnh0GTFIYCOuA8fGCkQMuzXu28PM/KlHenHkPC
AmOuMHmgEfN8edM4rAPKRj3VswABfRCD5OfHyV42GzBd+odPVJtdTLQxj5y5KhYlS1mR1RGL1AuR
eiTU5ZviNuxazmRiFxuj9NtVPlEftoLDMWwngQsNxeOKmnIGwDb5sWLGJS2n8rY07dLTbiNkmTcK
VJSctEv7ZIVB6Ef9IE2i6DECeA9vwX4JlVY12wGZOnbTYYZDxmjVBuUkIYsh3WQV0l5iaZq0s1S1
J097fnF6l+dwlc+44XNNYSOpOKtJmkKtDfKpdfdJFs6FtSYjY2o4x+rOOyaC+iRZPmvsRfhohUjZ
5RtyoO5/015aXu4BpoToVbRNusTeBhxd0Y+N8uH3H2xLrPe7nb3t60X4AvtNzGD3pomQWkyX/DFf
979KE+8XPemUU4GQHPQzP20xNVkP3DbsE50FnTv/NQgrD9ELagWUxWlFi7xnSeGquvyy5tuAVoPJ
iZA+lZkLhKaXoT4vrafiDOqtSTmh3WhkcPxvtvij8fwVQ4kDqhUEY6hl1RmDGcPgsRJiUpPNZFxv
ar2I2Bk0DhZ77AQiyu67GPnz7uLeSVzBd+qoruXZnMpFSvmkFq6+fledxs8LA1nORdVjX+uA/3ae
3GpANx4uQG4Le83mgXQFS73vlCjEiuq6ROq2nPY7W/xHjrU+Rf/I2NqQHvXK+lmHL9n1V6Jhb2n1
+ILMkb2r5AWQoZwHU8j2lmGtZ+yHqMufdCww933GElPezBEcbEHw8Bmd3Rp5HC/7BIHx1AOVlvUQ
CIRKwXnT5c2czBQWE6GNDPkzv3QrglcxVUnLX3ZER8P2JeMCbqOkhje4vM3ufVSq1V/n+UerOI0b
ZWlbgmKTtVE8DDYChAnkq9Y9sCsGR1ptzErIrcdfApNdHI9IBBVxrY1ldXYex8SeQgOqmJGhIyGa
nGJdyG49pUjtwaySIaA99eBsaJVRm6+BpEtcgtEVwC/oXfWfQqPQlD8fVpFs9+sBuQf3LCMH12qs
M6J31/MSQOtzNRlu2gRhHtsQULKZ6ltbw9M8cmrgw8dvr2+HRDUrA3TDMIMhZu/HEmJW68nD9A02
zcFgPUxwef42cVGFqWsxkAkrtYzE8o9PDj+FaJMc14sKIekBbsnzDPLtIN8wEwtvCqQRy30Gnift
JzhShDNeb/4fP2/e8k5Trg5d56pNTB54mquIzVVkuXWaJroMUTg0N92b75qGgYCDkTlS3o9oolfs
qCjNjzyI9btFU9Q9Is6UroMtqwyZZeY/Llf3FGwnxJkrKNrTvkIb7FPo625jPHshHSBTi+hbBxxa
SBzEFyP5OaZTe0Pn0gmoIlEOgaqQB2ZD16i7+xwezvSakXMhkoTafbeOMTCTlCs1/0R7Tgmhvi6J
iJXEg/M1j7UsbOrljX1Rhcph160xXTSfhdaw9AJW4HQcK8eigTRQUNEgLzOe3Ud5h0QVpQunrJLE
37IkiHB1PCtNNyMPi1YRAJ7am2qkT1ihlJgXoxSKVV7ecJXqmkS/4WHzOM2tiWihwFI4XovToz4v
kuFzbjSrKV09LmJUM4fgBSiYR9u68PzNknqN/QxCT/rhoeQVSIowDHWCGf3Yfc4Gw5gbvlmwJBU3
Qow/LgoDwb6WQmdA8OI0uORLV4nh6mn9/nnN2mZ4iOxVgcbMmJy7a6OeV/AWlDmlhENsx0TNjzuA
o9kXSWaprHC0u2KmG63JLMlyMOqi6BM75E5OZ1S+1wbC+E8mJKWO/wdXHyCbs+YJB3SrQYMN16qU
Fes77YcH3IwsuT1cQcWWPcv3r7xht6sTkbwvCDUFwx5Y5rEgwV2LZAlNOb1gpN+KLRVK2KCteP06
z5BrHsmZmBXhv1/z0SyHKsghHI23BcTNmSxpO+MKrk+R0AnstMUem1dKs0mmqZ85efOHEwaeHwcf
fPCO5p9CrrXalHgxvJi7Mm6TE/gD26UZ73PrVv80AOlx/0yiFCNZ8AFtWvX1biHf8+4hR0qh8YmA
miTRYQ21C4/icWTxwllz3mDQ0ObRGAmRgjCEnyNnpuStjvqjKqDKUp7TTVhLJlrLeutZEhuFAWi6
ZEKh0QJPSHznYrPOM0ryfS94D/dyTbRb7NzO5zdQaEz4Kai/SfXwTfOnbfWcegKrhtmFSP0eBdRl
iPyZ7zR2krTIIGMhthz1P7cyG9lIVj2+JlDtFjJQKr4m9arvJ+tvuWcF/hmXLIE9gmaiYLBIoGlK
DXwZD7NKUPSIO8nAKq4TQEwCaHO0dk4I0yq4baejmBfLexClzYMGSKVHdCTxf5JHEYCT9WvEFXR8
UV96ZKydPSab6lOc+HYZxmILeHM8Qf9NUuy+em699Gr1njosdG24nwCXKnBNxqqfwuwapMsoMkvk
WLMNGmMFpWSLVlr4j0OOlD34Jks6r3k+BHY63Yk6E9ub3xOGTHjAExpmNSVDhLnQBAfQpulCqTu/
/0J46RPu+snA3yLZcx4zzi573HMaDppbhGvRQ0xrO/uwrmlr+TvTTPsySXrRqXHV0AbBPQniAAkA
wS3dHPiF+c+CXFAhtrSi1Z1lT7L3D2AP9GMLn0bnmzw6QFpVtN+JoYSyhDRQ3bARfEoPQ4XoAglh
h1tQGEZJ8q7Z5M1LEv1zZV+0Wxdic19ELjL7Q8NWtYk+QjINqtzMYx2DwzSl3vIiph7d+oBNKRJH
PHxjTcZ87SUsyat1AqSIgT6D1ufT+OgetCjlB7d4JkXgk1WiSqyJf7WVVSLE3FSOjshQC0Q4LtNU
ExnJGjF4aTIyETqWU61DORiuPpzEMtHS92DFvUZ3u4YRND30zLNzMIPSGCVsgMrcVlh/7uPhW4aU
bumzylQNIlu+ULxXlYGG+CqFxWb6K//F5EJGKH39YCGXy7rYQwvkYrGqtHeD8y02wJPg46QDD4/5
bWnWsHUGzeJIj6vgQQhuJThcFfv8xY+oUJZUUzt3K9ezJgfI2sHxZ78/Kt6kZQvDG+E5SwfkCc6L
qL59TYmReBKXrWYxwy8ODdp2McbcbQXqpZrG/smEjxwAre6o6m3IGI3rRo3pCDeGoWTfXxnqy6Ji
IB1GBKpMfBeslwIt9shzPtAHX6vQWa0UbYulldbD54nN9gsEQ0mTG+n3PqFIsMw3ZMm7UsS/fdPC
vbjxJr+tTkGGWPsOFWxPjRqW/i+qePqcc1uraYt0Un4MJrnXhmSMY1bU0/W4m1WEJYrJqKcgLmKm
hRVqTTcTFql6sT/H3GSaxP6O27sElQw/155gvjmYu+SzVwaV+a7uBHq36I/Rduqf2XmLu3nZm7h7
s4kFimPyVu8HOXdCu0BeBW6m08scWVGeVhx4td2dhuoAsECSUncCHXZmBga0TDc9X+t0+hPqfbmL
Ch+7Im+JJ1QB7HRnFMOSepnyx1HMcrIinqWNstZ+1QRwCGpXgQsBPF5uxExV74opynqizZl+xcj8
p9CkV5x+a9WSB4hBzEavK/su0fIT0CUw9TzPWyGuSf5EAAH2e6Rm5FRVy9xY/WicbT8no7pEdVsq
UafQyiYVApFB//eJGBvhd5NO55MMJ8/iDA5DoVblRZcGvREEKPWEY3/87qAm7NdQ/VKYX6ZueFOb
iHIQxU5FhOBWIZ3eZ90or+KUlMzlgEBFXe+w8RGDXKvPH5oA6xx28t3EYa/R4HiG4J5enccgk2RV
QMLX0SO33Dp/zRlmKhbwZujLB1WBajjXwxVKrCq/bOOdJ2P6CBCW7+PnUV6ZW3jXptYJtw/2KUZW
1b4es546IsZfQ4xtaB+y1nE4VBj7A8tez+SdRw97U6tchJUwyFdNS3sActcmjYmuc9pepSfbZfng
D6RyeIaNedgY2M4XXhBFiNqWlTSnoJFhw9pkfZ3DQDWI+h9rJXM+TZ921qVy138CUHXZroITi5Fa
+kv9rFbr6reTdLB9E136pQHxUT034CVweMG8SjuOZjDGvT6xckZx5k9xrJMsgqJIGRgLzT20mErs
R8i+5hojDVYYbWOqrB6DXu9i5QhA3b/Z+Dhcyr6kXKbfaZVI+GWAWP2xRItkrq7im+DJwAQyRRW4
pNi7zTEmVQ1qGO5E3w09PlPkvKttYFnydhqn0M2kEAaOxuuHqKTonj9CLWGwDCORYOpj65fy62iV
4GYkklKEJ16wkhaW1rDc4nWvchdtph1yc683qYCFF5Jvg3A1cyaab3ygXo3Z2pNNL2uY9pMvmaT1
9bN0+8+6G/0DembWy5wi8kWoc/3B+DOBI3O6t4biiwfCSk3WSQscazCNIrNdH4CaWAurALMlTqoL
hPLsDRukZ4ez5j4KCBuPmoX+Du8IIuDxHOKq4X4WpGbYELGdQNNrQjRVfxhQFkhCW4e+ruRFwHnp
qcmds64YH3l1h4LLufsebC7Lc/HdjVMcBcd5Gz3alLY/CN/uEd96sKCMBvhu/BHzNDO6Q1y+eJBv
r5zdZBFiamuDr3a8n/0+iyIEmSexnnixN1v7nSBaetIUTYMGCDpnP0q/D1WVh8VcZDMGkLnEY7lh
9x+9bhVskZ3KUdRfx8zvCYByDJXnaLZax1RthLS4euROsPGvY+kOBCrHlqRYcFhZgcU4VNFPhMJF
8LOS2fD37mAgkVj7MtADRZfBWCEK8xZPUdPSoLmPfRyRmSCwnHl0XqnCerIw8Uf45rv8iY5zM9ar
fyyp24UBhTozVZ1zomI44+kLz215/x06DGHJGqV13YDVZ0iLtYM+Wy2kiscvauJ8CQ9HEfCF8cn9
fQW5fu4dutjdlh6FQbrIt2I1yCVyaY2eA/szDLnZJHoD/G7yQK4iefwXzdp3rcz13z0A6texnhzO
jugp9HOcyL7vVf69CO0DGsOoVHoJ3wZjI2xsSEminIMNRWly0J2EJxZ230XO2QdY6+KwVqvre+rI
FDIS2PGvuP7zIu5Q0otQNI+lOmeqhJMALxaYQray/hGOnekw5w2VxL7uDg+Aj9DbFH6DM03z782A
Iyy1ewLB0kLPq7qraOtUBMFunIvfZjRw0mB+V1B3c5W/s4Q9gvzxC6FU4bxQQm9CQBf6V0n6+9o8
wa9m8VYjOPWRQ3TwYcoJ8Q8uMp0A8gol+HTwRe5S771dgjITRt3cOu9wPSzHMZE+5DbxpOfKVtfH
DwWnp6i88TzHl6LHFrxGQ039NSz0sqU8SNvmYjXmSLXMdfw6ccHZNbTnSwLJWpytk9sf30GIP2Sc
ST8IxeUQAPNJCsrj0Tpoy/1L4/ddF86+d05UIPcC9GU07/IcHPGvIC9AQPMd1bqtwZhylV60KiRL
CyORlYUfWhoG6a8QfOMcM5NuNnkTFYYetJGVXlbx6b0i6QIriONLHE1NS8epF9/80fck7nyNyCrc
4BS28pvzkLpmSbyZAR2kfh1vIBu3z2m1/s2GAuITUlc0lDKZtIVJ3t3T7VAr1WVkxx0fF3R2ZEtg
m3kJ+Nd7szcbucMBNU4fpeNgXnrAi3YYmZppqimaGnbOCDgUxr9w3VOnXcUB1+WGQoqYtlByhoNq
RzXE/Ef3YAH1sc5JAPPmpfX9lbP92vspaoC76+mj1ea4y1pgRKZOYeL+ToJ0Ei9g39mPFnG78jCf
nWu52QuXo7/n7wB2dyE3j/X1qZpbPWpv78pZ4sc3EURyBDUZCZTZ8zksaLZBAfqoLyKCaXDbVi7+
q5E8NSYIQKFJdrqYIwkbP4T0nvC44Fgft1bOTUPPp6zg9L72saRTzc7gkg9quxKvRgK5PNvTdzSd
oeiEXASTOghtHRbS0yqCESEowZgh4KYmn+djLrRPpxl1v1keGL2EjcQe3f+QtiwaIkxzDYF2Fndw
n8AZDAz/2BCP/i3col9WTX/J0FrsUKa7yatz8146gNiJgQuboHvdvGpEHPBWql5+H655y6L1L7Q6
1cIBWE0vmhugsX6bVvzf7WydJMHOQENDgUT+tCSHfI5poo9hCWhueTBzGOqjdEI8bkfJQYFD5paW
Co9kuebNp8RvyP45sVm6fAH20qN13gTP7H1VADu2VK2y2F2U80qFSDs5Bgvh4DDRv/cSUpSRfPRJ
Ka+WvnmvjsFQtIE1savlOdsv1nbRnWyhx3bjo5H8pM60pMc0HpVm0uneTadThNaePJLnLlm70MN4
4h4/72OtJSqI9/xLjinL8SJYw2sGKZgBsgHWSoQ+/WIDvTOgc0RyDwfkVCgnD4uu3N28DzoV5QS4
LaamUTfbydLBOOPT/+x1cq2sCQSYlXuGbSf5ZcxwP0kAdNZRwuYGEw+WdblEo0RdGO454xCkPdXg
ZZv3aEIy18DImsONeOI+nye1GTqum4wAyxMO6uZ5M9uA1LyqBXT0tN+erGPqCf9T1tm2jvu+mrHS
RD+Yh1ZFPRVgfUw6OT1tpqEmqL+JoC+LZLDk7f4jm1RveAcr1D/iUDML1TPbdZBn1Tp8sL2ev7wf
X2tUqdyd/UZybD2JQvSuq2Ygxt7rrWbm/2HUaFyd9ZW9XbtL59wBwFcDVNxaLQ4UE6tIfUmzS394
YTOkHRKzrRhyiQQ8nxyY1zCub5VcbjclaWAI2ZQnvikXCW5YqBu6Eccf2zixn4802eVCHUuBVLw1
2crzqc5tvIrMrHw4fUEgMtfpnpIbk9fbQ42vpgu/gPHHWZ+3H56xuSiBbF2j3i39K7/SpjWBzl8n
prtXiPOhfpQ5i5ndsMWcLYzp0KXGHnFhKxFJRbhIgqZo7xE6YfS2NmSiWSL5w7wXFYqH/CkWw2E7
RUO0ZxIozGmg2aJetW0rERJe6IwFl0eT9S9/BsAV6tLLR1N0JkAwS6x8FhprP3i6s51mHRHednJG
4w9s8E9aD6FlO1EsJEBA/F+ant8tFS5YOMzGo8GNhvMfO8fP4tEPgLsqpZMwEfvbyITfRL5afice
Dvbzd8B/He/lWoFg862rcEdu5/8mSUB8iJpqsAlsiPkao2tePwmZg+vZnJrE5m/05hICWa+iLKwa
+6VowRX4X9T8D0knRytDlIUiS4xBHDSzC2w0ACX4JRfpGkULLDtbVEYXs/prr1QQiqqy4PsQBlUU
ulJf2EDGtWoERiaB4Peo3vTMq+adWID59a17iTOCjO6dZRtDMtIkjbiNHRr/LMB7DzSgrFd++zQk
buym38XPnI1/ft+ZewxjA3zbQgxGf9wnrdEjdVANLyEWafs41kcZ+0RvvMq4oRt+Ha8X80eUzEi5
3ECVEqB3u77GcfhUWYkxo9ejbWuTZuH90gr1LC9ABZq4B5Gsipt17tHN+6Zc5FyllaR3LVGanrBp
49QN1GdOwOXc+ykxLFlwNBBupviNLmqJdYm6IDXHq6Hhr4wiTmksrvp+BBU/t+f7uLJGI6cMxgj5
VKg7FfPmF6fZ0r0d6RTagr2ch0SzV0Y41zG3kAsEIKSHNKDAkRXspprC3iSJHua9fSFIydTQgbxF
5nwXLoyp2QXYKFdfXkiG8qaQN5FPll36AEa3H0xeZJq/d4QvDZUjJtiHsDfovIOcl+LovByGsazU
2WAysVYJNQebWjm/qW6uf6j2OCourYKhVpJ1wxmkglGIHRB1/D/1+xh37fVJ7b86/T4Zryzb/FGJ
gHifSyT3jZFJb0YLyxIuYftn0T/xmClRt1diGqnBQ+eTmpMwEqEomlHJuWdhBcWgno/dex+1FAqE
p/8bGIMwEmjHJAMnRu7ejg/47yosQGi1v8HaoNjWSd5R2NPpZdCSMjnoZL9KGt9+/+1bkeu5c8u7
fqCHyjoMI3GraLcwDuGBT7m6J7f81tgUAVbhWW4ibYxZKwOXmNHwHaiWuqC8xgaNSLq9QkwmzxZX
vCFPc45oAbpv/33DHealnNWhUciMobSsQWcZaCx5YgTSv0Y6zEl3SgmGMFyLhuaitA0URmZdrKnx
noWDiBvOTQLb8Swq+aDukhg7D6eztGW5qeuw01Vp0hW+M8x8inVidaLgRJhsSN8cKkWTee+xqT59
4W9FxayHXUov+/J7zw+cMbPbG9ZyotWIli3fVl5idp7009jtNqAwNQuSrt9Yl7sWNN8DtNugTJWR
RygBy1qNwVOP3YVt7ddWa4XR+OMr+AhUg1a2EkcbHuYLKdxh9YTEgPZI8Bqb8RiJGeV96viNUZZW
h/+/99t/Kgq7mLtbjeP/n0BjoP7hz55bpZpQi9eO3UvKq8v1l+rC56NVusOVmXs0qlSQE6hg0qJd
L9XylYGpZArTlN6I0+uEc30GatB/PViH160NGtYTqUKzN/FIfZRdJYfC0+pbCORksIYIssKZKHr0
tx4SY5T+smmzTSHGrTvKS4HLr/08vonULhW6a3zaNrZdWWB2Cm+UjO3w/lot19NgsdsV7nq55B5J
qxzT8HBaXv7uJp7BX1GJ26YzpFsJCb+eVBnv2ofnukPJ7A4o0Fu7SjaOfpOBAX1eF0vRxXGKJhOi
OWzDl3+uKrLfXcT9InTiKCzzUXHy2B/kFYT7ZaApqIpJfWYB+z9TRpX/YCGtrU0NpUCSC9L3y94h
OZXW00HGgeU7u1muUPGKq3p4lQMDdT1ib9hyVLY6x2xCXeopER3HHqJ2xlAiFZHEvgH5YcCYDt9N
hmVn7mBIxBXFrWElmiIZCugXXUN8y/s+YNg8wmkPp1AgypuCSwbOqJHMdqI9Z+8a5rcbopjRUeHN
8oryndPU8iFJWHH7EfDGMAvYnCu/HwPPG+8qPL/aALWcrVCCgSmSTPRUuJKASqV+VwGxTRukD7MP
4au8EsS/ZCiOMN0Sm4KuZ9oYp9q1HMo5cJqfo/eYwrb5+11RmHFpnl09W8k3U08psxFqP68tRSse
xnjLQTY1iXhcdPCWRuKXZzsZsGOE3ovZrzHH4WzTfGFH+vaQjl7BoGtT6pWOtd3zo1zx01MMbsEE
of27BIiOd6Fo8klxuF3CESCx0GvLswmgjd1lwg+XP7ny7N861TIplwPt7EGvlHyvNA1kZxPGHrSi
LMDOw9uRo1vOKeLDiMP+ExTuc+/Y5ljlD0i4TqTTNJVQGm74kTvgQ72lX1UAEnecC+2tQK79bKsc
IfZ7n3GwC68ADoJB3dw3+2pbk4LDsA9FWqffuM94jKAgKIuzS3RClo5VHiNnAufTbHGCBcVnBHfk
TOvebID7bKZPYL5HUSlhpn3U2jmwa1dRbZCg5d7V3x0QX6OJ2NdDo1jZRZphxbf3Gb6q+fsXrg/M
w8Q7pIfda/bJZRZaslT5TJ2usi8jR6w/LlGNpsC9X1HcFyBysfNDAHJZO71Wd5h07bNiliimBWa+
RW+Ud1uNS4bGzc7jkyndYRB402NjsCnif5cPQ3a75TWXKYJUEozi8Y9pSJAFSUEPcqcNMFqEO1QH
Fwe1jFk24tbO/R127p+0DRtLboicQpQzEdMi7+RJzxCYJYGFSeWVVY41i9sSdqaKvtQlXMW5DrXg
BrDmR0glPtV0y0FZ8t6AJwquYImmMAspF7Zi+oeQLVH33UD/Wc+uYf5y+0LsOmMFDPmotzhYA1Ng
Ns/iyrIHrnA7jiMLaL6T+RBg9soc+yr5twI6Hq1NAb+i1el6SgJdzFdH2n0n2vmyN3Z2I1jWd9Em
BN0MXYNbjdcYQhihurqZmxRlDiHDlSpNAOrM77lnsfcte651dHFNej5hLmWvyssE5hjpnlBbQDUz
EVDCS3VeklN9KPgusQXH40qvFKpU/LmBMuxNjt+m6sBFWU87IIdtXtmC6LiAfj68bxbNEblQULQ/
P6wQwxxwa4SFIS4O8mx9w9keIJG5x2mr3gTqurSHJn/baJVRBMHvBCkt6NFA7ukMrKz6LQ5j64za
47PccEZKkXVcUYL8fx68A63LX32o64Ma/6S+9fAlOe0RDbA4WU2/Z/C5Rg6IUK9d3poazFnzetBY
KA1reulwMDMMsW+42qI2JATEK1SWVabba6mJ7UmI/2gR5dGX/Fj4qahlj7DONSaKHbrASEJIiMio
y6HCbKfOR+UYyFjKsBhqzsVb2mEbvhog+k8weoZBv/e9BM6vgcSaa0kEt1Z980hUtrbtsuiuxW+m
8H3Apo+I2ZoiMBVS+SY3NDS1hjeVxB73KDJO83qmFmwvLt7+BAFRKe3ZorFztoBT8CkxoPV69xIT
0UXAd2QNDLF8AIBW4L5xCtxln3m5o4RcWBPIDNofTLJYD++tkrq5PUJ+nWfe/ZBdohWlWyQ9amvs
LRVC3tv2dftoNiiB+XFhqmiHoPNyjhIIv2dR8YIAjZs4vFaSxQJ/MDTda9Am1iPivu1HGFfXd+vm
hgJuXVd+XngVxyY908C56i9OA7i86JT0on+5Ln3Y+KGuBWEjFFM/f5MnSW7bpSMo7kpikgIvDiHe
+eUObbLu2tGJQdbAd9Pi+l0ynX7j2g/RFNMEoqdan/DSBrLpzkUuIN0fL/FdmVrP3f/MJ9f9/xcW
No7q2narQ7SYjpXED45kRpA7E9QzqL89vwKJZ3HaGyMgJyFDpZQiPxst9LcyNiBBJkaP0PqH30MK
Mrhz44nUZ9dBIHlkQMiMjgzEcT7/wht1beRGZ6lvNtjcowYzqL8W9g31iyBJnvshgrk3zv0cTe0G
aU3LoQffGepbSJ6NakabuW9jeaGZ0bVqFg8PbpZrQ0HAnsWvSugaw1MUyhdbytQvlrem/vBkS2uO
1IlrL7c1qMtiDh0xyvjyccz1C/QvHjKX/6l8KyGPOEyRiEqqdfSECppomn0EdDqe0bSgojaSiLGK
A3GLlmaHE9mhI3hQDdW2OJWu0haN/j9hBHGordgR6oThvBjnqFFeVEYAM4omxN4P8NqLrP5wLRJq
/eMVWrmGwSSQZMfA7KoKJTUIu0FBmQ0a3lJchbqkSaUIAfIIiwT7eIGSZHNvPGskdtSjllANJzI1
02sbwAK/JITy2gZsukxlz/shZAWK3u+6ViaaK9rBgx9WhRrLJaL5YckUsiePsL5Xzp9yvdxp2uUH
hKjf6CF7/NOm/PHbbJXkl06JS8kObj/w3jrJO2fs6N65dCI2mGhK6ManEe+t6KG1yPBbpjm2J6Ru
pQi04uPYgEJmgc3xxF67Ub+Ss56Yfaai3U0n9EzduiZJNtYqsADxjubNstIFY9I4T/Gt87FcjOcu
xGb/gXLJ18MQIa+KvXNx/BHFWGznzxKT91EhW6KkqIh/vy+q2Upn8UsSWwYdo5dy83Jwu3y7hh+H
XhcJ85E9MNx031yxjQEc8oj0PJK2fsE8P/jtJukg106jDUSQBDTXsJJ1N7qv8/PBtyMIA7CpaQt2
BIag4Xzy/L1Rn2DNzR0Phphys2t8vZvxT/+K5Pr/6+zSGi0zNl8DxlD/NMn0PgpeC0FEzBNpDiwx
kCHV+cxtFEhg9XkXhvw3y7yKJtzWjSWGW7d4JI/zDdMCQKpureEuTJ0uRUlleZfoIBuvRxEyv2oG
YXEFjqhceohVLdHdlT3IL3aYKVEpQgiM0u+lNYl4QOU4GyCEowHok2s23ihqUeG7GrXCbBPJCNpB
EbY7GYuRHtNSoTq2EqkGnQAmM90SqQOx3SChhWLVBH9PE7oZh30ivJvSix+jUTkmpVbjkt9xDe17
HLbhjJlYiusExDSdCc19Tcu1AkLBuYeSRbyZdUUdPjEz/9SDzUUi5fVAUi+hvyS5qp5RFpRYAe9C
aRT/hZhoMkrtTmTD2DOVYMQbPjWqLDJ4+hYKlsqQ/nFeJRuJ8tvJZTsIYLVccS8brSg//GsWFYB+
9jZVhxlznXJxlJN1sdTH+PSH6ElY17hH89LZvPJ9PCSizKBv1/zxCBb25IyXvPqHJspJva2x1ysK
dRsso+JA1C9FxVf22vZ0T1YViK6jktbo1mw1n33o9fl2dFVZE/EzdHTd9Vm6AIrYriU2WvjfRAJ5
GOxUITpI0MmJ1wPayyskQy93wy93OzbUYxfwpGlTZpa+24wbJn9urK//oEZiwV5zoES5NTrrujGS
jwLt5lTjlZcHNQlg77vFWhHijJEhBAxvN+2CfUWUJSaUMdXN5uqVREWpcV7kKTSTW5w8hiLU9ZCH
msx6uA0g5Z+aPsArsLzSZlNBV7HBh4MvBYXqT//QLGnDFpZlFzx8/WQDtO975Upl4QtBQ8JDtNXb
phAUQYyErRtqcp6s547Xb76n5py45pXC/QMH4eKeffCRliA8OxuGxWgTKbF2UUMz2IZs6RJnnyXc
qsFnAlZaMyI/vD5NPtv/CqUdBB3XQ9cLPahmj6/9S/Mhv7rbzNLntsG2tdavNHxd0I0lYa9wm6iY
gaTnnH5QUGo9K9ZhhWJJ41LRQuTzvJ2DI+PqxdonYSFlL1jfBlZNJazlLegsi/N9DJbPrprBg01Z
lYIp1VaBbI7PErm5qKrzHq6lL7d9tPmOX3R7pBeyZDOmxdAlFZ6LD47cIiLzhMwRGGoourOZNAsZ
1cJjyFaxBmlHHIjChsYrrdsJR1oS5qKgaSivrXTcxoolMT1KeEuw1Cdh9oI5T8wVvfaHGL6GleRl
zlW82y6U4W9PkUZyDLwc2fnbSkKebEsdWQeQTrE7xVmyCMsda+Hy6wwoVANRGODEN3CF9+D9D6IB
3uItpKOHj+wHXzz9nsWV4NflTdIlhkDAnjskTNk8GoPZqcNtsE3hHiZtSOqHuMFU8+8PfV5zLV6y
xI5sLdCNEzBkSGGJmW/OWpcEfoqzZfvfOmK/QjshvjLqWw9AkX5IQiP1I3NcvTr6HaeanIUeyH0R
k7plxXNgcvgHHrwOnKT+79R0itLngmjxr+iSww2ME2RgxdWnb5bli9cFQghDPwtH4acrCpAOwUAe
wX4rk3r75MrLOmZvJUW7wUQqNu607wcfRy5HGVoDCm/Q1hU2OqloWQ/MAdHK5ABAsTO5ZS2casPB
1kmU0oW+cSWnMXypcgE3Isi9J8l1BAx8J9FabuGiB1djpXmzYVD/qLe2w839ZqERxxWGUcWCd7hV
tJ9aWk9k4Lo6dh1FHtLzu7nBAkahskdwbW8WWinHBHw+U2T3q/K3Zs1uo10EtIoPrZt8wjOYtfon
Muo3oEWEOhGbx11NzsosHWnFCSW8lyF1KRWAvjLJIz+BMr54RPQJLUS5OpQWgcfYC8tMBaFVSHV9
hsotyTqjZDn7b5vvphNLxkGsGVt8v2wTQh0okWoGvtJUvgsAb/OjtwH5fnNVTHsu/th6fqroFiFh
SmmE+MQylwlWZlOyrHqkWILkJltafIoX0fY1WrmgYEjvcfj/MlL7hHI/IkxR5AuuchkicifhJwE9
DJM5Q+ZxaW2biY7UzH12o4VXkUCX6suUXeC+vcwQV36JwF7gYpjxV7GBHwGHF5qyyak9dVxlAhxD
su7kJj/y1QmluF4U9hA6cZljQ7ML6pkvJV5dXCmWM5YTGU69gge5ntbSkL+9sMOuCpC0tva/UYQI
B8PAA/Ci6vwASTFdwZHBPM+R+jAsa95SsOTqzRE04neHwiOrFhuAE1ZGKUeORhSCoeFNCYY2KUNO
zojuQLpD00QpCxXOdg3/RDiXFGMkqALAWOuKD6X0a0SjqWDRt/pm3iFN7Fh3/21bQu9WvZuI/17O
usRdwBOtdipOS1XnFpSsCbAg2DRhj3/cu+omGGXUcBHnQu4XigjzAPuKYLNtReRnAioo2hDf0c7S
mW2+H1UbR0dL9Uh+qZiOtLop9RFLDf6nXU2Kj6cUqoBCecS2MvhmUJXP+ym1kcZ6Bew2Z86k4z4l
3KgreBHWxq1dJe1pXLYxTHOGQGsDNERNRiiH3U/qfpwVrjrezMsK9FONwFsSIIGpGlbmSj8RIryh
u32ps4pi5gK8at3l/+49va2qcSpGXCbKdEPfVvxw/EycQFtlSL9yIcMXbkCwNRVlUcHWhsU0yGId
hBORK0PoccDIjJVcQAaXl5igY8InTV7NYet9OWjA3WFK9yUKN8yJ1UxYW69sZ6Shohftqj0lFA8N
J+sUY0qTIdMvgskXtdsnBduVOQBVBv0qpG4dbcJUZr+Dpmh/YdkAA5bbAWVbhVxMj1acOHtdZOfT
qabu70EOUT7YFq4jicy0iMZYKFJszwi2Txrkr70d+sj/Z+fSu5gsaJAom/S4lk9MNP3s/Gk4GTt1
HcBzmZNATDZ+WJD7jx3WHCJV+G53DNSCiqYgYogDm1S65WysY5vw1fwm558foewWLp+3FlGNpJ02
UbeJWFNNuRv9w+WYmg9b4HeK3JXNCSetTK7Ocl7sI5E9hWR4h5GVScQ5OScaehSxlINeyh1I5VZA
Mvu5GsJgxxL1tm5aa6kGmL2PY3M6NZrCyOP5CxSu4cr9ixQiRI5H5jZkqD3nLdpFot4GC/96M2Am
BNFNPkV+YcttFUsoeuNEAyELcu359TR2EEpcmYaiejG5mGUrsBZB9Ryx2SuhrS6wE/Vrf7U8LMmD
6TTOqW2Jwjoyz+wipC+GzskJtrjdBqiougCt6ue0UWRi3DsuO/ybm8D8IAeza3B/yuqqpF2kmzUX
FKjatXho3lwGuh28fhy23v1YZQbUtaPSq3MLKSWgLrGcPOzSJ+WbzOklb4Lpv5TkjG68AahliqoY
tVc/mgkUG4CA/VbhQJon2tg7laq+WseJK6qw4GANcNVRO2uJFM0sEFrEeV9NGzveat7JE7hFUVwg
I9/WywXcVbJYFbbtr2/G6nQo5KAmVt7XegvoUqkLFWBmCVTeajP6MgdOWkpK1TZOF1j+yaqU7gvd
XsN8kJ6nZsoru7AOhShGKtCReZVR1agS0Hiw3jEEFvLzcx2o7ndMRJJNtEY2a1xV3L9EOWCjnj5p
j795SQutMXzkLy7RXYDvtJfo3pXmy1Heq9Z93VTEfcq8PIMZkm5FKqe4vVZhk5l1RCgZJLXgMFhr
pTID/+H2t9T/xGbyHG3SnvFMzzf7fdxlGQbLa1iKugXRavyIO0PEE9sMtV91FGFA66MYBzsbpzXX
IWUWmKm5oUTJVttaa3xLsKzV10tY8BViHrsG93RojLPSFNSIk7Z0kCXz8n7bM2Exs2Y3s1qVNWd3
vv20wfm94T8GpQBnalQRjsfHl/qDfzOPgeyxROp5yoZncrqRxlwRFwQ000l6U7A8P8ToNxXgIowK
A/UFgymhY3SYBJrX+RulRnmKVF57gjnqGQTHFkjxH//fPTiu0WSYq04yFVBfzfcFjFrr2rRjlC0D
KJVqdXl3MJCkgFBLqFrRx54hNkl20VzMtxJVYMnOxFl/W2ndNwjhr6euQwJFda17CxCIEd10G8HU
l6OL/wMBTKh6YZ6x7UHwIgQBg0bm/BBZ9bU9B0wxkT7z+K1iprfINY4qZlETZDkCOqOZYBh035qk
+NeGCwGps/F4p+X9bPpLvaJ7XZ64kc6eLaxBqFNkBPtRf4rkG5+R0VuZbJ9LV3XigHOxumTmrjne
ef0EyfOjzPET1/nM5Hab8JfWf5MldRqW+l5xgvjU0qdgo2FXyiHTt9zQhAdNv6FTuOI9mUXvHZ+x
Qz93z1zVpG8E/Lac3s7JPomwjedBjudCKeFww+UHVid//DFQ6bttZXfkjhHBdPIuGNqgLiYtUwfj
yIH9T8zc4GEA/H0N1VE1xFiQ2ttZvP1QfkHk2V3Zg9hODn5ehob5LC0thWlUNzix2/6WiozB1zAy
TRKRLp4EvDa2e6R+vjEawygRc5yLiNpqkl6FCqEMO78ZhJgIx9J3oGodFiM5PY03aMBLyy9URv/0
gfI7UkHhEFUx4d93ObmkvK/X5mKeeiIsJUtsailOM4DEw1WXqhqRDBU56M/XNNkEeiemOOIw4gKj
orWaEaebWDAy82A1idaVv7Y3W4ZsLg2QPw5PyvH2ZmoAa5ODlPXDH3pNo86e7hFRrMgIodT1aUya
c9d4cp2+vx21Y6I93cxUuSSxsNK6QzW3Cvx6jkiBXLiFnRXAwdJvNa84nGz/BHXBVv1PWdrZMSfT
g+KkvdG8GjO6/c0hfsFlU/Ufz7P/V4rq+s05V82spzxu0RSYn3tXzkoZLG5a2dJ6WFlh7tsCBVuC
gzA9V9Z6+SoMnJJrT3zaeEmOEIjhq1UsrfxuYmHqIHjb0uLHXSPPszKT9h2YQ9cUZlAaWT5h3PQ7
D1gb59nww+I0yYTGHYTIh8UcJ+05ERsfKOeV9sp8RLuuqCSqqOixGA4XxQ23CSHsnGg5TAz45Hi1
plg0usCPguLW9YtDViErNOYewkDjXuFCCaXVZGKvgLzS+1+VK0rn/+/QbuEnQ1skaBaAgcoq0+dc
2IjGRiHc6WNnu180wasPhR1bZ9mi6aWbMZyYUFJhKVaae8Ihi57IfevQLiCfuaDRjuunQFWlo1Y3
7Ib6JybV4WZizNEZbiJGm0o/ouJTMsVMVSVzNU839s5w3yVulGqS2jyh8j6pOlhP0kJdc3QJ4/uk
35KC4m/5ADK5HW6TuIXmrvcwCYkumoF6S7E9tTgM9EqDzZfOUA3fRqqLtfj5c+xn/+vJ/wGfCVZu
CLvZZC+9mweRZ0PM/kV/6xspqV0uOd+WRUYRM/+ZwfD5oBNuQYI2u9GNBUyJqod5cyGCdzaYFpi/
gRqMRLssPecW5QUF5CoGAzjLWEQyM/WAI3isMU3dVje1fe532EH6xqCf/41SevpgP7bxCyLipN6J
hDJ1A7MfFMSNy0fCkLZTEolewbGEVCaHExPTYlOuMNstEkVH9WCO+SLAzMx4vw99QG5jjbMDkTbl
k1TrB1Y8xbqdw+B+g0ChkVjvAW4JtZr0HbOcKBKftQ3oCkeENpO2Ti2eGYMFo1L66PhzHG3NYuFy
HUNCyC2biQWIjgYJ1YgG8F2z+jJcTzfgoitMLTrX/El+023KizrNDC+CzPL2Q+9/JaFpQ5MT9abT
REr7AmYudHOja6kExk37XdJO+UbVPHwIJKHI6bvs44GEr1P2shYSomuiVU0s3bXtgqSSIZJLgkG/
O74wCjwZtHK/Ci5fyM0Y4HxLl26lHxzl056IHW3ZhVF8LsPYS8WS3mAQRiIFcPPS9JDyAJVcyYg/
g76W2ggtZf0x5JM4PX2UIj76ZLLkQ2J//eZsZ/oBeZc3gMFF413K5OMOgT2tHfv+egkC3kaNB8re
zx1ms5gsYmTXDFnClpdWpVIHmiGJdVIGBiPBQAa5DnuuM/wv7O0Gk8Qrov+QNDiCScqDQmf2f/z8
GoPxuV0rpd4Cseoppboptzgs6Tt/HgLnjhvBfhBBm/uyTZiLenilYD4nc/Q67FGddX7+7PN+2e/+
x124fnptHp2zW+AfDXab2INjyskUw0doXJJ8Jme+0WVkCT8VuhW/A5ASQOocJRAoRUnX5jM925Fh
39sPykr/2DUujQR3Y+QSzL/1zXNvbXy8AbVHXDaRXNmkdJ0c9WdQqPh2tnjKYNeiknwrdHrdomqh
QT07ayCAMhAvQImloE3eK0oMo2Su/v2Zkvrvru+NA+dx7ebjBPav27lNO0aF0DZEtZG/ov0RrqUV
dNsvdJLFyY+hL/+eBWzV0qpyFM+ItylkqQ+6isLU29rYZL055yND3f65n8WJN7ZZZZ3q2Ha3RZTm
mk99IECIq3OTSupjxTHu1XQZTOOn/od/iNKgrnsrxQG3H6LD2AlISnVXIvH5zrKFYPnytD5VTptj
5VOqcmaE1CSHsk6+ntSyMN3JLCOB/csGXWrw/BjczXAuKsHVRfZLFe00Kta5LAJZL+/5sievVzA2
Jmdb/en6JnSjhRAugBHowmFIooDECiSvejXeReKFCLu99nvMXqVDJ/jlJOnUUWfFLSKS2ELTMKUw
77Rmh6EmD0kZmzmgbynAqkhXdqj4qNRKNMdNN9ZHXYjDZ22dMcj1kSJzc899Bux7+JsX6WLcCP20
KyPndyTqGeXwdif1LzN9iAKTBUY3+YexSf640PilZgtqDiqiyjPxmksCvV/Q7GJpGXH+rZw0nKMl
IYPX0kIBmu/EdZ45vL9/NIhUQlczBoqZix3QF7xno+0ofbqIqZA+A5nGvAdISiOBncQnh/umEED/
ShobEATo/eENfirUFtirvUTbKhv9pr1fY5QisqPwIu1NUA3b3aWUFDhgmuP4L+laCWprijqM749E
9TubbyL85Ke0vUAhoQ16RLwoZrd3t97olsUVqiqexBZuEnHOzpFHNvUMhFGZjINPevNjY0mkTfX+
OW9oAQ6fwCPKd9LZRwuqTUF/aYL162yTy+JKS8OOeyHfpc02kyhbU5gJE902svFYTMWdHl6UxwVb
hr5/6yPC1horFF4831SS+UX9igR75y+O8mRMBNdPczRjzoQwmk85kBTFZx/fvhUxsDvPbePQNy8e
glST7FXFwal0+IccDM0gkmOEsEjZTF27bV9U9JVrCzjZsDwc5/AdztdpxpOb9cQKTG78mMJ+ndyX
10FbXZPaqfk6bc/mew6NsWrLIGrtVcSUtJdIcH9zrjntFYuP9ER1QPiek76yKKfHS0GFhEKPhcfc
9PsHjh9PGysbHUNnabM2LWbBlcvRXXD3LMIMaqesE1KM5XPJCi2X/3KCWSEBjYwI3csiRD9jQgqh
+m2uGt67u23blLxALh2m1/ksD/W3IRF3bWsZK840r0QAf7sbxlATquQp9/er2S2vMi6844sy8NpE
yhX/6DxxWzZKr6vF4EHoxI1g979wuR3tUn4xEmwGCPH/cOBkoj5W+WzpfJ1MH9btXSWbdqPv4Jrv
HzExWI9o8ad8wG801RP4DLPuPT6LW4t4kEpfus4xwXV/IxOgLw3EGr02q6TRhEZU68ULTl7utaGj
8vCnWuVrJkjuKh6sH3KI91TfOgiLgvWnlDx1IafxWQeOTO9AZZds8z4hewg4z1+v5HKg1t22SXex
EbqHzBXKBbiwSbGNV9ChXG3QWkvyVlz2pnzJ/0YnLCbjXQzYo0MM/I5mB6lEfIhgDmd7DxpcbinA
PD/pc8yv59QRzD29jlug2dvWMvycssyFvPTBwUHz8KVaxVA1gAD3KJXbLm+JI4BduKCkd+h+SSyG
b2rcyyEQyxvBr5OH9eDYVoUOgD7WzHTP17M8J0CBkqw7B3iTvRfQ1B7fTVUCM9OJrPUbaWrUGcVC
K/o94r2CI5XPjYPYr38w8zPCIlvH524zHt3v1Py2Rw2qZ9eXPomQgO4f1cx8r/dOS70k53zP6pna
ycqSrwjvOSqQd7nvoLo98aWsWj8iLQBf76juIqT6Lenfn7GTjqUTPUKFiEhoeb5Z6T9+MEY8JdGW
w99ubDnO/HixsbEidMiUtLSrM1GwNVmQ+CJ9cmeBw/IFRuLgRZ/ccYJlYWeFU1DwTAxiOfDQ9YtF
E+fHYSsDlCah2yaygCuVgk/jLiNypQNydStKt0cJl78LdgCaUzn0aTd6dL5LlGLdW9ZABXXc0tCr
4xRsYuOIcPM5MhsZ94fk+A1M+oaOykeCEd/Q1WROet5K8WSjNF7aG9FBSCHCigyRyn3daRiNEE4R
vOi/UDs7Yk3d6T1PnCAqLJ76cTVft/NlcscCBmkBDAL/fgy7CKkP91WV1Lud3vLIS54k+lloUqJi
wRLOGN3jJW7zTZWsrnRdoys9Okjsrpocto+ErpwjdObyVnY0fYKqL//o8anGkAN01aJuRrQgP5Al
jsaU5aDXFqvyiSeS8qsR3nV+P6lPsBT+jtch6Dj5RbK3ZVHTiDuGeMwz6GFDzzQS3uHRtIVLc4eS
m2FZHFbTUWMt3X5M9aa7TbcI4ZHJf5DNt9XBQEFMC8KO7jU1DL+ttrDCblrUspfyWTecGpnut2ij
Pl0p+hz93QBYxv1QNThY/ECOFy9e2t8e45UeOzh3VFYKbAZKpeIxa8Xl8TPShtia7MlkD5DtYodC
4I4ViUeUHDIAiUPtfnKaAjVp9rgkWRJ7fSHjdyaD2PamFQ2Hy1i3Xk2Ldt9NZLA0rMTpdY1w8mCR
/Go82qMW6dD1JtTCGLwveo9SGE/u5epHsEQRwxRcbPJQ/271mk79ks+qm94ZxYPLHOr8LbZ8xyAF
WmBPhZM3ESfWwthzVPb/oxZqtUn83Rhr7bm1VhcOHKX4OJdOdvJwaJTIRDuAV6FhAl6zYIoyJxNu
wcYM32/F2ryY29WhaA1ToSzcHjZt6xrOd/+Foxw+2Gah+bZr7oafqAFZSvNAfyFx8YqbGXup2f59
830Ipd6fvrsJMF/V3XyZMjRRvyuPSnG71OQzewNh5Ps2Tshl8gJvCVmhs1jl/2bsZtV7SVI5Hevb
vrKnWN/JrzHWY0qS4nc+MOqF73KXYeV0eSSs1Sia6kq5awf63Xv8DwFWazM+ndePfOJVZsPYakNm
3HgwrTfpAgzt7amUhNPsQNQ6aWCltUkfKWjjOLMQz6H65SdPKUOqFXYyUvj2JjUYazCGSJB4FoVN
MV1kWcABvIVFncV+hIVkAyEP/6Q38nKQbxBuk0euZxTQ4t5RKNc8cULgdn3tmslvoFjjKeFstYx0
npgBo0PwLJ8HqAwkyT7YXAUc+sVfq+CtBIaEYB07AWNP4n86Rex9fh25RcM2MbR2HtsmLnpxNFCq
cumogPXYrSzfjcOcpBLb+2aZme0/Tp16BHmmJNyPBvBI7+SeXBU4b6BMHh2K4P+EiAcnxncJvOUk
ZbKS1XPYZmlejf9N+Sinhrpnz7Q77rXP69d4nvzrwu9/RKETQ1EskoN87E2h+CU+R+rhJVQaCDfI
4mH21NDK+2wxTBVloZjwzS1tkPpvdj1Y8bZQVa0Z9VaS538ZS2FeToPnxuCjwrnu4euogOVzyA+d
ykAJP4bX5Lbp8LcCHPOWkSiJy3BapHsqwxBHeHHrbspZX3+gs3bSnmKsRNLJJlAyBlhqCyE1NO9o
5SuDvigDBsvHQXwInPZBaXsTjCYZaWEuCEvn1nQORv9K121kPP+oFfc2WPZ9TKQJbtfS5CfODNeD
WKrKUKY2+2AaX7iRk8ZD8bry2KQNPGsoO4SN37AD/FWWboXzw4W1Ihz+rfcQL8tO6rwubmgEBGjJ
CRkItUe/7mZJXJ2Gu/NXkcft2SBJRsoVlc1pw7rScHNczQAEtbMESSjorZv9Aq7TwNk6B/VbEExH
Mm4kZLhgYqoD2P6LKdRELKdeeXVdSjW/Oqi9wu86f7qsg4sgIVjsNdkeiGb/lUUNIXag1q+ckwQV
EHku2X96xP8cgW/4niSFnHhjCAvc1F5Djs5NwbGp4Q+KT62xPGIG8Zu6l+I8phHpOwgrBnSSISiI
/GRF5W36XzW1hqnVYQa4nGHiECwE+rn60HJovOeMukgT9PJ6n+koRkVfTow+vocRuzUk1QO1KLzr
FQejV6pyU8C6E8ECu3FmVazcmq4+Yly5eARRWbsLnYCOcV3uaDaRjDRsbLvUYpWVu5GQgDyKnGXS
RZMbeUVT2+5FS+TqIMInEwT9i0Vba71Nsit13slciflHKYD1Ac45di4FEmPaw/aZwBHMpuop7sSz
t3cJ4VYRxgHMunc5Dfxj+uXrqzSiFW9QDGXkWrFuvCMZ1ytFDDiv4igEgPZp/F0gm0O489eHOFjP
P0cLMQpp43p2JUHN7g+wxJsTbsr5FlsnlblryhGa7xKfrYWARJw3tLn7mXHFedFl6FwJNs1pBlHD
53RkMM1XmbS7cKILI/W5cNaBoVtFKYL/evF9sFtmUR93HP14N8CIuAHKIZRq17cE7hnT+mKBoMGm
NuJOpkB6DTwQsgUhwiVSv6zhjtBh8UrJiQlH7c7FJalCDm+wDK3R9GYRgxWGZvImAfqbbjp4VhAD
9ZrP3jYccFlqklJP3QHWVOqCQZTrs6hYgc+eJgAsw81gNf5i52cjlEV9FVczZic2J7zEBrjkNiex
/NVcIbSquesEQfWY2HT3DdcCivYVnfldB1URnT1q4Agf9dQK+ZBZWWwqdZ9KnTHG6V8xnb8h2gBq
KX2kB++aWDeDK97Kv3HVrnKLfPqc7H5nkUQaVwKi7ptGvI9CERyiUwEpKAA7v3QWzqyFQgLS1gty
6/hpgo0rZeXO7lsCCy2vBArNG24d2o2DVjLon2PO4IhAYmxk+4M1c3gsb0W9j1unXiGztk73In3K
3pui7ltBc7r6L5FGQuR9efEUst+mm4svTVyI/dWJYzzQTKrswoSWHl9BVgEOnKCPDqsCE68tIO1/
rTBpQ5xbg/xt5qa/8sSauxkSCB/bD5rQLbqZGcwJrIrBZa7qhGLVE/iSWM71guhXlW03sPs4A/PA
XnJzzxLDyG/qB2jqL7i6VSxTN0OkS5n/8RoTwMaTlt6etMksrx3UfqA9VCZxcBksmhweEOjap34L
sIGWFMXpqXlMdxkxx9RNaWNNDH/dVTyW9DZSa+y4W1kStISDx+cRy190HmpUFOlRMQQ24kf7sqCs
9x5IM353jVwCNmnA3pJ4NBh+UIT4/XJLgriO8Xnjw54/D7uzGFGBfVyW1orRj6fvenn3MQeAJylo
SDa3YEf5GPaq9pSVAmaj2XBGHbuCKCGbejI2JeWMSgdOUcxQZrUQxlp+IOAy8IVbvptsOaJBVo3L
oi1fYh38nn1Zht2cYbugNlymvfHtDbUB8do2NTawpGMFswSHV29GJDGLD2xvv+WngoSYetsvpiAR
1s2wcOyu8EcwF3Iv9MprH9EIDpVZHrgCpupZdN+5P6AcGh6Q1QcLL4DK9xFR3iBY3nUmJv3CVgBl
wQp53cZlsNgKjNlk1DzNCtcUbLhxLopNQR5WQCwxq+Pc16GnO0oDIk9sCvrg8oJywyS8aIIh9yxQ
jHQ89MT6M++Rt8OhW4LpcDOns4Nn+uU2mDi4Tu5taJQD6wGmv2HxybF0RZsgpryI7+LhIpIfJSoS
aP6UjZ5aVYJn1AZS2YqrOyUOzl0tAtpk4sAdxqRaCTiafjkpNkGFw1lafm/S1Z5cqe7OOiakpQ7n
SFZgtigWWLTMN7DKqL9H0YI15lYvgThoU21Bm24LFq3OSx3lCrlDlfWSb3lseufN5RpvvTBJc5on
KRx/SonIJJfQPZrggr5Rkg1UgLAoeaA29LSY37DA97rbH8Q+Y25XW+qTXGDLiyJItnBepj4N+nXd
sfBZnajJUv3XJsWDIXOr4an9K+fGkVig7oyBZPWEetWd5njluOHeeh4Tli3tR5US/mC+RshtkInW
GJlYqRJmFwNjPRfbMpoRB+K8HQn6mPE7fDY+L0hMCCU2zYKezz8adr/6o2IjL616tLvz9qltCHYN
n3WxCacteGNUOlGN/eujipCzrk/hOmKEmKRd/1ONXtOA6hP1BwBXHaPmdcY4mPbTsS+Wgn+zYV68
SkgShobjecEkKCtb9Ea8g95hcEE8vksF1OP+AyHhtkoSAL7j1oc3FnxqtbFIlxNSMlL7YeCs+gQK
vtlRaWeceGOZKFWyPaEl706CnyOlzr3LNQQyVmlT4gGRXv8fe3LEO4ypROsZmPduzgLv5hvNww5G
E9vi55r+EmchIOXQpDP4DhUC1EPkXDKGzuiuo7hUINeEU0Uiz9UFxkNN5sctBKPDvwI2mPZiY5j1
rF9E1w0qlpCJ/lg73rOsC27nf4zwEcNVaFOiG67T59BtEmwOTypaqnjWe09KBWkDP675SJWUdwU1
WrUfymEZaBL9qF5Ih8ofg0QT9eNClSBlbtYDMqrboVOjrpUKjmOkufCn01iSdN8Th8vv+7oOcuiF
WTOQNUXdtXMycOFtsoiZlyGx2lSnkDbO1CiXyjzHsEUS/4ErlRiC8b5r4tdzBP+Q3WFXYI2OsCKV
LgtcRsTMMsyFt8YhX1F01NO5u2ajXil46fT6+R3AxZdRd0VaslNysHa3f6ueQysul2Pj9kUECATD
3oXS8kumMeJoEtjMLRHb6ScH+ldwfH5EzMERWXLL5T+8ZHfV2FoMs0656wlAvwlKEgX70GX6FF8w
atT4Zd/wXV72oAq1CRxLgPZAhhmjWK2INFh4xBUoLBsuf0zVa07asyaBZmrRgUXCQj3ChlgOIxvD
psLgFAg/8QisnujPolqo4DDdtmkQLdGAEez0yLm2sNnoPbB2Yvw8rFV3l/BtqVgcVxMnFopDaXtR
oFdn2FJfVZq6JV6xzFtiMXUrvANAE2BIvEvLafM7GoYtHAZhCn98wFq9L/91ry+dS91D3av/46BJ
kI6UdIZ/0rM3v18OYyzFQWJ+nxrWOxe5ByDyKG4zB8RNWG3Of37feDf1Wl1ykRpadqfVJMT3Kqbr
4Ww4U4Ytd1cs3BtUxqMHakuRIAglDl8iH+NMEztzD+4abJgNqR9fkwpZ5MN+WzJYrENSiRrArIdj
ztZJ7MSnla2gGd4JPjlNtcvHEsCJCCD7uvuxcWKBarKlrbDbPizpXOOrvjQCxjWk8WUphNOLqJVa
8AtNOi6+927B8Vrwv7SsA0gu7GGMLqo5HcEmqYlbYdFdd+wLleCAARWCQK4RL32cj5ESmVFsdGqr
85si5fgSkUKFJkphxYFoJSS+EGAOrl7hcaMUwInGtrq3GbvKKcXicjyoV+yYArwjrdIIYunV1BsG
b3OxWTRYcniY/q6ZxMKWpzSsaGm9e0TzXM0clXjuMWLZOA6s4e/ZUg4LWBOGeqSc4vtcQNDawkkW
NaEYrLQ0WujqXKyeUJvP6cjRFuI4HCUdfxsdbTcKrFgk9+zl9EORjQmyXfcd2RoC1JFoeLTXWhSu
sImSZBMCid+qhs56q0vXNmvmkJPrRbmGIMHjFxViuGrF454b+e2izi43b7XoWwnxkmvqyUbxnerJ
tSKgLulMIU4Fpxw/IGZeWgvVaFcaSqr38hxN2hTW/Qt7nt8R3tyr+hDDBBVA94h8IRN26jXGBF4r
dvZu5U1eJJ+nmwjdOB9kJehB55kJ/NoDYpDhsnPVSc+90d0h6YGLz/uYydNdsTdL4OZSTTF6g2QM
EPKQ2GtCcZhXhbwUeMhRJngLQ4FhhNghIQZsEg+8t5ByMxO2xYlNm0TYZ0WrtY8JDWX8nLW6wTSL
Rz1ugL9a7bwu1LTpc3i8uvNpG4PlFci+EEQ9tGLNmQzAtYyEZQOp8fHrKI1QdCwVb3vV0ak4pPRl
iQOIttTx5r2gsXoo8Fk+aR8Ytb8wJnhWuIKPc99KjsBYqk8XKoy7qpDaH0caVLxGnPzt2umbKmOh
yPQIwyhZcMcJmV0gg5GduGoQ9v1opU5tE29STw7IHoQS4ZimWFPwKEYS6sKAf1zAluJXeSpX5j2T
WvGaB8XE5nIM95lnOBxEp+dWvbN/Pj119fJAFqolKzFYOYTvkt0w9G159X81ZHu0JL1Ju8j5qgl9
p/aHkwOfzSGbe1wHuxACLUMjOkEpsfnDe6kmBp9t1TSv1lwUNjZVPQiK4PUqOuuFHRKaCGDL0jSD
b9W/Pj+3VZt2+OX4fOqLS+awEGllcV8R7PjQC0I9T86EH1KkaduWnDimydXCVojID1yAGFHNRsM/
z9cmeE9n0vwCyoM8cAB4dQQGAMpN4R+zn1TTB9NX7dZQUlOKMmOtu4bFibd3B/gQdD9ehPMyYJph
U+H9vbV31iUu1zD3a0PTjXbUz6YnqQ4IL7wdIUlpI2NssoJy/hseUfY26JiR+6snFIQ58i2yOSHF
1AG3hOH3b5IdXHC2t5h/lS/BH2yjGkze/jKO058iBPdv+hUejwQp12eH3plUM1bbQlmsbTdwZfra
YWizWzfP4x3b8x3iM440VxkjqUP5iOgTXpuoKZ9m8yYcn9SaNB9eGlMW/Lgf6p1YSUbk6BYHpf/t
UplH/1jqDbt4cvbO/VyZFazYMb/vQK6CIwTSWiQ3jgRCHMfXoMDFefL4BsBZ6XutGWbwEHsTFB5z
xLDFeF6AgzZciwSvDIpiSF9VKThWJyQBEgKGsPkhzUq1oA66WGvELXusaPJfVzSknNaw1uvyQGv2
JPvjcdKxGbDbWoRgdu8BI6n5nYmQwlojKgymbsQ3B7US9UBaWQXVzOaZyOP+ejoT4/QHKXZR/Ycu
YLt3lz2oEXykmkNxJ0jkLvWJS8mLn3yvIw2xkhDZ/Kr3zCLoPaL0qABCDpz/GuVMuoNgdQ4FnSVR
47RQ3bOb/FmIkRwNrw//o9kVcOaiWFrvUzsw3Zm54Hm1akjezd5VRrnl/nGekSjyMP08kuJCoXnQ
/5QPzJyfOBwi9p8uUQ0eYJIDmb8DfsqLWVX1y/m+mJhoj7bJX/PUb7U9Um7AQYiog4NKt0Os++Pa
LA2Es+dC6vai77KyudR2gaQ2dbJTIHVaH0nrkSYYHRSU1qXl6apF2zGbBZN0/QHBILMe1WzRpmtx
jVlogccknO3gzdhGG6V0p/QcukrBK2jQL99fjjT8bMfyW8a6PoZwzLf2/arZyMysQGdp6PEKnpp4
op4CnTpu3xryz7Zj9Fan//IzdyU5nUwQyIMG+SDXAdzP4jkFruc1RZxMoBHZH/Mao460WC5/V68b
Ss2sJdpla5ZvkWsXH5wor+mlVPU722TfVpCD6hqr3SLNOcuXmgHQJynFmvm/O4rJK+R7ac93nbLg
UjOTWNUPYQ2F4rETXyl8SqQZNRdU43NFsm9RLPVdQ6olGUjG/7EulRt6xoEouTbx2wZYYd9YavRc
Ti2xDkkvIywv38oVSNdRJuKtAR/lUjnlgKhTfQnWz7BpVcAtZ46OQGZh1Gc/WS7vZRa0cOC/XV4T
/hEWJWh58Dnb0PXhHB2fkClyMhYxaFJJ+8UCUBDiLpoEudFNaDUBQox2UMvPIrL9P4SBVi+5paf7
LZ6IQY+Oycj7LO7w6GwQvXGSI7fopAV8E0A7zcJ7TQwjDv03r1iqbgqSOTqTEU3jP29l5Ao4y5ni
E0YvtebLbVHxI2Y8+0Tf6xGaSsqtFIm3nev+nMcKVll3q3rfhhIlf8paJ9IZWt0Uk8VOniMDfufV
1/PHTpHayMpXuqVe4wmYMkKlyT9P/zvqkxGsqsXeWx6t+qqSbyPC0u9xDR8Vafo76vUhXfMcJzW+
p7sXIqyr1XhBHfxA2fE7BmXllFzgqsJM6qnRRVMvfntq8E/XC/0kZAjszQNVFm7ZIQ2CzOeiszTN
ExZlKQAEuEZD/VZcWb6lojb/BYmolBDfD7Y/Z7KZx8kz2QR51FNlKhjBfjZQ2Ll5MnNbBou2yYRQ
x2C38XmIxqNDuA1fTpq6n81jzkY+8pXFCzygBO+7k86WWDvun+oPhVLTZPfmNA0bg9ONuX2fFJDW
R49NRqeY8wjDsoV5JzfN4+PIRLK3xMuzFT//lie7tJS/5sWV6yAal3siS49MjBbVvaiKQ6V9NSTw
mJhINYGLsOBgx8ELkh1BormplnkfSBSX75XLZkDdBJ+LWlQ/LpyhjpIusuzcA2OqtjSRijZBXmG0
3BI9/gmDGUlmqQ4lCGGBXqjVyVWH6gProoZAwLliy3gCSspl8cq40AD7uGPFuKJQRZFYUbIZNOn5
OjmjlzGLsbI++UoJrIkIdMj2yHd5VbWMKFwU5yqQmMgcMrljD0JMXmaFufkCkxlDfgHcADvSJcBn
el5r5RC2gDK45b97IVSsPgrF0F3qVtjz/vpGS/1mgZb7ynLTgp5wmCVdAR4SZlkiVu+r4hLw98uB
3Nb19wsY1VxXC3OlWwNZRm5Z68LZr8pe2EU4sRXJFdN5UlrcQUJbYBdHaRdd38dc0C1TPHWWVasH
lE4thdKxBYaDGrMztJkj+C9MYDbf5xtRi+YmH6ole22zsPs19dIEh+cfr0JQdkKTw95bjj8DvmWL
zbDXOq8P1LR5Bhe7VCDe0mjDJh91C2L2CXH1vpa5qAtPSa7qfInmymOpmsdFfgQIVA8r+qE6L40G
HFt1viVIIho91KVMqm9GzcIZBsSURp8NP1W3ggHbEX/9N2e1m3CC6Snr4r5ci/ksh/Cvz9EWyDqK
BNRbqYek9r8L9R4X+vNLgpA7iXThd1Ritf6mCt5vQdy+x8ngXzaUDVZLz2ToFLasiM94pDbX6uH7
7wrrVy1zEYftRgL2Ncj2DK6ssqEEWpzaqWbf1HiEdSrKBsn62vxEJlH7dl8Sn/zROZDhhu8aAMyK
QFlh58CnU4uRA5rRIACb6tLUgiL4q1xymjBJ3T6VPgO9tL7ncX6u5+J3dewb/XIzl/HIvmQXF4jo
1fjfp9NCGLtYeCaQMkuxTPOZNP9UX47yZ6tQS8WOF+EUM2vHTOMf5VvgOF53cY4hZWVHlHR95PMk
/mDXtS7ZRDYX/NCynCHBOVo2cKjOtVk1Ni54VCTZXwLBw5XhMB3kVC2Q0L4981Nz1P5w8lRmQLIT
5LHn2WwzvCF4ASRjd/Q0p0n4Ssrh1fXC/uc2LsFRVsQ9KkUrqXy6LUxGpwt7qcfLw+FU3o9xrUuu
kPmXgzBdhihWUE4PZOFjzjoX8/g1SGchUXR/Ljh/f1G20TI3AdeI6QGoCHKwKr78S/lFia4pYBNs
yvKNvPGzUmumOE/UsquiOpxJvjcV/sLc3IBSAe1QiFBRbKR7JlUX8Gp6f4JT/h3waROXPimz9J3/
ydHvvCWQEmxNbaaetCdlvRCR4ThoohJXFJ50WjgSWwylZAEeyyX/9PDbcfrr4XVLPnx4EjhSqE00
nTPp98CDbUVdndaqnZyNlgCym+4JPqiMBdGBwn5F9FKraHVghKhOAQDxVG/+F4qdLDVDSlwNaCoq
Yn1zbsr+XhwbixSSR3z2In4FAoseBNeSbqt/J6LBWsn2fkNkIC/lkPHm7eEVwXoX2T1GIK2vwrfA
Q0iHrAcmgoLnBortm17Big6lWEmjJUKIiDPwLfYxci9JhxkS4GTvTtqwPVDdqmyKthIYScQHrlH7
6XRiItTnaGX642X7Ty3wFTJxnlY5Btw6nv4gg+1ZQzFTY4DNuh58dY0YfXLVtKoHwNSUFS7SXNrg
hGj/g7qdND86H8MZi2NIsKZCuN8byfvcddLWxC1+SzMoTYS6rItiq/RTD15v4joe+yxo3x+aN67y
XBpFWumMIGhxAfev5ZQxO45swrJpte9o89X/zHR8UnqPsJKnVaYicclPt7ePMA50yVJ32NA4oHtP
al4HROVAPItUHfT7ToCnQZjwYx6bxcQDAOaWwj6t7NyhVyFgd4BNNJbwmBxpWFBhHzuZU9SPc/IP
NtYlctCgtFbEmfPbjBpsjybM8TgiWxnP1eaS8C7+bIT7gm3LTo9yWm9yq7ts0JluD/sse0v6n9be
9CfvHLh1zrJ1roW1iczQ55omIjn8bbxmaaGmNMCEKlxbLU1BjmZCTWG5OWZMod4B/9YzB6NJWPbm
iMIdfcuYKAVU34+01xag6V8MqGF2UAsFBzKl4hhwLSGBZchDnDXGeCpWME84GnFry6cEATlhQAdf
Mhm/lIeaXvmN8iJWpbJZVuO9V1kIPY1D/NCxqTRWhe8/+7EIish7mHFu5/TEfnI3BPzrEg0M3y8i
v+qPuA+rNYt7J2OJkTWbxIhgDfo1jdL3YTZYmuvVfO+eVtrlHvEw547N9KyOu/Z/hFq22CHhowri
nynJqOE1c93oBJFqeH+mGKiclqFY9tlXO+gdIpyyTCbgSZ9q4HIU8dVwsybA/UvY51u0bzhL+H8g
tQ8E5+LdnNQpLgXFGpM4imduFGV9Ib2X8uqikklES3fHbUPQS3NmhVO771aNuZ7UcPHkR3O36fkH
lvmSZPhyQTe0+cEpZ7o4LOkwVgxDPASLfu5jWOWQGUXfUCM4TyiPFg1IFJ52mFFsQuJcaqdivjLK
G/AnUWywk4qmN0u1ynitniwRcC6YCJd/fMS6V5oIE/LlXvDCJ8DusF0EEkY56bvcOp6dpKKZsYMo
v76AbgIByr4riGoPb1VwA1Ckqd/x1nQEtSG77NnsgHDzObtivjDodVE4FBfnQZCC8PC6RgrN1Uub
bV4CXN0o/8e0L0u1qq25rCcEUbScAnf79F07wq3sLzhYzyiZIFskPVIh63Dj/2JTieUqNj3TCB4n
IAG/0gyWmNST8qzfXCMMSe3V0C8d+Qhiuf7TjwcOZZmnqMwij6d8qZ1i4IKhYChYins29t7eTW6B
H8WCylnOEfQGkrAi72+D+6yoNVDP0cPSxxUfknz9sh6Lrlyr1l/G6Yu8hhqv0mSeQeTd6yXWa+Jd
GBK1viblrJ33b0SYKhUcdpeaCqwNx98AOcOrtyqnKQoznSaD3IrtECQ8FPqheslg+f3jAf+aIv+A
ue2uHNnHLQtjhP/U44RjTm+yxiZ0GGBwDAEdCRqfzvIbQu+OBD6Fm1uqxBpmgwseeaQdn0S7Ldab
KPUJRrY26qmf9sq4EZ3pjw8p4TMkEtb4JnlYLCi/2VvMYL0ueLc933ajPsCM+Crrp3o1KV8xAtdq
4gVchiFDQM/TappLB+P6cwRboLHb/IAhwvWB1a4hLwBZTrEa2BAVYnaWwwnYWlgiez0/86OOeGBU
j1UG5vegIMNzi2B3yw5N3mnR+tmgZj/F7vkNh39LdvK+wUv97o6zJ/Mck533DViCJ1V65aZVmc9Z
t4BxNMclgWzLRf5Ozzg8hOEV0Z77N/2EWMVJgFWIEU9taEJvD58LEcPj0KapmMvx9i26saRQmHJQ
aRorWADboSODo6xd9JJUWW1kSTfUfUmaknDPON9ekGzKYWQbn4mnltyLDxAZitPAIcopfjvkENsK
oiasD5jS/jY0lft58eOXGZwaHgDRXOA3ivb+GeMH1L7FEhMAxPFCwmk3W8R+E4dLio1ZvkE1shc2
s7Du3+vCCQZG1OQxgkOsoyEGntaC/pVYjncsDw/AwoORSTlmEzs0qcjEPfVhyNnWTR0fCSkgqRDM
dy4OgKxHS/viDYPpTdxmNM3qJ8JsvwvioA/TeATV1h8ZCIROll3AYtM+wjYIVuHZGXxVuKNfAN0O
9OlmRG7kioaCleE94GqUGfBNnU55PqxGFXJdPiiFr/ZsKRiSvqYhX4JtViPi9BCfGzdu/NM5YIxv
Z7D0B3uG9V3rgpFGJX/f8iEaP7ESZwtApbwoNYDV7oaW9oHY/5RjXgOfmOtiRYmDE8YZKRIKkRCH
IZJz+lQnvMFVuodtMhEedWAnnOsYWOGlfo8iDtNIKF/TiM55dQyyD+l1ZUGgNiLMBoQiqaxPY4gV
0bnZgT4ancsnTRh/z+6ERgc2HMmtZtg6cOM9q/3vWh1WE0+2CelQevl/0mRj17L0rLhK0O3ULxLO
reSAS29moRqlLOl6yYUFIbV3NnihpI5Q84rXI3Hdk1OoHHfGbulAgXhwR7p0hpG6ctbwojm2NNWN
d9vlJzU7rN4TnzzBNqm3iyc5pf60KXHvb5URHk+BmoY+nbJyXuJRUQqJlC/P49UHlwH0FkI6IL8r
tlB00u8G+YCLSWRIoosrWA7xn7Ld8cd7fOPEnTL72wyHR38AaRanxyk4dKhE8cQz7flfIFRlD0pY
PVO5VCed6CfpHhEzFt8nOWXc51+Oj09MTM4oAHlU81RiJfhccwtDzV6TF13oZC5f39lo/Wv9nFsl
sA1WaNUKsoFESJos62mbodmenY5D+7mGZDAycnZ5mOx/JRBoUC5iTmGBgYWny0vMe21eudOJGgJP
WKG3o15SsthzULe2hZaABXSG1B/ocWv0ShPECe6sZ7Obj5TSUf/1gzU3y0lPG5EGGhfupFuZoU1c
dee7kLaBwgapwrIlsj38WTc5Es1/oofgX3RpBh9IaXXNqJf8GEKQPuUFZqrq5U6TCzMFCanyk7xR
HaCz9PglZfOxLXtls7xZQ6WcczY/ATbsK9Oo2n0tuUM/WfF1nA13Ojjfe4yBw8URKjseU4gCKjVb
47TwSDO8pSrZ2zDa3OY14h9UuIYZnlzOIg6zA2LV7yyIp6lsC66ha7H7QjyLBGuKWyOFfx2wSWeR
QKMN1y5fs1QxMkkRrm42lFilv+iUyYsr09z3quQ4Secrk1QHEQ6fdWzIBn6DnaO7IQLyj3CPrJ3k
lI3QexipWNPc8QseLkWxBeQnHpulMQz6eweZG9OOGEhC2ugv4/0BBnvmZ/mT8KMRbaaUoqKBzP7z
NnvQNy9Fr4GGFu3FEissEuW63x1Vt+dtzWQhCVe22aMsjPjpE4Ww1lNZ10mEGGIPnY0f8TR6i0ig
TYvenynHm1gsVJtDQFR9+TxA+bUIr3mvEULXa5LeDqVpoef+JTaARlbWx/+JJWJKV/5rUJEVhEmd
Z867OHcLsiak661TaxqE6td3dCXMf9COp6kRAc6tKztIDHJHqNMsIL5cM8IYg2rf9WUY12J39oS/
dypZvYCepAn8YrcCuJPCZBemVIGOtXV8IggEAF6VhmJwRCLjm7aB8fb8EG2vozUiMF7q0U7xFJQ9
5yd8LGYShtG4yThF3ru7o9qRxEAgqwa1eFcJF4yahzd5SlxvXu+MwL+t0/yRLhVeBCWx43dE8nkW
Y0CLsOm5MSNjAON77u/LWlPmyBMvH7BECeGKG2aLOPQfp236h7AEQrj/tNIPLCwbLEey/d0xrlEm
YyLRYQaJyOyOu9bcfXJOIYtuul9/OPZ4dVUN9gwyh+3k9rVePmxSpxwn9EMawpYIisKoargnOIwu
y2EXqHcu/Gu0OCexeQVLbiUJQ2yslBv1BwhNyYz7n83LK8hfmbHywHWXO5n4iGIZlOvo/sBXMdDs
lIuETRGKw2nx9bkp+kWCCb262sNweqjGLGmpd0RYKy1mTGIX1M+VD4vC+lgsyVidKxxa0RjiJRkH
VL6UP+fNfkvtQ0+O9o+4bjLKt746f3kCZ7b85Me5pfIMs1MiUIDQu3D1qfqqh+8IFGxCV2ycpE4L
ICdwXhJk5YG1R4+oCaYZGfH3qdvpjNooCphPtjTaUFZLC353lrI58Ds4m64P3KBnhpHz62dtwjpx
T/8b0CSkuqunRI2iqOFUSpLswXC/37wffpSp09BuEIGeI9xLNf+iXDHcnt1uQyssLbnetTDCeDOt
UdFLumX6Rksb74mjN67kQjJvGmAgQ7pYk7aT5s2OPHHN259RkhyJF0ImA7UTzA4NDmYIETc03vJj
itTk26g6eXkdOkL62O+GF94EomvEh5yLAY+AU/k8vWxGI6xGbW1JPVE/0RrAOGXW5zXkRrQMQ8FU
uDUMCfBFCIkHkMzxhfssbSwImEB6zXE6G32is3T+eqDqceyIDSkUdMAVxdHLIP2Cf2T4A8iZmuDy
e16BTiOpR1NJgw6MyttslMYfBX4tHddNT7b9Vae2G4pd2T3qh7366iBHDVKXlydLR0FKFXRiLopG
WA5KJ6oe8hOXWAs4aX2Gvv2YoH/J635WJSZKh/g1OdbOwfph4afkue+7kUDkAOzZjv1q5t4aj8wF
qzt2S/ozeVzjwTt/iCqBgPNXqWO7eM3+VV0BJ6sdohUBuKUzI+/wO87PLbLvv0qZD4mVc2c4/lU0
QTG2Fdbli/jSguzhaT8PJB/aypGWw9veo6XuKeZzyTQ5PtnK8unZhaHL/4ggBMh85R7XmX93FtwS
fd1xWrFwZ/zhIvfySS7UVQ94fyoP9ESO3yr4XyKOV9oZOIj4b+uaMoaUOQCVHKLo+J+Cpqmp/st5
k6f/Nty1CIH56BE24h+MhAm7+BWKxrb+1k+eh4Eh5eJo0C6aCwLkasXixcItf2+LIYyi0UsaRKER
cfUUxld20tCsIW5uAhe1xqq3m9nlPn+VRKsirh2cKRyE2q6Xt8e38LimVJHF5Zad/x7faZ7CEMHR
ysQ+kq8qvsb1GCEVosMBc67Mpf44NIFNC42Px4zFpZ65UOuvst3WrGV8xoRIgiwM7M038iOCrfWD
2sGh9HO4NattEN07cng2H+5dBbHf00XPTafB3WokAOsoXgiDSmvTNq+bYt6+Gnht8risUnFbGGdn
/UoR9FF+yYSar0p5l2ebS2wsMVWazMx/NAyzLgsN4SBfrC50dK6y6Odd08gNvp8hqr5ChN3CeoLu
subiOhxqLz0s+vHU9q/IA6cNTH8llYPzzUnNHTbJ9AWr+CXsuallMeUKE+mT2VuKqJ0Q8fBMiT1j
Wl6C4cHquGniD8nSDuKTrSAuo221N5xv23xv5JA7skVB7/zyuEYwh1uPVz7EH+JIbgUpLOyfPVrd
wkrh+Tg4Fi7MXOcH3cAyR6GCuU+OFuThdFIW2fbiEb6874AFq1zRUdFyZN2qiqjBhyHHj9XK6vFU
Yy7OY7l3dNyLHqhRnHlIVk3KFAU822XsrchPtIZGtViq7ZeQ+S1bJ1F1sDHW0wpGoVfSv//+EBUP
o+i8Ril+yKgkiod2kvg+O8q/rGXW1rvmjZqn1tf2zY0fDKnyG7/4ZkAdpU/cbYahDqfkE1tLNFB7
McAmhMJXk4vc4qrFp3lBr27DOch5ht3QjJ5w6kHz/3anayTPKungdcF7UFGUnRo5tsrDldusA9GE
2v4q0RRJ1pvNhw5N/L9dhV8kjn617C8h4N2uQ8r/mEnqR8QbRaeN/8i9dxysZt7bGYOak8vJyGeI
Xfv1LDungvYDzuVn8oMr0+6HnznxmuNuoNBuuc0RviNntcBMUVEPpMxKdvhy9dgLHEdD9E+NN+Ut
u/FNy1Saylp0olF0OzcOdr6huUuxIES3oFEhvErrhP/sdBsW8Ia4BnPhXiianXqg7ZbnxXc7rlb/
qSUat8K9H4VtkuOUPAWLlTQYwZ9hhXEwytzNTu2cuY6R8t0ug4ZQOQ1xaEsm9680v/W04UV7EG/L
FVHnQ2GJ0Gxk4QIgQnlzBi4sVK/5j8o2FkNvKREKJIdkQadIKmgTvIGaokqW22jjDW0w1R/LJ8jm
C/nd5pfIRsV2bcuDEna35x16T0xo6RBJByMF6j8lL9tB3QXdE3v+2OkwxUwwZMSgsEgkh/M/2VqM
NiDp9knrxkKbLX5J1HAw3o3bMgng53rAIwzhd6+x8zI4XSnh6/ipXI7ypjnf/Ft2DgbUZASjiN7E
pkvemuCapUzz4McdM1LfEEuTvIAI33JnPYFXd/GBjmXK1HcJj6ke11Ujqy/Jt6KZOyfw8HB5Rt0N
BvqesRKHkP4Vyb0pwAblv7SVSrYPot0vjgdP0sRWX4osPECXy0oanQJ0Mnu+OvC6rpyHGij+cLzE
GNujjNuA5GnXlo4kRnvwutggTxFs6ovRdCi6GJ6GkTSuQbCAd2qIDGBVt6waOGJeLQFV1RrI2Gkz
U4DVRwoJjyaFqBAPQxQmfNE1ChHAfWrXaVzIf1Qta3NYAeGyCPGtlWLO86G5tmezyt9bSWY5eztK
Ea2YeUXHgf4iUpNCFlft1UpgEu6FB51AWnlr53tt9qUdPR7LdJX0krIu1lV1PV4nk+47Dw+ndPYg
Qsgv8UV9WfZzwXwQp9+LRm/UAIYSsoy1uiNDT4aINn+28jygpW+ckijxXmCI/zATBeROw1ooPqTV
Fx5TgA7CLsoPqml9MbruZ17LH51Wx7A2oMN4Z/fsQmuNrtuunRazOUzbcipne3OLhVmViyUgq2n+
Mje1Rfzm4B+T5FMiymRw148UN8XAqA4dKY/Go43mPC4RnYOGKAn7FCjfyVnyQiy1aV4CCFV5bdNH
6624R9btqtPO/3g9tzz/DdBmmv9qrZ++WFQr2vwhQrTL5AGFStbbI9WgDDbepLApZ1W0/rL0I7HI
jzl9zt+aC0pWpV+KDKsAdBa8Ea8yHQNRrVXQA0wc9D8mj9q3x2GYBOlXjbDFRldOUkFmQ51YRcAh
RBh/AMaKX9exo8R4jlsgdh5+s2d1JgDfKj0fGO1I6LByhCJf62sAXuhU8JUNZWzJEMx40LFBg5Bj
+fQV3FXBLGqYfnvCFFRaYgt1TFF3s//n0VAED+z9qSAory5JOVPChtTv0/6BpmsRYmwOXR66XSC8
WWawJFJJrfpuB7SiEY9RScAP5xu3HPkNrEhLgOpFMhLGyC5fkZ7qr/hPKEOIi9Yq/QERO89pjVEt
YwleCSEG4TwU5gO3DRjCTK6Y0pRZwnXjaoC1fhXtmGUWCwp0AG1Oa8wXHjTXeNDf44TBSJblP1gi
J9IeD2K21vNkMBNNWHOElT4bXV3/6ZZfBHZYfQ4IF23lv8CkovOZAPEm/qVxZbWbIvLJXrs5X7tp
KYZi09B0Atr3DyhbsaVZSCixD4pX+6kMvOyPVAbu6rNN/S/HcrtLwZSJIFZMRp13cTDQokp01Vew
76VPkyJyZkvJx4k7bl464qihuEAVQ8cqsCcUW4pY4QSF/4vzuLWW2z14gwRMQ1KriiMlMM5rpv8m
QHmlfJh87BXqsAxbRYtvoU7+OyqfJKgMsuRyJjcXLLGhLT2+n+VVdeoawQkSikU2qgltNwkOY/fA
Tks0xqX1r8Nj0R6oI7rcbA9x2rxgO0CcZPNXdhXpZFlrGk8CJwfEEq0qvxIWOWJZnSEAu/ABx814
1CfesxizUAC4wk6bTZZU4SC7Y8fGuWcHi8KId8sqonpBAyfLiEMDCKp+Z8/Hz4Z5KQdKlMNSyczP
qpCLWi8rBSo6S5rqO+5Ttl9BR/DkUwWWOQ1jO7y/dv0V0uhYQbxlBzPGPdogXbVuhUfY7+7nqh8J
xB0VQc9KYiG8kdnRukYpqgsmVUV4WESEMT2hGdvur3i0zqlVWK4Xn4EsaZhOhnl3Fmo5Agg7o1/F
JK61GDE+A357AKKofNyYtIC357zT0cZyeDkjqET8FKGCylYcy7pQeUGugBaMyy3ZWk9Ka5XdIUT9
tgv6SodqSeRLyi7WYtdDS9Qht+3ikYQynFzJ7wrLIz1lb6qoPMBNLUm98E8u/IQoQ+X3I8frpxBY
vBMTFpXX7UlAEM6KkLNy5pr4ttMkjSFZHMKXPuCL0Tgb14hplUjtXe3tAFnfM1dqFGXOY96gUD0p
aiNWlT0VggOO4eJ1VuNCpcd6MLa57E/s6TaYJURAj5Oa/jlFT6IwBbl8KWVBKw2JnBSaYSNI/SdL
kmL+lTsy/rSyWIZroJZEfGCJz7Md1EOfkhG/YZxc96qsj0c4NH9ZULsmrM31BoIULPrK2COTIwZO
tGvzy6s/+cOGn+YNCa6M4wBEcG/lrwcE3DlC8pFSkcaX9o3SM7QUOMv4zM/IG25s6UE6IJFWySkq
0/UpvJwz/QM9EZWC4dqWYNyg0kv6/TITYHuqGF7rtnhiyUHA/U2wMJI6VRmKHq/lZnncH4Q96BXu
x9n+Yy0qsfljdoJ7GZpIPegu1epvkV0pVJt9I5BvN1dYf1hKdFzP2xsf5qBgvQW1mbM1ikoGEy28
zsEUGNFahqCNre8xdqRQehPdd6ezrO5HgS5VXvOiodfsnNRhGLimjaGvk8ODrYwUS7wBhE2sqacx
M1hihx8i+h4Srcxu++GrlTcWR9xFICs3hGiu0MWIYtLse/4Gy/g1KT0ruppIlDPtYoSDZzNZj/j5
1+bZ4Sdy8PkuEt+3l5tsgs7WjcRJj0fr/YopedLKW6Xnftz7v5562bwR9+Hn7P9EJoJBhKifyTK/
5YarEATMFlfcPV0m8L9JaW2YHZmYOw20yTfjbsiLvAB0voGAXfT2d3h39iQnvxVnmkpBBo5px9E0
qkXkQJ+7teibQe+hHnRqNRdyuqzHqGSFYmyhx7dFekseKPal1YgZGyTIVGtX7m6SqtuBODHzhXD8
ishj9tOnJnD2mHoBeZsrJTW63XzVcP/eYpI7wrCSkbzvwbFlnfAaKLCzUdArnmSdL6LZ84dYel9w
vlF9wjH9oKCjzrwKj2x3JcsdbX43z6wDZ7mNHfKFTxV8UM+hz+pvmtEKhLBCyco1/Rv+L5T4uwCY
IPnzkLb5imrwW/9Cs2KgqqeiAgkOnSH/wCSNlq3q2jHQn036S300OCD2nTuaVT9sk5A0khiWQvjf
cd+IxfPshTulCVd+knhsVSTvSyreS+spKzMEXM6HIaI43IUrGluciYLk/wkr5Dr4cx5jBO4lsCcD
gyKK8RbKV9K7dXHFM3jHHV00P539PjvYRfNHWTUIdgYDMZMgh3P22RVXHeF0g9PsFEhnrPpn26ng
3V3FHybCQn5ANUQf+kLwVb3XXEuHr+GxQl3blEvd5lNWDdmr9xsRZ1wIN3Bn08+YVTQsF9+x3yTs
V+PUqcD78/ej765npi37R2P8r7+4skHrgD2BBm8pxM3PyHCugYLpGb4NI5x9LSxkgcaSYtXaRZwO
/g8JfVNdjsUtdISBzO9XNIn/1H2t2xRKh9i/4QFYXjF+7VyIeCzrrD5Fc7HhfqBbIVcJQj/haQnj
8fj81QA6/DOzKcSmTzeTYgnW8/vQiiFF2T/uq1xdAx8eOPNfMCcH5dnZRGt5817deUxDo6vyzfXd
spe9+i5s7N7M0HjPt69g9YQzA3pGTVbCe4UEwEMEeBJnXk3DMfbTl0kJXg839O4TT7ioOunj+tOB
4/s19Ip1YkOP/fwTC0uC+1fKSTXuej9StmYdUinXh85xsbWuA1kUi0//OZfBt5CHy6AidIBb8AAq
Kdi137U+tbBNkC5snZ5+3AalymGdcJMLoFM19Ls3r6mh/2h/eZ7stxfPVSeQlD/PhsjWjIoFSBG6
y8NA5ApF2DN4VrtYdYZ8ojJh5Xsclifkk0nkBo4PVay7D+rFc84JsPTpDQWK2VsGSlgNIf+Zh/1l
+Ydj3yKjSoLHPLDxhYSZEEnMXxgFTsEvfTeU74bE8fgyH4wGGRXZP/490F3Pns2rnfChAOeIYVOT
UdPkRBO2Y+EwMDt3pnQsIBnQMEheD5bbcvSLAC0ty5rHdgqyQEh4dy/MzoEACMPmgymxnAu93q8t
a6w3eywtlsCdJtcKCqFJ954yYtZM62ANRBEYVstTpnr3HTWZos3AhupP/ejDMegS5mCBNVgCSkjO
qa4gu6k34otL4sqBF0AZ6YHc/N2VBIs95wMsL2hMK+Y77sdTIgstIFO4Xm5SC1LT2hICwoohH6Pv
RiZb05U9P84Xk7V/msTgzz0WpT5cVRikIlsEEQRTFZjqSgmQChvYNmGkfynKvb2FT2gxIfpK2O3v
o9HVFYgKpmGOMvSuziaLpRgWuoP8Kqd02CTjgKBBdcwKpWgXQE6CUqVAA/2fYultLSwKHIrgmnL8
0XYEWHquYjpScafThHdaFYba91enhRwFF0TIfw59a6P3Nhgg8NVnClyZc3wwTevuy42YdZQXM4eO
MEmaBazGRxstWv0En1/7iz0EYiXawS8nRBCVoMrcRKsVrMqyxLPwPqLx5xXseQ9Wud4oxh1S9dwl
mbgXK8iE11jhUOnix/hTnA3fJy/FD1+4YxruX+/Gr2XEapZ4i8EwiSjtlKtHKW0hRukHsai5Zca9
ox/Xi+kZK7eBYL522JKaj0Fp/ih3EhzO+6sh7Ff0ZVTo83gbt/VL/yggykqDkR/5DwvIQum2X/Qt
aCwyYU8CAWlIc6JdKn4ZC9B9Jgq5YlpVOi3WXqO4DzT4mOoRePikS6GU09C+i3C8LgXQvemKhJdM
+0/2uEyeqGNoKkYBc6Py5lPajnNF6cRorz21ySGC9c0Xa/8BLqx3IDIoGANn8aiwRdWz2gbfB4iW
I2YHE5XfsOX1yGW2PIADlxJygVstWWiWOHeTBhkePJ6LqMkx+4MqxvJ8rb+yLm8Sg631omzUWWkE
B3cdweeDWaWZ5h3fzdpu+yNFeKoQ5pfcV0z3GZOMtPMpnAAlgmxLUhH2Z5oaellqk+PO7Fs+yV2Y
ektHW/ALFdmV9CGwvGmTxxdE230uDpchbwHsD1xlhS/3McGDK2s5rPdf65N+Xze2C57PsqUfiGGb
meSva+40LDnHx7cA1GSJhY5IuJ3+KdNZFLYFenAW44TFuuvIYT8nKFY5MTBgq1kAPZtWCkfYMYEQ
p7evgR7EgVxBJL6ooALEFQgfc5msJNa2s7Ag5Vi5OlXy0y84+Z75OcF1E1ugqZ5MemJ9cdP2KhLx
a83KSGzaC/DCIX4aZMQVsZRvE990jhYbaxWf3O1iK3TYVtD+tpd7id/GJbHHjC7oV1KuHlBzjBPz
F1LHkJlQnk5PLUpyg4q+uaSY03cJk/wkNQlj53opv1s2GRaSPwcdlHCM+t69yJIeF4O9U4gRR0+i
93/b1LBo/64Uh4TWME9/4WVFuJfxbMydZI52akUsHx1SzOnnY8rwpFgHbiXex7PH2i9r4kf81M/7
mTnCWqSoPXD7Bmf40YTtZ920HdWbq4yRmdu2NQ8rsNHxQ2pU4Gyzqm0erJWQ/0NzZL5Y55to1HS/
vkxWT4eCack/ucyCptdegVKGIRwssT5RzaI2g1gcKWGn1HriVZscT3TgeGyebx65Kd9DfxADa8Am
MOV19ygsV2F473p8itBDdd0P2s8X0k+ZVOfdAP7AeCR4KuAZlR/Rexy8yzxsYKN9LDNL4dma0xkQ
VeI4ldSoeawn4/+7w2rB4+mqLQI1bJra/h+AClkStYmoh3q54DZ7+vp7K18aYpBUfnHeeMmMRsLv
4qgZmTqGDAzBeYaqHQKE9Y00bIHvG8hl+k2pDpJwkKdf2N/ZMWhcLO+fSTCxThrFlleNQAtX4134
DbtCQVy6IdquvvqxB93SNjYqUN8Rs7+pHpdj4q9usT/yp9xBsH/QEzd9DLsJH3/no0eNZtRPgUbh
/dWy+GjGMUP0P7eeSL04op0D6wQglt1KYjXQa1Zj3fnX4nADrv2K6Fp0R2jhyGEioeZN7ivzGoOU
42fCS32bB5vLq5Ixw8xnLzH8VahvqlYwQILnEVh04bGAZJFVIl1RbMm+LoMs4ZpnylFAGRUWnxl3
k/CZYpozh96bpZA/CUbPmmA1WKJ6nqYky3gFeJWVMg2+Sz+64JPBXNY2tR2hmqcaaugvWKmAosj8
DJkp9V3WPMLb8yOEekZ0oLWsi96TFNjAj0xEO89Oq6UYrvqz8IHdltm/4EwjOmQWwGHHbXUWByEU
VlnFXqCQSUF9eHW45/HvTWhQIxgSAeUsIYoIsgsYUugXtJG+bhYj0FIE2bRQPTtgt25PrzeB1bCB
8XZS26Q0iLXPo4n2FZSfyiNk976ceFBI/w1WsNdrxheCQkrQbYoqXQSpIBjAt6JoxRBlMDkgcl3t
bBG6gxDOYj8asNlG0xHlw63BxNxo5CSbHqsJmitT0a2MvGx2ITCZ6yEe9CmlJB7FUWokc5ChAdaX
/HyDR5kfpC/+PuDh0TiLa1Ue1rNKVzyp1m7EQdSmzq+np8LP3CWHX9KX7WIt26Bsysloq2lrbcKt
33pkJfrRSIrqERE3gjsCqabifyvxf0rzko0XXzjwMxEd/mlGxafiXI1kbF7vrihiBx+ZH8ptCKit
PeqjTY0xb6yJ6eBvH7i+Q4G27zmaktURPKD+BfX7SCAcFM8JqrrVu1F/DmUBGULJLtg9Mzc46D6n
YxL0Y/HBWxaBUxG/AcnnJnLhhEPFvYRzalG5UMG247wKCmcf+ttIwb5vFQMIVyo/BcUVtyh3dVAu
n92qDX1OOcSwBDz2CmO1gg57xO8dXt5j1kHEyLr333dQ3iGXiz6czUW0IBfH8X73jkeSaVUKywaH
e/KgPcMEq9NVjhwyxy5t/2G4FWd/fcxwPMrwzHuUCD7WEXJl63l5saeL7CtQ6X/JHapJ+D6uS5Y3
JWKS+rbEZ3W7UJ2Yaf+I68qc0NS98XkHfL2aqhl4mPqE+4RAUzmyBs+k8nIoKMcuI/MrCTbX3r+o
wK4e+8vSWbm0Ht5+3ZDJ2Nshlm01+xurEhSk1cIFJvvsfoxQT7FkN7nlFPffQyWh5wZpA7aq7y0p
J+eUGU810Bsi3QnI/KJ2PHiRODzWgJ2ia4NtN3nN+Ykenxv+C4AjZzWV98MOtCliyQjfsGURifQ8
zp9mEg0TqRnJiaqgFpuuylkcRnMzQbfH9Z2ZOC3Gs3zA/6u8WfJfxbazoDq5CynTXmMT0UlAHNsA
6FxqiR0UgzjvyxB3qpV8a3vhOtd/vk2nD3mm3iHfddwl+H1u0HacLShK6QUFlm1eEdfiieMaRi+E
keFH751xnwlcoX2oqLufUouDBBCGAUnalbn0Fv6pUc+R2KyBvk7GsyTjTaNfG/WM7wg0CCv3shTC
MxT240KWesk8+NRKbyLS2AgfqtOs+A8KqosHvYYHs5owg7WEXnguKawSj2r+MMogof8VV2h43td4
xdCfnslm0kPFvv3CVy9T1CIAdPS6kuR068J5SrPwihA/rT8hwHGOZTYIOvE6wqp9w6AEoVC9aShM
HepLWZl7pe3eWPVNeXG/zRjpWr1gKKru2Dh7S5hY6b03hhlcHR11N9rtq6UanoGxVIWfq1F5Zg+l
B8mwD5aMXOf4MU31VSc7AFUQBmC1b9nANtZ5I4vFuKOn4z7ydGOXu+mfzdOHwAkHPIhEGM13N5si
okM4+XARuyHEoEPgverBWANZF+GWhSxQaiuP3ZezwescTO4ziExe8KTYuntkOKyGii1rUtC+UUNT
DleXfJ/a+EbRUNI4vZmqBHkzTXycwEo1UumHq92WIVTMyC9NEVHWsieZdXI1KosN+X9Nj/QJS6Ja
V8XtRgb6h0hhwW2vYi5jqGPVWCvSbi1T5L1kEosLLFxINvdjp+cY/ygK/le/OkmwmrGnh1ke/q8g
wzSeSKyd6QqJM3S2GZeYqR1s+lI0voXJDLg2kpYwZt4GR5FRrjFM+xwdkqi8qVq4Bq7qSoC9G4xb
oABwvZbXpXKm8G5dMnj7Mu48Mb8tucnGTNd5uF8MDl37dX5X5S3LHd9/zSufSPXjqKPXCDDDagwO
WnqIXTNVcqwHDN17UZWRjBQQGHQXUDg+xQLfI+KUt/+5VUH9nXUAcYcC5WEEoj6OlpijW3r21EqB
rH11I9gXfedfUZDFpqZEYMZHHSu/x8opq7Nnv8Iq8vLmklHft5nzDQh2hAfWEGmaquXbWCYrKCn8
FeeN9Iu8Jdq9xqk5TCV+2n0wNdPUBYkEG9f9zCBaVNdOSQ09WE6MTKBsgoCMwFRbr9EbkQkOeD05
XwSWhFK2wf22Z4MELvuCuz/Vx37HkZBuVLdoxweHq8hJCdJJfWdHtPU4DZux3KxRQgW6AQQ91npS
eZ7UfH9aCRiZiXzNUC0M4rI4jr1truEw/sUmNdYwT04GUvvvO4VIvSvC96haUR8s7UWPRXvop8QS
BZpnnPbtXORCohpwzaOm9BITvPRBSUEdiKfZtj5FET1N5dmB31QqRGSM9GG+a0ZeUaoKmXPHhRWB
Y3SyrAv6Bq0TmT1amyeeF6l1LjT9YE77bNq3veLM+e3Ik5XAA5Uyj0Hfv/+2Gwdp71QPm+QOcs1A
9XrEUArHE9WdsJIGR/6BncYG1XrknPaTIlNG7aSPSHrr2c3at9s2G/RVJnVfT1RT4hzC1KEFkjpd
AfFUNgl9WQyJ2NIOQG7mywHRPTTLRjI5gcds3s/ifhbaD48XlCnvzWiRdDS8dU6VeD8Z7SSN9W9x
aCH8IBaPf4vvn1KQmwhiAWP9e5gB48OvtXFHHlATWah3JmmaY31iFIE/CKT1iL6I+yPRyYRjrvC6
6I1uLjbXtbfDmg9oO/9mQBIOtrO+zi9s1kKyhPLqKfG+brtGwuA7NNWDcaKuVSogXSwzD1VoVXYx
19/co+9qrsGJlI1aWJLGEQM/oT3nPzdEym4M6ZJzlT76f8xdIOwRqiNP9Ehvitd4kbGGpoHk99od
qFvMV37z7m3W79yyz25SDJv/MHkBuKlklLv1Pj+KhhNFMUyLY2MW4o/rcNz/Pi3sEtxYcrbWgM8B
I7V4hzFueiGawHtcAZ5Pvte3q0YnCxjqvSHV+i1lV2JHFPlEMsOCY3JtVSiRz5NG5e52HAS8uZBD
N6WixNeuYSkrJAw6lKjEC0JL65/n9hk/95pYK8sJsAJDxKxA7eiMuVfItsLeNXZHcS6vZle6FMsa
HdsmxUWhaaiITYiJyBoJqBo9BIYEfNkNCJOuQQVMeYz5zeWr+RBQiJXUbbCixJU7mrS6WCWiZc3x
t6J4WYB7NWC0nFPtma5nlp0QpQTy8cDiMckBpuOz+eI0Wbbc2EOf0ZktraC7bt51chLZOiBU0jJm
f2RhOw2SZMoamgvoAZ4e4VyQxTQNyl94XPgrk0I9BDKrfP57/dLYQi+uDgPm+VkD0K5Y62mc9Jph
qrCc2TX4pkKDKTt7vTCNLBBWJJbGBVEhjzZ1hJZElkguyBs4PVNUnp8OoU+XTL4T0jlXbG42CDhG
C9wMYqORBhNas/LL/8sRBxoxz4FLEvkUXuA/VGdN5tX6zARNOzhf7CGrcnt0N0L+aOfU7s1rPLMg
xiugl0sN1TKnYfPDIM6njIchWFuc0Py4qqM9Tx3VTFrovpEDsH6JmUduILs/W2pAMUHEy+0U7qmH
/kC28Iat53ZtCAMzDtlUlMOrkrklY7hNa2wq5EfR79YZToGE65C83n7sd4omaILlvrVI+8mDq4KA
+M7U+9kNtTcZQazXxYM9Ci5CVW0M4jmHeqHSeMYUoEXtsz3suHkC5cRs1DPKqqynAqIdrUtTyo6+
ldWldxqRP5xf1ICuQbY33uOF2Tl6LznjDbLlMaERWBwR/0Pw2QbCBSN8IiJTG3tMNVLOQn2JfYBN
5S8x6w4b6j1pPuoMMJgeYmYY/Hi93PObDPBs6Q7JJlEJM4gWZWsIUvaSa9YSCMXyqqBn945WD2A+
9h1AdLgX1aXAj7Okw6B3eaGZENyQJXp68N4jZRuVnHzi3sNvBY3ag4D/+k94oSw/uGP/lCUOW55o
C1IFxU07wW4dR5mhZxmkXsLyzWCSAPjW3JqjSFVITgPF4/5KGJ7afAkr389YNjN3dxoKEM7N3CKo
pbxIMxckYAIEmPNOCPalx8kJAoPtZlBvQ9wt3FJTgTsXX2vYzC86rv5P2GS8fBkDratrirkpH9B5
f+Wo5Gj7EllWaN8RqdjRi34J8xh/MTwwU2UNlFJDP+co/qnENdh1qdu3oCUj/UnYWhnEuqVGbCUd
pfVLAE1ZeWd9AWGkSicaz+efgY388x6XE0cMRhkTy07n6KjfbQCPh56P1vH+kiofYFPS0iRpStzY
13MNQXYh46JZM9EErFI5ruhqJ/+WONn6b22se+r3DyWgwWNGulHANKbflSExfr9BtQImYZpYeYfX
E7I2dOQbbXsc45xjHitYHFUohZAcV8I4wQRencsjXGQiKCF2IShrH2ZjyusG0aEiNThMaU0PMeqo
wOYWSxPidDZtGUT2EctegQZyPSX6oIto7u3SrO2yMozGn/122tJHBfBCDeEtXtB9z8CPFHQQEbAU
3BxDvdZ1vQgsIB9tYM9c/2eIAmSQMyB2PVINSQ6TJDZ1bq78vvR+ymw3pWdHw17mINkDsymaSbgB
Mp8ba0R2MFCYGz6UKoE7sbb+J8xcQp06KcQQAQJSfezdZ4qd/jEBhDt8bLlmdrYkz8hpJ6nHImHA
xXJ9NfgVFW9gDmnOlmVjUWbBuRA3OmEov7Rwpr7P2pRT37vgHdH/xlsWfVFZrgPfu6ujxvEZ9z1o
htYZx514XbnTLYY9SIoA/wutucKATBF+LG+KaLuKbex6xv8dJkI1t2vnAK692ApZXzePVfSeb53d
Mrvedn5WBxcDGGQFNU+1VluAoItOgSAT/ls8yZ/6jx34uUXCD+tE5F+eIVEVkW+ZiVLsf7NSxQE3
pBbdHTmDSpxVyAL2fcR7qLXXGTzLSxfhcF3c2PxfOtprOyGq2ip7+BYXpS1vyj+XCEKa4cOzTiqL
sPCZ3/ra6fKR99bwGQMOYIhU+8Eg1JUaKuOkVS0vkfdmjuSYPQMCeErsU5JxUPYe8mFz606+ZAtu
SABxQ2KPQHkNZFWfICYDK9PEPny9n73BzCn9GQivz8rrxDIk7oglDpFLvXK5pgMm49Fi6OhDmHZ0
pcRqsVZDxlQge0V/fkgYU+udMZ3bf3/+3DJ8DT8jp2QeRUcVztf+AkQPt0mACwgqmV+TvWOf6sYn
4gI/O2pOcLm5ttm313UsQYLMkz/M/j4CjKA7x0vsp/cIQL3q/O0/h9q7hK6WNtoCI4vXvwvQbnDg
XDyUzc+RKScaCKzmO4VAdVkOnt3P4AuFMD36DtSeYnEDPvWMVQsLZqoeyzObkajqrufSKlJ06pcQ
setaMx08nYIbAFXZRFD3PyTbJ4Jk8+hMfgweRP5XsMO78w7HS0FiUhKi5ux5VhwVFLCHIC1pJ7av
i+oj+YflaX27xlDfJ7D7BTgtm53o06HjkQ9JIWYtjHk1+F3QW2dVF4+bLn5mF5R0uTvEdnrS/0X8
WARxHVAqnR1ejF0KDEeH7xHc/Eer8SUWviEOhyDD4waDVV404fsw9+Nsnvt0CsS0s/Gr2S6F4qP3
AZ0hFuZAGKklFhEqotu+aeXrFbJaIW7HC5AkpB8lyGPkif7hogGeLtZLeKdmpp6EhC1OIocA9xz4
bM7E/fmQCLo1PGV6dd1rhO0A03TqjVlLl56E333DaHwBF0tZ1zcu6cnkEZTNe1qyE85g0VJkW/92
cXYzbDOnG+W89wW79e3vw0N0usPO13+/t0psE7KXKNQmHlcjafdyvyvt1bZeGupKPQMmdr2KSstz
Fxt72EAIKUNCdEfYkTN54TCGlPYCdh+xB+QUz+yxP5TkGaCD8Z42hh1+wJQl9R6HayPH/7J+jpv7
CQd0WO8y+wvyFNX6Q6tojvPCHrNZASC1w7yZqmzUqFwSsJc1HzfTE3xbzlhTVfMi6rUhKIpRIv2O
OKoN1TfaL7dyHzkr1WGexKdQVJEdmsTfib6blZd7oeUUSe5RY8KWsaNWcy8fN45BhwzrLsDWBUc3
p22kz91gGCC4hlmGhc+RMXJhWsV0GUz+2qrEoJevEPo4xogE1atXcggyJ7BKQrVgmCi8bPzGvDn3
G6lShmAPs3w/donGC6CPN/2NpeZQwMkJR5c+yNBewSdq2eP0VW3IKv8Nofn8Ho/N1j0CgPm+bSXh
3nUlRRfgRk5Tgjb701CHKpQS1gf/qjWMukoDurATKWcAmyUYpNB/QIpbNtckpa/jTDriesrtqgs1
YQeImbX/IYTcyvTdqUcv3bI72t3qZvu0O0FE1nEPGmQrTlQz0SblgrF7RhiOmrsFPXcfaRzSRdSz
DFhqVY6RAtftgaqPqUhQpghzTY//6znUK1WprlF0kFIrRIpuHD71CegOV3kqgvFkElBo5JsWZMtz
tKFOcx5g+9i4WbT4eyBZGyhHOcqqAXqIq8sLlCCGpa8p8FKLTSoYgFUwP0h+WJZHgSJWiWwHXDAY
oK7vOcuiyTzYe3ncPBHNTGLgQVseeqxo2tf3c5HGJihaJ0jNK7rt6YHSJ2IjHSA+efOZpxEgtz6g
6kSGUtjcxw+UGxRA/A41qrCwk4w6uQYN9+j87e1ueLdMzU78rBlpx7D0Pr+94C2p9PtqeMw35Ie/
YX/0/4XKShcPHQsj30Rd7CdkkH6JO2xO/NGgzuZ/MEmxQeKM2l/928pvACryMRDXzlUY6FZcCmh4
Q+sYgxOZhIbLQEp+4b4qRSuHb1oCkOVsEHRoh801SGOi0LUJOh43viPcGF2JNH469ER8+flK4smZ
ZgspqNbWljC42RISEiaRTqM7DKeFeNd1eSoX9fwvqyY9s+DkicygnS3HNDye5j7e18XJ0EH+ZbiT
gbH4DR95OoKUL8cMoufUdjAVAaEeo/j+D0qp5+EXh9S+tv0cc9cURMN5/SgI0g4xQnPWSPf6/6gp
J+S/mfu8iEMBVwn18SWbWrXvvkZ/DUFgfAzUYrwLb7iFye/kaIlcUS1u+bbM/hJhaVQYtvted6pc
TPW4uqhfj86xkbfK/WGU3/8Il4Vo5kDLYUdALk/n3ClxGaFYuExqWgaA58VGTJJkBznJxklKmjPg
k54zjVaSdXhA3N3Juc83upcw5veWRJm4WK816GijmNkK2+ePX5ZN03VFgSnr9Ec0K2ULHsK+HsNK
VvB6zozGK18TPv7S05Jg3FDLoYca+MFapclkWt6umpGXMadgC8mn6byaPGnNgqe70kX9KZ1Vu1dW
no+Edxdv3HB/Uf7a/ciW+rzJfINNMDibvASy0gKCMFg+P26J6hA6HjYxnDlbIq7FJm/phP89rLMJ
9K0o96fl9CPxXBxSh1Mp2cUSFju7QJEPOZkJVtK7r7njggIGdaXG06/RLtuCzJp72uNEDOoGzE/H
JY0YOQka3nFIwY/455cQpqxy777X9SPSNGBVvNEynrErr/NP2IhjsbBbnzwnkFPiL0PUCAbZFNAI
wOGVV/SAashIL0kItoZzFjNh60glY0n5PvtshJuye90j16ezmN6b7EXIlqvHuTIS1NZmLf1hEga5
FsG3WQV22pKCYcbfrRNkVg1Em8v9WUiWs3LMZAMHpn55ydI0Mn+VN+5JjYW1RbTqiIoW/XrJ1hWZ
QTMY3s4CCxj8g5Pm15bDel+3uu7kWGll6lB6HGgrxZAWP2eu6xUbsITg5azhu1ZnaUiKJnrPtf0K
kRb8a8Oy05/OnGsH8TNFrjUqGU4INNFdu+LpUrm5t0SHPokmDtZSAlHz4h9TqgAwoIIAUWzLCOKF
ICHhR946GUYngMPuo81r/0PRN02N4WFNTPsS0YrUoQguuweAAp69KFGbbUv+dzBM9HBAzL6nlDN4
fcM3wCPo+81gF5O9SylQBnpW16FKeveuGvBB9QrIXiBVdI+XBhvvKHLHskzL60hGjhPTZ9PyEspR
Ul5B0bItuXs7Ig4AjagzeYurqhVK1couQs9d520GL4dSqisd9xzHJPZv3X1VXLs+og5qG28q+M4g
Rl5PdDpY7IT4xJi3ZNHK66TIXDpcsrqCA8Q3FzdFTTWmKT8ZfUlSLUz05q7D5BjNx+MVpJ3VIADn
FTVTKTJKGzpzE4T1aKLZnh1jli86Y6dHA9Zmsgffxytp5Hq6qDBrdOnTuBhG/4QRrN2RB2DhO7BP
fVf6SSyxJfpgLRU/FhNntdbAavI7ub8rbQdIXmP/Ya+/sbyt72v0FabmjC8T45pTh8KtpvVTfdvb
j5hIa77eMhcnB/oYO8lDQKXsvEeJNk571VEK6YUMLunZT2PnJaWTlx21o5js/QkWnbd5hCfikIn2
DD8/URllN2K76TlD88zFbt8M1gFBOjSvftXm1upvmq8ntSi8jVGZ7OEu+ApTYiRue9/Gt8tOGaje
9002lRPeOVWqi0vgk7+F4Bf7oj6TXfWXI59ExZk0C5lRVj7GC7dTPtV97txdCwOpOBz7Wf0cNN6J
VP74KdNmds9fxJI28OxGMdY8i+GdHVliqI2nEE1T+6GdckWMCzXcsBza3xqD52R12cA/9WcifQTt
O2dALGlFvN7WRzcsakxDpOfLeBbQXWYczqimziOUCVR+2WKcD/xNg9sbNNcHfhpz2uop3gzCkSrI
0+7zfYGr4gOjYfhCeUqOC1y2SuJk2tG6bpBuqkRrx4Yu2fTBqVaDMAWNgoXBS0atai7L63L1vGLw
rfSnRv26eZT87RS5vJSv3y0jApRK7O06x/f8GJgygKdFpnoFug+DvjdtlPNuzzMSREo2I+dIle+2
QM4W4EMdZ6zm7464OjVeCA5oAe9Hve0QA9RO+1B9aimMYS3kgKrSeNtUM4yrYH6a2DWKD+FKdURU
ABZychZe3wRMlb+O9xPJZxRh5KVLkPdZOUJikDJeRT7aGkC0MHiHtedi0ZaAxox6otxZ2DIDlyH/
pZ6htvpI42KcYfb6814OdfEE1m6Q+HlAmjLNwYBo2hvL3Vm068NMqu2gQhJW3bVvQh/oUsngO3EJ
tPzFmBQpG/tE/wfNvu2mzzYOC9MSwti8uy//z4xGiXumD3vKUOP0IlW3rFeOHrHzl9qkMo9+OzFU
Auw4Wzh/RYSb1n01XFwJMdVD3tF6qxb5/Z2qIhqRRlG8tkiNR97NBBNqMwy22rL/RJVOMHLfkGNu
RKgn5hmL7iHouaVvNEbdblMFHuXcXYnQcZgaJfAYpxysMvnjkIvfutBvKW+c0Jg4GviovPn440tv
5AaC+csqeFji+YdwlnIgywljyuOW1O/lUULkAPBvr71NNFmvI2UGA3rJCx4hbCjmkVCxhf9CQtvw
/1Zg0bKVZEGeeWlpilie8RNju4Mq0/gqdDj1YD3jB8BU9E6g2evx0w1mJoSk3rwACcr996Zxt5oj
PE4jLaAghDkDiGhC9+XOn91ZCbOJssZ2HOAOiXUx6Dz4XH7W9EupVo1qcTqB8P0qSG/K2FPeUIk/
uaXQAI3x2WNX3bnv+QZAQCaIGiAPjCpMH9kqT5w1LKOnkxy8yKesnB72LPCJR/e4DropHR5e307y
ebOGv8uxx6ftdFM19fxVYpizY2y21bXG5zx/hGGjp6hJvoYcRtNQbKsqaQoonv5XVv1O1zd/UlEt
JSO64LFWFMGO0h168oQqHc1ouSNXhR5BOS7sBD2IX/7Q9txeyU4lEXElH05JJ/STLN6CCwiEFu5M
18EHKSLRdOqVzdBZO6QuKh7xn+50d+eO3XhiGjCawy1uGdyh9ppJuNUd2ejTJFRRvwZ5ERMD+EuA
M3pUoua6NBK7cmZnZJavjIIthdcHmk0GP9xkty8SbeqmVH8MHJI+Mag9Unjv5u/mGbpCgzlIkUqF
XU/pF8roX6zoTOl7EhUEC3f0shgqywg7gQ6vZDH097l5Uf+HKr9EbBmndXRxcmwcuzBempG9n/4u
aMjYwM26qdxW1mlj2khXUnziq1LCOxylRIj/ZhKQE6ZnPC8ANDvTEwr98V9t5UisLcyDA7u0XhvB
QwxXdayLCC/hEwkvd8YuPyyva8IHdFmHxvS6aRxtRc+tC+eUQdYmLRTK0l1tuuofjIttu8wru6TW
jLJUWvbckDt5pR3EpDM43IrpD/Lz+K7YmcPKHRzQ9hvbbljTJ1hH5Pcl0L5sQwmK9/+sX/TG8m/E
S2x1pTW2ZjKAneG6ugvFWa6DHGFz02AapC66W6OkK9NzuxuwuwG4vcQB9PB5BvrWP6iIrw1Rr7Wd
o6RM01WZmU4/EM1cNryw84OYjFCEsu1jidaxeVxYM4GWuTsX5i8UB0kiu9tCMSkp8LRAZSLaM26h
gwJRJUld2KINBw8XueduAoiLKk0CMH6ykloEk2BccE5twgbpLTS/2TChZSdVZYYtyQRzNPFL4iGh
5elNoA4k8TwOon1z8uhxbAw4StI1HL+zhp9kmzvBbWpU7TkvJ+j0wKClvc7iPfKiKntONeAy4j4U
JJ11VcC8Ikwuu2Zdq6/GOvFPKUNLSacXdualm7hhSChEPJ5zCxsoP2teSQTbIkSUPI1BAxIu7+3F
N1izFDTbyB8ocm8ejy+P2ZdR4E2K5nr8v8DAU17UkMJuErAZfflRf/jjtrwqCb1/WrL1EZPFpmhn
UfuCeIBhp2Kus6hZ8eeKohLhHWk9BGklZ6nShbXPfCAeBRSufrwMeQl1xKrUMkHVhgLE4u+AHrsd
lothmh4WwAYUuRkCxMHsx3+rNXS1U3hKi1DiZSgyyz4P0VUHWVRAwUlt1e0SjQx8xVa1TwKmKF9B
zVRBsVcqBpcBG+cvb6fRMvhifb46yKoltesdix1QCtHEn4sUW2FJnGZdW1IfU/yvlSYSSfkBMSSd
1O09kQ5rX6hYQKG/zZL1ohq4YH47K/1jNtWK+Ygq/hKHarOGwO/K72frKdWw4Y6I6ITRrVVI/A0a
42BWJzQOI0lLMSEh8WFNNNzOe5d9aTq2x/t8TFBUkeU1TsZVu6Vcddpo6TOUvRmFV9Qp0118sgw6
/2ig/PwSPdgmzFpeaGBcYYJGo1h53vZCQYe7bYoVik69yuaYxej7FhUFYc0r+oEk00uFbpZ1GU22
wXs/hl37lMpLz/HEpjj9ch8iza9p92n7N8gyuo23PAh2m4Kcs4kW2a40U90aQKhfbmQPzyVTAGG3
eCrrLwk35MknKSU/N0aQU6xGuXYYCKzCpkY8fqt3/9jTDgIk2/8v03k9OE/XuRcTx32wHECyvPur
Vh8B6OS/KhTle6QOipI6yQPTcgG1DaZ14aLt/Lg/HpyF9q4lfdG86rIDKQPAeZXyIdR0g+f8f7v8
wOWh2boPSRun1aZQx1XVdgPIQnGrYsOXFbgba6q+gJKLpv710HsXWhkugKfQ2MsrRgaE0oDXbShv
SecsnVpUt/VyozCDz7ArdzYYtoZ6JX/FJZwFHCs2f7Ho2z7Wd1zzwP7rKMZG6qVz6HXk8isXvY4q
NFFYldDzb0Uo1IVRoYwbOWvppgHY2T4AkX7rgzNPm0e6vf//5ppY4inXOG4D8SOWvcZ4sfT8eIJY
175YpdEgLLUhMge0wlnQgMWBm/+R+wOEFr1Aq7tCbKnMc6G0YJC383iwP73Ju8Zc+uzUuhsL3eWa
9RyGY3qdEPTLac26CDv6T7Qet69lnBMv9tF9QFoVbbbEem5YQDuBQu5xD3xxOnAAIt6UNzEU+dSb
blITQ9kBttJ9K5nIalwdeDiFCDOkqeiCTnKpXvKuBpnNCiYDq8JFifG/URKvVlr6Q2keqbwQfHsT
cUstC0KsoGsuMz/kgstoyrRHHj0zNG/Kjt/GBJmHtB7q/v+Xy+PT+QonhgjMMFprRO5R9IfLH8fU
sdZ3U0mj6YIksy9/zsB8aRntgjmSRd6nBVnJY+PilosbjCCp48f9ip8aUUOpQButaIyCixb03Qpz
wGlE8YlAgibNa9lvTvDUEcisc0042xYUVgbv6wsC8vDPpftbsqN4bFZypaGmgOc7EusCi+zK1Gco
Qiv1ExU8wHUhg/+UkQP6hA/nL5zrIihA/m4JwNgKrBglyHVSwJ6YPG8N4W0r0LjTConJZwyZLfDg
UqJfuyEB3I5gQTPhbM3cI33F6XxEbAnH04rbuIrox1VQiYcdW6slzH4aNf09kW3T/zVauAL+PEqa
7Gsd1XTpeTAkZsv9QW4QJQH+yxARaFUxw/RnOyxb457ea6tt2Jlx/jSgM5INgPVrfFvxvkGEA4/0
Ecv9yX+TuQxVvG046ONOCm3qNcUT2PoPDQb+/awb00nM/MHm3lsCjcUivNI7XusQMIkG+dxv8eOx
RU8eyQbTzpdby62WRW4mICfpFtuRs46s/C08SXTbS3M3ZR8MJTUzj+hQtKaYgmiv4BLMuIcHA+nD
vePTWVBf292a+3eTwggyG/OK9vZ+vS0szXStBbEZHlZ+H6euPqsTZimJQUm3L0TUArgTYFsczBYv
2mt95rr0GrrD5HX3IlrRbqLUl4d02wyDGnxjhFpEiXH8Jh+depEdy6fT0lZGbc5CeLCIJ2ZhMkwi
NbSZ9V/jPH30+P7QzQ2FzXhcHyysGYmqHIsdaHz5U2kfaBQuSTfGDod48GDcgLgVLP4F+nTIRiiZ
cBzw2iMXtQf3PDIjqo0fzuR2nFa5Bkz4KwIb2TSrapSzwE0HLmaBbvHzdDtwNItMC3a8gghOvkDJ
gbJvaMLk1ZjiFATc04hh4CcvvpBQyZju+lC8Cgh+GQaY1Hn4RfJk9KPl8L4XQRfRFYDbf472RjcK
9s5KbXociHOiR2A4BuXfgr6X9ZxoU8GcnmKqNUI1Wqg+0BrIW80y3vlJglQZ0eZhXbrV3bvlAo/J
MsBHFEZHamBiVPrZg2OBW8LFmV7I1Cxakmhe3dxw40wYOf2TWp3PDhRbBmgHU6fLofUGY0b+VPZ3
0yK6ZDgJjv18PFN4qZBY2KNSZso7bqvDTsRwHPi0S+GaqjyWSkF4KvBnROat/5uwju6a8A5xSxTk
w+uKfBSR5HnF3gWTEWNTgIufQnUtBR/Thoayk0cTWy0L35VqwO4DJEAgLaNzQlFmVvA8Xe+mWDR9
i2/V+8j8TtduVzPJSrDqLUn7LjHU6dVNbir96pX6yeOsNlw6ISJ3bkKCNgk13+BiAvphtJ1TKSax
pYIXrip8E6wkjRKdsdkh7XDyHvgVRL7r87NepvWiji1NvYfeqmdVzcuKqj4Fc9KVuKNJTja4AECL
stzJav2rduJj0R+qqOP9Wxi+/09qIJbZVgPb4cVYJgUz3C85qhrBY56hUXr0e3oeqlDaeipetbFs
LZ7r/lOpQt7Oo3WASbk+9K0VS6k3L/p11XwFHmcwU7F1EZ2uNrmKTJQpViDkMSxza96tdeVDY7cs
5TFLqFOCrSOp6UY37fp4wG9JYMjJqYzmss4P3/35Qbk20Qd60HxBkDq9ilnhxsvteFGQK6diQEWn
XJG+xITuHnAww7jgg8r4Xw296gvolrygK+lreOtTORAjgwLWe+dTKthRTQGN2Aei1TPerA+3/sdt
8capIesFAUlOUCtQferLnQX5gbeqk8LC9OlMKFUtRvFfhc7fAEgpLiCh7C3T7Wg5WpsFm2FfaeiR
CBZJ6p8/6Bh28EabY7Ty9ww/GkhaJ5wFlJIEKRyZqwYLj7vlN1f2sUKuKhXT6/7x5FVyzTeghKHJ
cykw1DV2Bj5M9265U4c4llJ2KlUzxDvX6s0jI7CmHeemD/rEgq/B8CwRRIEC4NdJRVXfvuGQVfTo
tVy7s+ikA0tZLe8m/iTG4a8IHQjxoP/Zt8LUrQMq7Qbr/de35PNCta9rRKDc6L0cdkm48zDBsEVv
HJD+yXawribEAV8tPvIIM2MWexpx0KJu0PehBcMa+0dIfGJFYPxz4QvOX6Coxd2VJoig+sTd/+eq
ME2FGXObHJg50oCHxaL/xhx138/Q8yZWk/gbLGtpu5jS+9kOIaWkN1h6qzlDVz1zTlARMW6Fqq+/
Ljz7MmZBSjrA3ZElrErf118+c+LnNBi9K/J3TrQ+ENyNgj60IKi1/WfGTzUvfjIzVIn7rli5h35B
XWslqIt6ghCoZ2fwm8DDcOhdR/80SvmYiSjQX5Mat/+kS27Irc4eGFf6X++69Z44oUdTvJjtAcz9
CWuM9hJzTC4AZwJSz9YJz6vcOPcuv54XcZZqEnrMkJdXKw6u0qwCLrsnFI5w5u7XixhHyVALOGZp
nIRGKmcllN3Oe23t0bZbC/vtnCyThTvp5KtZvM/aoTQ8YECElCTQH6z9gfh0dOECeQlseYOtAr4M
wLcIBpvc7rH6W7hBSNS3VqVgdruzC/FeBsv6SiOUCWhJ/CJrgWrMubwqhUXVBaYkxRbeh5/rI/SS
5uced0pcF1iYy/tIsBr6uX3tEV2I/bUz4lFoKbAUyniz/vV0jZOXCDSJCXRSnsBMkFV+yVdlJlvg
/J9CDG05ljvXV1F7xXSmoxBzRUxbTFneA0ts6dCb1Lf/Z5Ld3m9XEtYRaRZUvUQkT2tq9O/BgnPq
Vklf7YA0jeOgZ8P65LIWBOlNkI8fYAsj310E7t8FvAxbYNbp4jVTg54SH+2H/v0VBfsCPF/aahwr
vIssxpoTdPOl+oVDZC1mVGxcQQKX9OdpExUtKEDxzLXRKrElvRQbXNqN+FRiuz/S6OQKlB5LqI1j
EYOY3H5W7TsjWJqPSkAgB+nznOd/eVmkiob8cWyg3TdXHkpnbzcb6BGGCeg8ILhYopBJivZeD31B
l5G+pGrLbIaTC88d1eVEJXIE9nMXqu1D8ToydBUURsCXyvPvy6IQhXace/TJftU984AyoRjNjK87
9KbStl1L647Syz81phNzUhDhVN136eScWduubKt7qi75DQxC7fVaSq4DbNYeGCwVfJi+iwl51djJ
3/EU9wAD2LqZ3OPZvyPkuptKzezVPs2jscTN/6lO0sbx98vy7vjV9R7P/ScaEdozL6nP0/I3wNBN
bqkEjkG1d4M1BmZtdT9rfe9U5quP375AlSNAMYj8Rgm0SRJ5kvFvM44/CghYx8rltndva08JfKrp
Wj6LUDhH41TSWJv5brr5Dl3mUQ3Wy5uQ0vXLkshmIdV5/A5fiIB8PYVYVrym8O/h1T7CVBFSLQVc
N61Vrp70oWChsTM3lZ1dMBlYKAjdWEYptC+oSQZ7dcNS+HxWLyyAYL/Vd/T2PsWvyzSun/TmUgid
NYVZePn66uIFR8CpNDhRAFrKYmnnkqSCcGkUFiANLsd0R5Ol1qtUYsu5XvtgflmwFxT+ItynggrL
xvVhiwzpeo8XhvX2lNtnV61PCl/g3ywpoWSmySZ4mi+mOkF+mVot/f+L+id2C3/oQWEHfZnfj/jj
Xx6ykPPDTkvkepAOOJdryoeyuFr7MYUgdbL5uEtZwy7LCZ0ldHf8t2xyUl2uoJcFHpCfB+BvgR7a
BMcFquyz4LW/OqmV/v+UAeHKTwNSs0g0dUi+f9l6IpKHfXdqGNPrYU6f/EmTEJPcV0eHgiYY6qoc
1/axTE5oFFENBy23BZUFje94patRXka4NrmS1pRxroSdadyYKI+f6b5wU1rhUyy8aZRD/Z7hYcYu
sKF2r0wMPlx3tW6K1yjBjj/1+9Uj2g2vGoOs0jyDQBokGROm6G7EGw1dRh0QUuePSuK1LAeJ6nma
PJWvWlkh8nNZQRKQXlmJ3o658Bcn1d4TTsmwMEyyxbhq3RIGt/jYjvGpGLmCVGgxhsPSqbme/SSt
Z2f2WsOF/p7zA9BWhmkbAREj2b46CNUAAekVNPqoJUC8scxY7qNePnP+CfcUMNRCCOy0OCoV5r40
zBXPZY7qh/XTlwf3V/vfZ1upe5VlNQFOyneyXgMC6j8CNOVerYpMBjZIpUmnqxJO5HXasa9O0Laz
BB80NF6fR3g3TjfU7SakxIu2bNpev0nY5P46bEEjWPGmQXWvDlZzwkA6gyE1NQ2tJ0/ei0jJQHop
NrRVVeD+KhkgOYOGfZko8Mj7RwktaOTvtZZy5gllVEiJoQlZNSfA3So49g1EcIhOdeDXesQ8CFQ9
1vuHa5VCk4B0wkA8iOGJTi+sVDr7xpmnUhEM66vpUe+BORtM/twEn0FCrkpOP0VPSTKlljJJ0t0b
guPIup0bWKyES2MArhxCCo+Z+qEwUKV766wv+I9YaqoISTEzByEpNV/9hsVk9F17wTeMDLyPzQ5L
ncmbM4W5VfDFfeSHqVMdaNPVNAuP/ScRsOaY2OjJS6DBqQTPWt/RGMsVPHiSGuzAytU39T+hUJNb
f9wpI1nDFe/LZTGLakNHXu2Q9kb1mVG7UkN+kfKlpotbbZ48T0jd9WAAXWwXUtIikJXcbTU3gqTl
mpQhkjxth4P4A9RdBw0mlRBO2e/aF2eBfvZvlIlQ6/CtRxXkkfEFgOPaz85R4iDOkmfvD6CmuQZg
Xs5I6dj+yO8mLDBtY0oZ0iZIKinZsCMToQjQpD22RqJxlHBg78Qu709gtyAY7abKHcRAb+vi1sPu
+qsWGdYU/pP+PzsHPkgORnxXCYbx/1c6+2EGx2XQ5dHQZBvzhvn8S57kkheFPVIDXF8nqC4ZjEMl
gXOszFsJrI+5oiUVuDNS0x5+/zlcKL4MRqcmjK/GW3LZ4ecZ8BqMG5XzOS+hzPKRorUwg0p50asY
2XaG7Ti/9SSF3/E2o/jGIWdHSkgfDxxmS+evRaHGuY8rdaPkQUFDYr/k71lj3IcbcDV9+I0raRu0
dLtNgfbSH4v6u+75l07GlHEdMMUkqLXFzn0rEwWYqToy5WoExz8X0JYRBII0/XJV0yDIuKAduHe8
ePo17I8LI9YlqwwOM1wWm6lNf7LwW0pz03CrTATXBHvVXZMQZw9KMGMoz67AMIpQIf6mKGhCqFGD
gJyahwy9NbK9hoRI3dtFmthQXd5li/zLwmnl+gfADgiDyHWfzE+ZgMvYN08r88sbnawpLNWGHuD8
2fhGxuHJzm06svnJLSVDpLrCMVyLE8hAdofkcGihwlZsWyI1rvTkt5HdKs/iDaVJbrZ53pZVqmgq
Yvvhuz7rLQ4rpDIXPJnyPkDlxLxrEKEGAuHL/DCU1LV5ZkHITU2N3GYChZSkh8bbOvqV+GLsfT3x
/DCS22REmDfojVssn72M7kL/Ag0xSNo105FsW+szOJAV2jtVMwRbXfCH9/OpKr1exzIFCxWWTrWq
+NIytiXv/ThqYe5rgnJw0weNq9cmFUfU+9+c8zy8Z9oO4RPzgBhisxiO3q/jdg4agzg6mEKnieTT
NoXZIiyRVpdG8NG4Nlz8rW2OuiGr189keKyWDDYgTQj4xwZ+6f9rvRva8e5CMMqWw7qqxSc/c4Pe
KNExJd7E37oU12W+eUui0nCG3gneuvoPKWqYouixR06L72SKHiLLvZme6UEfup8Rzclm+7MWOQoB
5PzrgyRt/LGhi1RRBIKBt2OTKbVdpT38bvBEdfiyiv5VLMgqW6BEOGzp12xzJcmvjKPUL4fYSLe6
BbfCuVmQQiNI2Zt5JJ09US7G9QY7GC2fBfBz8SiMgXQLXPmQ2i09jf/xWA8Byv8HIC5j+3SBsED/
t2b5eCpEe+zu+muXwnqtlNU94ofEsu1HB9kF9iNYOtyUyAI3aOiOWN/DS25ntOIcmL3BJrm/Mftv
8o8H+/vezAZSibNowk6SyHfc238Ka59QbgAvHtMPYx1csy9rkP+vgp4C65SMDy7vlAElwhnhFgph
W/69NBB60TaBieIOfTDQIOBwwVgDocckQjlFzMkwWZIXfY3auqhFn2kKgHfLwXUjqiNpQsOlZLre
mZHsmY37+YTqo3nPQqjWQw1GFuFwy+600xdCJ6C3ZwjoMIjeN+58MJv+ddc6kK7NARxwLHIiDuL9
SQvRHo9Ie1V2XRB2mslSYrDDhzhIkJ76Fa0PriorUTL6WxN1vxlzkOKe0e3l0a3CqWNmv5rpNB8q
Iri21kyGpDLhtM5WdFigbzG12KmdUYPwZ3kvqjXGcaAIFHMK3YDEWhel2T+X54PZhUsF5Ml/xt0e
g8Ffv1N+k0fC4AmAjzizx99AJv1ZUxc3ZDz5hD5rqNYrT8vd581hio9zQfLCRGETl/3fweubNdMB
++tq3vpuRlolNpDYHRH10itcPlL2Te0VuDIXX1UsKqkS/CjPIUrlsQgyYrEdWVy+VtgE/wkSN5xP
NGBsJrd8FYbxuy9nfIp136rCgOFPER6Ib3ucwcjTS5h/DE1wMRko0oJyXOTsS+c6cdqGtMa8ow77
JKz+dGl4kJVr5ZV3xyVaYOuAaXRKAlCOI1vj7LUqQnTmK0+y/XB/xWrqW7JbrWE10y+/DB+Zy7HE
8vm6Hrg9cX1RNp/RdqrDrIlkT+f7YrZf9J5NvO3zTD9PC799H0WfxsylFNjzQ5ic4HzmO86MZo9n
2CWmvVQTtd0003t+2r3TeTMXyB414qnDnzt5gAi4B3sNG8wcbI4rEfSzzay0OZklxt0h0V1ZItEC
bkO1rZFWD2ETMGUVk+34PawXcNfeSE4Uink4JgdT78Knfto4bd2JlPWGao5VcRrKbJcUAwm07AIE
sYGW+76U81s2rNoG6TuafV3Ng/YLj8LQICYTQCCjsjR3q3uACHDKzaTqecCPgN0yQDcDk7+7htpw
IGomDJee2Uo0ZA2cvMuChoKAmog7BDM41U2R8rv91GRLr0BuYgy3X8gIzAZhqTXWWaPgNtWT2RBF
DgceANsZpaav1n0XTkI8zX91QRqumBTKzWpscrW5rYwXMNXFJpabaJkagbOXUI74ajnrCN8InTRG
U5HlYeZuGBn/YS4LEKlHqhgZjyVdf6MyELH+HHB3D+PQLNmpv2WSl1ZX8Jw9lJ2+O9j02UqGp6LF
iavbV0825eQLEKAfKJppH45WSUC8K3/QJFxh6cKJe8gNFKE/f47u95A+KUtkNWRV/e5jJFUoL+nD
19XxXYNkWH2SsokxM1FBPwUm2Y6kIK8wwjozWkzH1wXGjzudvj6nuDNe7oc6YDf7GD+BbCTuhSxH
47LgWIvnapqfNtIgBYnuPWO6YSY6a5YpczuwCyuCM+bskf6H2GOX6mxM9+k5i25WV9Wt6e8Hl0cw
KHb/2TfqQfSHbjKtfGU+QwWrZ554S5lrQwLd1pYgyS6B+avBAG33X58lKENtnvhdbWN2vhOrbfW6
H1F0/+iSULpY83k3OB38UiM94Ylj+YDOBWK0j/LkuqGcMl2AUGEUtdiuGOciGn8FyfwgXbKmUMMP
9E921CdeJnDSdVh5Nj2jOQhB1QaAhXWblpR8/h97lc+Xfm1zrmyUhK4BUm4trhhCC1sw8v8svaJL
BhbGwoPj/hgJNiXFoHOmGCawde0ME09Qp3LkM5SjgQGdNQcAy2tlAwpXZpE1oxLr3x9/VnPO+VjF
BN2YfXPkmLROMvfey2hrmAzDu+aGRYeaQ+gV5TiVISq3QCNEMnHg+TJFhXsDkMdYVD5xqW6pzvx8
p1bQvmR3N272q2k2Pb0rhQDNBcbADHmzqtetfYrbv+gQvT1WRFuPNnS505euYkT3mTNMy0DynB9Q
s6gsnnRRI56rrCP5j3eaCCorIgKkwQObfQoluI+fcAkTW5m9hik+utWAn7JDsiKBsYT1UF6+XW00
GQlqjMpw7Fl6tY0oTm4wPMxX8kz61HKk2fJbBtWijuDJA7ncxZsKXU5kzENRjOx1IozDzMoT1yQk
FEnF2IOdOoo/DVUiUlfrHiOyUaQ1kEjyrKr5jQiVaFG6Q10AJRIiX5qzxjcCc6Q1+MEGFQxDnL54
veVtUOlwRb2SdErwBNJP505XD1CRZTGPpI+9ohFy5HBaBbjlxxkkllzwnOv9oogaug0ehg9UETi/
7evu2TBd8rpicEfiX9lWderkFufhKIFhO0m1QqkSzxG+nPNUaXO8n9Cm7WbSQlc7Ix2Cc8vHKH/s
BM7URiFsrxh/WRfK8qy9/gZRozaZ0D870z8arfaWvxOpNOc3lxyl9tNF6nUeVnM28Fdivf6gb1ro
nyfDeIYxCPd4bQ0cBnCTP5Rs05yJPKfic7ITZR1EgfaRe0Dn2eFqv5JbCKPMIMx2kdtIgfcaeTsJ
8MRlghGEMf0TiEUSa0IqwT0mU8tHY9cgqFDXG3+sV69Ci2ieN3rTt/hBpyl5ToJ7fZD99+JpSlxP
tvNe9AVehIl9Athvqp2NN8K9PwDO4Xzaavs2daMhvwVyp0zYGqoeXI+lzk3UFN9cZrB56ZWNhZKk
MPzaEC3rcxRg7GRQnJlbJcbidOhg0JIVENK/JZm0avY91GUTaaF4BaVkATJ3CIzuCLcevfBA7DDQ
ORmfkgpZtzM6oJVoabCpESgW0nR0Ze5UqXwseDp/2o1Yhh5rL81GvQxl+uNPLm0MdATluVVBaSUl
eRMZuzabWywSxKLPat5RuG0AmtgKgF0J10nt6ubWmr90Ujx6s5Wbf1TdiSaB1xTbTFPJdeJ7MMUr
mKmcj567G9wXfQCm5DAOmVzMmRufQpyAA8mRH5gle7thpep4irNHtg8PXLEFZgDl9HWxdvzhOIRy
oN5l72iSly0blc+DJuIaC3k9/pC+vh9DQ1sy8KPljW2S3ozelIm7AErRCRLFGhErv3Fcl7Zyw5RE
SyK2xy2gUNm6PdZ7Vum/mH3J4ALMFV1GpP6lJnTYg6NZ82MD3dzaENEMOQAsd6nYV0jx8KSoXArd
pHUvbVhAIXuMQNcEuGkiLooj0MjMowSF3PBAGssfrOC8us5BMpEhRTRaC8FRhh/oyPaQtQLwc8nC
jum76JdEheQ3MBP4EReS/rtMxQmpkBwXX9wALZIQkCbt/antH4AS9ckLnzUc5wpj6WXQiTJpxRuN
vPh33edWsMLnX8w2AG7nz7vLVFKDr95vIryJYtfXZyQFMYqME1suHtsZiR90pOUapfcvURthVTNx
cubswNgTtf+8DpUiM/wksJYv39oPoS/rMm92k6PF7U574zgMboDpLbLvK//GUYmoURCbVNaoLmf4
A6TdNaMIBlCZGnF+L/uHnhf1iq+sPmUHs6zeaElUJXjc2gJU97KBtI5BoMkojtMzQ3zqLnvdHTll
2522hr4A1v05O3/Iu32NB8Mlx5pA/iQ1QKvK/hbke2EYe/bIIDG8MhVnM33cU0oZpcO0eoE9m7V/
Zj0YuGkj49Rz0OtilT89Kk5rn7nrO6brbLoDkXrhHdYFcotVGQ0mIsvuZbcvgNiVDNI5Ku6gY/wP
tQC2kiCsytx3z01WWevRiVWBl93hlWEfewcG1MYRGSUFi6GgTP9EVdaGF6ug24PCgslQz3zH1Mz3
r6CdlGLZ452xAVachQ5Gbhj0UhjPm+uRRGVM66zSE2Xb3T1GSG1SGX4OOqlgW7Jf1DIH3IAICp1f
FbIywD3UQgVqnyNlU9uJgRnQjR0Vr7smlE1qVTUUP2YXn25ZU2KaN2lLYipMO9KLowIKRakjRBgc
6XKQM8jsB15xvgcYJyn2X7RpEPfPPFsW1xIXCbGiQSDv1B9P/ZUWxZxw5SJe23N6OdhXRrEG91j4
/S3nUQASAsZADrYY7Sx3ehGb/FAHFmIu6wolyKTEnTrjtCUBexPNTJrRn+9CHpgAsZRrlYPYTuM0
F5wDZpqHiRdpjnbqxMqA+emzXVLd3eOdX0U2A6fANJpPvQQSxyluPqnMwZHOYInPFEc9D6tJuYEs
mA1mJ5lE1jlY3XLReHt5RzBuc5nBJYPn2TCcgI68a4782zkxL2hQSKXzj5CvA+vLq4ZbXhd8Y3Tg
qtKuMW0prQwRVqUFmvM2csExOtHOMbhl0WjeEt7iX2icntdDOEsmq03oVl05vJ/1RslqcaryG/NG
XxJCyw8mWOx+O2Sx7h7QtCeu/xQY6lIA/oiuxv4N/4y9y4wzbBN9lxC0wfk+azOdd8eJpSgvOEc6
BZ2Z6wVoVHilYhcSYY7A4LFX15MuakKJs8ySUcrhV0NOAaXZETlKC70PblsSMq0J/NkBpGkf+3cc
6Uu1QpPDyRT7oFpdrDsTudYyjPNoT+4BIb6rMPkBGRp1RBB0HmVoF6cnL+fV2kqnHBxHNYPpXBZ0
GvYyN7QF6RRIoW/KBJF1PU/S0geNFoXwcXz/wCngJBy9CHhXzHCjaMaUuyg4oubOMaiXJPW88FX2
oqOu8l7KQGFSH85oS3jDNRaweloYteRHrx8z72pBnIw4qEd6nkcqZ186hKkG08zHkG6nJc/VjmYG
iqkcq3PhDq4qaizQpQ+9EjA7D0YD90d6KjyjRaa7bEKd56BAhFRGqRawqie218AQurH1SNpL8byP
exfhQut07nwfbnOLMASkF8e04mqjpERUtM3l7XI1b+H46BC95u6FHDdvE8lbXWtE8v6YiYQKTPom
henup8xvGtp5wUqhvXY5vtAy+c6Lh4QninPSCd/tQ3P4G5PU/6PXwUy272fo3Wk01j7g8tSZy5m+
OhGMuip7vftnhrXz5rKh8xibBQ1jZztXE6+hUzbqK56wpv5Kh/en2eXFfTTpGNjIj1Qw+KExSVLU
PLiHOBZApRpcwBjrCT7BYftxL78aiE9SqP0uriPqoMzVtpHsUz6RppMc3U0bkZ5c5yerW8n0gD6m
qSPdt89kN1Cd8RWIBAC9DtixJ35DmarMyATJzV5pXBOHpNfSKycIF9bhbnGItyyAnKamQFbtQdNh
YsDdCiOs6MLppg2a1OSVoUPuqiLzo0InKnc0+4Kju4rSnM6M4IsrgBCNgu2yn/iZRL8s3aQHLPk+
OYUFWKQwSEwM90Dmn4fhoOj0NypWTfjJkASFr9kJr+VkVka/zRAhGtYCQIS5u8oaYrO90z+DaHzt
E4vJhYKEPKvk3PcTJA4A/eARPfeVgpvT29CNkvldSR2F3805h2zd/9YGigZTkt3IcYx+DD0Lv8L6
KjoMhZly7GuTnaWVnIH4/PlND+0Bz+0KAI4uC/ze7aH8svGTVVPP30gk903YJb3mBdIbx2GfxkEC
at27rd8sPmQxFde5n8gAdExueEWm29K4LLhvIG59uJ4ELr30uyJM/JuMmroAp2LZTOJE1WqNCL4X
sUwqn0dwUB+GeI209KZkzwIpbUS/6GUUbdcIn133WcImLhyp5zpQqzwk35k/Kdtxsr4G+f4NSNv2
6CHDlPocA85Mlwt5LV0rzgJX5YHTA1E+ZWHfZ5yR5WnEZpDjcJLQFfjJzLYYpexHrQ8MH199hvHD
mgAbs9tZMZ3NVjnP/JNIcCcMA72kjD1N46z7fgLEscOor4cQp33RSWvMdh9H/9FegafHqIGQjHoh
YPrJbAEJDnLKgO5tydQv2NHxwhoFzuz1oBuFDrAFY6WdBEI2/l6we/7tZyL2ZuP+nAXtcxrtwzS7
6DKoDSgD89IpOHhwiF5F7KCPagtEHjskhOBXCkDpZ4Z04lgWAHnC6tLVh5Qh+WuLI64JkVJFZNvO
5qzuPdhX2SHYomokpqn8et+zcIG4Xyjdm4GSJs4G3gaoKugDc2sZQTdc4/UQ/Mvqc4xqkLCajB2y
lBSeFBLb83yPsklYoFSV2BoEvySy7rcOh5WxXhaG9oVOfdpBI/XxJH73yqipSGk9bTW3o+kIslxV
32BK8n9QO4GUdvIMLh0fyU51QocNNnqjUoyfrdSHRi0qoS6uYy2bPhcvMw35KTksEnESycFnre+z
tLNoUrBBabc17mfmMD5BDDYLyhXVt2eAUnDCqKU9e2XWhCQJk1L0jfEKiH9vtiOjg44iWxUPfhMi
a77bizGKoRlyjvqi7L9tzI/PiGmZvATZ7XhTc68PFmqohZEk4g0bl0seniDdRE8wkJzpVlXxcWd3
Yaxo59upmspQFNVOqXWFbssKobGn2xkBMGpGniI5XCKEE7gPciYa+T2mw84fWtmglydpCSTtdItg
pb15TH8yA1JwVRNGgCQUXvDy9/OJ3bBEDXy/wkHZfPHi4RTgojcvslgD2EAYQ2a9twlLMeEUmA3V
FypXCYi/9rZrcuSDs8tqOcFsIv4DW01wwJL5xt0z1nb8d0cVOXJvzCbnDRXQz/Tmo71BNPlMGXJ1
z6lYe3PuN0AB3gAwGX/KKaHq2eOLG5kqcDAXcdAVb4Jq42sJbGBVsgmTRoI5TKerBz71vb03GWdp
1jcoO/HmuxMTEhRMidC2jg6TZ3hOY9JkzQgxyGRVZ1jSrWJFIss7r0Ti1QUeX2h5CKFuT/7yndEi
Q8ZJBVZCtl6bjQe/3lO6rhMZEPPiUa/8tWzm5VvH9EPtTvAKgIwWQdmQmCWsdQC4AkmHzMmm/FwT
38Y/+DFdTCp09wCVnn9T8tRFqOZceU0yz+qOsMFN/kVsSaUyuIiDWFpU49T4ME+QOmMhbKzjwGbJ
9WqPSBHi0xh3Z8v7JCaULYMkcA2+bFPJ/PPfDqFDl8NlSLBeD/viYNqDX3cfSBuAVT7ikFVJ7kI7
oJ1dyXlzX8QMwuyeN7i+0g4UOIHsSQjM2c46UPhDnsQYFd+7Kx8EvMZMiFU2LvZzwygGyU2zym7i
GLm6rGNEKIuWqORo5/ua7P2SaUlIMfALpGd21nMZGvb6o2rFibUMXLHLrtkVWA1yL5vTGRoKqDTx
OKDh0HvI1pS3Xt1ptc3/F3mbBEtfmJOzwJqCOpbCXkn5NPqMWtPKbJoazoEYYVgb+Z7hoOM2+KgL
jLHFpYhgQzctGRziCHusHXmdAj5309HfXJfmWn7gNg3EXxPPfKSOl/2syYFlCvapi84czvi7C/uv
8Hi3jv0oXVtMdCKYQ1X2sWLO8v8fgo9PjP4iJoRkHxGKGd7R+Oyu9Yn6ISDX1OXMUci7/ANHUyGt
8ZJDLmiuJRODHeSUQyYtwpuHTqnWs3NirJCFXPGL2JEr0ZkVfAmJwrx4tPljMXSkmSC37KYWYPy5
bms0K7at97KAg2CFamFSFlTYL/XPmBQ1YttXovVvDBJ5pfyOavtQaLSnl/1y9olW/VDLuH/KUW3T
Ev2Fsm1W0t5qivyErmFYLgGgUss7WsfCPS1l4S6eHrkBENt0t7FZWmexh3232Iz5LlIEP8kyze0S
7Tds9hhwlwDJ8U0MlQCeZDw1GtfB1CpDG8R8TQCCDw84jbUmbP6OPei+OnJTsy73l1pTTLk1RAzf
ZsSRpDL9+GPsIlFQyzUYGJwEl/LO+kRe5Cd7Q63Y/OxUKeZESOGViIYot7yGAUchgD16sVhiAD/T
57PvwZvVYSQGWOG4It+yrYqkTpqXZPto84eaGZk+uHnYplDPf22y4MjEUBXOdVtnM2s00l5QZ8XX
z/Rt/VRLW9xavJDvP2YrdiTwTeRA976qs3v08DnU4iOcyzlLs3KBWn+6qLkbgAtBTYPpf7ai6SJT
L/o8w8OXn+xHeJY+G2Hxo5dlUgalL3oijj9dKlnaB9tzx9VYNEghwiuZVjHGJCIBlqzdK0BPBv5Z
pbnZpTAJU98CVKM/ucRDF2TYYEU0xx5MH27YhEIyVVDEZsmnxQ/n1YSt8t0EB7HFOUwseLcBn24x
YwAURdSGA9KsaenaYBUlHmfDEQxsDk4cuZ1gP/IWP/H/sWKKHnTXrFXKUbSw7cCJivV1fndS63rQ
7Gn33usvtwMZnXAbruE9j7qH9LlHaQHYQES0fFzJEs9jSHsAfV2uAhrsP6I/oh2bNqpsGAIixMWL
Fk9yAJSLu5j6ltHq3H5dqTBc5wWmNjqByPq38e5SEtYDQSiXXpF/dTz1hYMp7Pw50Aqs2V4SZQ4k
3YOGBBkF+ADLnzs86udbx4u8tAvMYGh7uirLwQCHCylAechO/l+7XBT7vtWLHLue2OhxsxtOKbT2
gNbvYWYfEWqs8E1fM/paL8SExSK1ZPmbk/anY65Gmf5xy9k/GE4AvwqWVUBwaSiSNeCZlt79cX7v
a32Vdujdw2/dGLWYR76nfynBmkoD6qmv1HagOnfXaNbckEw+M2sbsH1PHUFZ/H7KVRgO987e7qjD
b85mJy2aUjZGULXzKeC88vZBHkCAkXmI9Xn/MT8KWyA/9lRFYgtJaQqP870YYSyy5dQ/4szSf8r8
2RwCypqixVw+obe+lJ/7SZCKPKEIFd/VCEYOtBf1B7KcNcI8MEpx58ueKO85R2o4r8PJJnnD5wy4
nbeev8WMtKZiN86b1t1dSW0u9aRrPpnLCItBHnvWjQ6a+hFSfV3SOmil+d/uJII+2AC3qgLrO641
0i/RtBgqGEbI+JHCHsRfIK/QKeOoDTv0qU2yDbTbi37xBU2qcZc3+/RD441Mk5YmmWfg8RpfL8ie
W7SiSnXTucoJIC9hcoVMjtFV7XV2Ryk83IKRHfcYQEHi3bZcwpnrWHO53nfaKUpvMr2zp2BvEepv
lVeHdynRn3r4kACreMBSS1xdE7GE8r5y6l2nde47rmh7c0WWxxfblNDXJ6lFOPvPnQDk8gekg0cJ
HP4zY2A8sFmac1mgSv/mrZPS41ew9rpLDeH4iFgYSqzsRFOuYQg5WB3k5+k8oIUAoZGkKxYPhwyJ
RTUDbS1Q+e04/5qLzVKJeqJ87+y4CY/V9Zvv3b5tX0yJh8sbknBA27nykdXVUyzrA9ikIjj5Y1LU
yAW588CS7LWOU2bMreizbgVQapGOKg8pJzBSd/+KbImdvfaC3qs+8SAE7zvxuNcmhVSAEKY15dpr
n9Dr3Xp5sDS4kswiNX0/jJvj263bbxxmZbqogp34SezWeAGaB/8twyo7s0V0ydGg/7svU+foifVs
xBcQPorIZuW6W2aJufBvNwzfw25TqQIc03QtaNLEBKcND2alfVWKxui2oaLpBsDMlYV6b91t2oiq
b05ktl/oE+EYzVoORyY70etk2Y/rsvj6o0QQGovZyRQ3J+wDPiACUcKSQM5LFv+aGM6IASZoAgQD
2lGtd2XKs+PluucoS+wO9mCwdVBzO4Vf11AzD3avycmg3FB1KdUqUH+qL7m6rqrqTVYMLTGxpd0L
eZZ1cR8dHqX6oHLnjKH7RwcZpbxULtv+rhxLGhmERHQ5R094HO88B+b+UlaSh3PFBCMKmV/qtKgN
6ukj8c3jlyoTSiY5wUxrkMQwnFHSd0Q2IfLMKhhjTvuAMlTAcq/D2R8cngg5chux4WDuJMWMbOTU
qa1tQ64bsHK0F2VaAIdDjqWWDhjTA4XSxlA3/uUnfYVyJhRUT7bKFLFVB7N11YI9ed3WrLy+NZXX
550T5+Z74fX1wf9vgQErIcOaMgc7Dv30UeCAGhdHqNSWZfX7APQ2LI68hDnm1gGYHfugGokCxqoJ
IOjFYktc6MdpcrW2+ArfKbeFQIaoPUITpANO9OJDyT9KtkIWYQ2UTDUx/zGVYcARfIv73w+ayBIq
vJte5artkaiIZbOavI40hbEgP7Zagp3nTiHRvI61dw9mmzC4kPT+YhOkgFUH+aIR/b3/4uyXRVf5
xq/hCA/dWdJ12BYWa3bG4JNu1Kc208IR6ZpaQ4CsKHECfxMb4bzddL52nW7U6vdW00a0LgFhmsvs
SGVs8KyU/XUNA19ppjExI7mlrIv5aBPG0xZIHxshnVQ2br6JN6TaYx3BQeYrZPIiRsUXQqoLs3a/
FrSacexYG7Es4uEqVQqTRkTQaaY/WugSADIVyWuxpyP9GbP9gjxrDQdya6wAEtIV1FzWPH2LR7pH
ILOWR5Yy18TpPGya35CAceFDrx1PlGbHXJ//Wrk5emW4lW7DGfyaBMYHOIIHvwjdvPvG9yZWIxSk
/lSX8Eex/YV/C0ymJCGQkQStbsYiIg8++0W7XyMES2zboM2XrafabkDJRwXtSxWJMM6xtoIpN8h1
/KfsLb8Ve1a1wsFgF0NI5RJoNDRVPWv9G7sPow7rlkWmqkcPUXvmEcZpGzBm3BVuUDuJJX0wlL/G
Yb2emnUWiJhvwoFU7BgtXaTIFeAy1lq5tLnl/JbqEmyg6bPZjFzEvnJ8vbPZbIrRUh7pbY3ISDq8
TnWRKb/LElp/DDwWPj8oliIXHCP/nRNQuBiVll9XgbW5AxHrUBsT1d3akt+WoG4D9Laz8TOQ0LyO
Y5jw858HCWqmB4m5S73Czb75ht3Mv+RHCyeFexLdDA5QAawYseAv2jqpUi9vPOVY8dlpkF+eav6M
0KuK/iqzptfP+wdLpkaiLl4dXcD+QG90WMS8VNzw2yzQLyDsdaOfLdBRl4mvNsGrkKJMYhNmh7Ds
VmYopfHAvvfPqEO3CW7nxwDPCZz9uCTOON09HJnZE/ch9QPfwjN7ZJCUdu/si6yhrmK7y08ydLef
ABuugDSBitYUDwxLBb+Qh+Eap8/qCzYTWbDKSyjvHJLUED02relLOvcR3J3Jhe5A9y8jFHESEYR3
MqG6/mSFA89AVgm+70JEtDuJ0//wYb0iQ6bVrc4tEfCITR7hMr8mVFV506IPGP30v0TP8QWkMb9y
y7iDYL/Uc2j4/iWGZUCDumya9cbIpmzkji4bAmn0n7HHblEE+N4YycUvbVvUjIsZlmmLIfjXC+Zv
DJsPRB1sB5mUnwAyxvqkZSOXY6JLDe1yYRvP3y3baxEzoEc/V1Ef9oQkTBx4RMTENao6UG4Wk9ND
9PPnTZgmx3SN0VuAAMgJpT6SrIMjZzrftNOLJ0HmdeXNz+2hep/H8em12FT/Lx+x0Z5nwd745UJt
81yWoLB3N2Tea5TmLXj+YQ3h6wVibBD15j4bEm539SdYo7UUq/aL4LX9tqRxDr/msYvq9gtj3IAu
Le0a+fRrsO7XYPZvMhSelAs9DNy+wgK9l3gvvH+uXGXDdu9N5dZT8J4L/PbyqPbmleR75zrBYDN+
Dxy3J3n08t9YhpW7Kj/qtgH1OGO2ooL0lc3uFiB5HZh75mPzOrNWM52pnD1jQ8VPUlG6pZJ7/aGf
kV2TiTr0thBBoPqFQ8IRJDDqZ+Ld8n0HR5o+LeMsa9Zt6+mtg5c8P7eTM4ySC/viLzya3H2cyFrN
CC1Vs33/l6fCIGEhIa9s2AA/pmV9azKb/agSv5XwZ9qaEICgnZjgQcGNokwj4COLZS3xDDr4OLjh
wkbbSZemp/RUqclxGfzrXr/qdlRE8ddDVJKxnRFbSo7MEPqiPlEApECtjkXdOph3UAIwoNa4T/B0
V+Sj7rZMAjrrt+d46VrSWb2/RkDNXfyoP75cSvF37aD2DLCMYc7pOAgey9l8Bgl/V4Fdfqsnf1SN
1Pyt60Qoy37XZa+AG4Ij3QlazLXFf6VHF0bPoG2qYxyP3zNANR0opdqAqCFNFqg0Yizqln1hf93k
K1pub6Kuq2JOYQ+3euOQrznhtDMljSxo+v5hJiX5yfV0Rt4FPWciiKdYzZd0IG5DUq9B0DLJXt2C
cUJf++6KmvTMCdQLZq23PJ0UhDKK8P69PGumta8YRwwHZ7cathsDjDIhXse1BAbfLhJGjupI81Nz
l6PJ9dJUjZjEhfdCoqnVmA/hJM+mwUz5EAuYA/Bd18d+ZX8vaudPQ3F3ireDO8ZdZzzvRmB4NLH0
VGt09QRpX4S3jgQLAAGelBbILhq17sGFFGhbaAu3Mrb2GQZLHu2JeewmpOm1Vf+yIho+8s4u2Et7
9ajO0ccO/mxmkhjnzcd5FTp7COa0xedSQBeIJG6Y1RQtslsPzdig0lZ12UcDvNdI+kdDZ7gNEoQg
dqyAYHiQ3D0T0hOcPO6COc3nWRRoz1yPrU1V/h5/0oeG0T0Swh06xuAPDysbvqRAtDkYIH69zxRa
gSouL61NmQ/t2LJp/OObVvjjWE9X1DL6h9yZm1cfjFhwOf5VGcP0sRXh2GvIYpZd//T9h8emPbLG
w4dtsTKH3HwQImAsKNg63yIvo7cEViHLL54XvghKPLUIsyhx4xWT2Lg3iABp8Oeif5bmxIl4pm6I
yjPOuldllLa3SBdj+LV/skxaeYvAS3/Xu2yEtQE2UKFWQ7SLi+exaRmTKPhv0RcISzCFVXFGFw0v
wtX29Sbo6WqOheN+VdaLcE2vqrQcUIqImIxdCr0xwOAxJr+LBk97qIbhFzQkGDN+9Ar7vab44lyw
QikyVmBXXOMr8B8rMIzdPEKYBvg9D79fSp6y/r4KQsEnhWk+UrF0S+74eeN7lcQlXtBgTYDRSBfX
ESNCQjaIlOHnszUINKKEwH/gj+dorem+DlFLl/iqLHvF8hf/dmM2IM3KGUapWbhIKT72rQGMFy4Q
e1qD1f/N3aXi2kfjdGD1Ny6kxPFNVdkKwZM2koXWyfalemlXAzehcFqUlviz7m/MuvE33wtp1v9Q
D1s32j7oodNMTR2Gc1n0JiLQCDXliEwmMrIwxS4vMMtQt4ygZmtJ2IJOV0r/IqkBbA6GMQA8zeLc
7tJEidbpKmDchlL5CEg2Zx1yuiZEoWj9WGktgFvT/A9LLS4BfaejGUqA5PhII2M6NrHd1EQyVZKU
BQK/cLyqWtrvvt+pbkmOgm2leyx+1vkC/t7cjGBztC2IsQYoC1q7F9fmHbqC7fUgeT1CuahpyZDc
9xnP2i4QjX84a5lX/jefHcAVX6GG8L2V2rL8RTnqxAPSIVXylJNzRhEz7bHXPxYUx2oZaMsh4Bgy
KzBh/MMHiRyJf/L3gfO+dc4jwoITjzEcGZ0iBrmOR7SY51SY7UyY9gNThY9dbDFYsQVawt3S/chO
Ge5WEpsVAV/PGVGJmuCKxazfeiKuj6CMJut6p4BnBphNXRwPAidDBqMj3q1iiVG4Nx0W0MDkq2c1
cJ/EEU3x24p77KqXhwWzoJt7qhzZ6LUU568X7ZQrceFKzgrYu+f3q12OKZsLukgEeBiFafX97GVu
EUEvs5W1srUz1XpxQdb5v9QyrGbF4Xm2fPgvssYHQLLBDOzHvubENgwZ6zq1dmdVPo/hfMwLHofb
YvO+GYyjcVZHiciBDk5t1V21gYepqcmgsL9oyF3X40oYw70zPvEqH38reJuqCHXBjhvXKteKkF1y
hFFf2v7QwxHJfMM4bS32fA/nYNROZtYipt+Au5PwT3fawI9LOrIaHAaVVfw0PquHfEYWRQUIeNvL
TRBXH+oIWQhUGfWz2TRo+06gV1n+GpXHQ1ZfuuUQvrI4QMatsq6kWxSkVPP/cBU95WwHaKHi++vW
rK9D3g1bRahh5fF3s43xhi72Po6ujN/A+cp8GllvSheRxx1eEK2OOY3AaOrHfoYmxqdxX9s5Zu3x
HqwCAAlEfkHDXKOOXBPTJFVDtfYSDTTAd0p8hnIhyLewYxcOzki9i+UZZJgvksUae4l7sdUI+LKL
ptcpYMvrzr6bqRKLiiTfOAzv33Hi4ueu7iarlREKG9hiQ1uDMoQP9ZfT1yHC0meLNjp1ZkGzzWKQ
8QBwStS94X6wdNk1bTKt3XDr0nEOYr+042YYi7fBQ7Oe7S06DjLwcgPAyGNXqDOoPVEoBhnyo4K1
tIufcEYWRtq3r9SMUz0q12KzC4GWyF72vJl923EYxaFjm3IHKDdfyQo9q32wO6OVRFv31LDV4i6v
rn8YfV63EMERZ8Vt6mE+P1LXso43hxjZJk588rc6Uex0MvANxNl9pxqueC6inS2IZ42/TSAtsNAt
vnLinm58f1t11wOirxhW3i1wTlE/DRiPgVC+CWHqFBW+Vo6vBcSFGljBuCtX/DV5urrkScb2vYz5
rx4GsU5ctBC3Dzv9Gh/OxB/m6iWfSDZoFLosjw4ws2TQkTc6dbMc+SRo5r5Rg1V7tktQFsQwUi/g
07ScSkUqJAje5SZpCpy6BS9Cl0qL5UT/PodL9yIOG2gAyImYKRrCjS1OJhV0qZtgjY42J6+GwlP5
f1NKkmzJAwnScJg/r+tnZv+qNCSMvTLIvr3704l5KeK5g3OCS34j2eNZJnzzjh5hTn/s1cyoPMwg
ly33LZTf7MjNZMV9/zz9M+fPqf0FRPA3FOV2v6g1IyD+UQ7HmHRi6aWTVbIHFeavgIE1ri/0G5ad
M3Vvrj2BmOyEdC3jDo3RivfKwMQM9DeD/VzrtuZK/9PyoN9h3+5kMySDiiMFZ7pxKVppPqPvrlk1
WtNk76CbBlJ0vTKbqIncudcWTMvW5kyl+jTuS72qzSai1fUwepLb9OIzAQGRNwEKTiztMe5me/cw
f0A/vP1WmJVr5z7u1oJfr9/Q4NrLp2iE3yjJFI7hmjzEniApd0ST9GVlCNXTj58wlsu0Mplz/jKr
EPZ6AwUniGlgbeFamceHu1TPwkTx1DlYJ6FPbctuDyw2ssVaH5Ps+imv2/eVrWplPDTUtIQp2spT
ksq+nR5n8vkb/0FrsRYPCz+fMAu/TEgaWyZJo2n76DZM3zjNql5uXaK92ds28NHLGySCTIYA72lp
76+cQC6yMnbJoWRdl/XlxGSChM7yM2pZ4aVih1fQ3fwI6KUyA9ERfcQg3FtYajRs7XlsvL4F9ZVN
3O1FuU9Xiqeabair8NROAWZNLgxb7U9lSsmPsx6C+G95K5KD2Tgji782q/HOTsr08SeXHxI3H1q0
i/czkYKlqidIaEVsQigca1nFzvAwFNDM8ApO7ckJLeHG7Ozt2y1Qs0UsMVcEkWF7BFqJZS1nvfd3
sZo5YpRGdDB0p5tCGBoE47b8BzvZEpFEpxwkIj6TtI5g6orvk6M+EPZsOCL/YWMiR6KnefIs1Dfq
v6w4qCsqEcXRVdoJWpgHIWRnwHY9mYPvh8aa95BgwirZIFSMi9hHahjm+XXxt7jRbsT6YA2jFafc
gtt/wSF9ZSchJ0CdNG55uJBGMbhr9dnkd3eQk889HcsPAxyMe/mWFCxgyrVQJ2D/Wm6/ds23MRtB
7bB6E4EThHp//RuktuzWxzYVPLUNOUMcLIJTUYtgdYA6HGKw/kZ5RBlN3KssW53Uq5SJwN2k6e7W
dA/txr6+3owN5ytKQRAAmw5WShSmV7YdTmsb9PfG3wimhoIN2yuGDbBwFTFXeP0U69TezUH5mRje
IGDE+72zfcnoP7pYrnf44HIUW9LeLCwVejN+KGN4a4N2HG7rBPei1Y54aMoQuJq1MwllZ/by2BVV
t0qJk7Jk3e+AuYyLPR37MeG8O4R3QsRaCkceOnZ9Kai4bMilDZERqs6l2hJfQTU59TSitmtZJfOd
7qf5rZw2vFFOHSy57SA7sPAuEoNQihQyJBTny9zOxh83pdpkDxMJffgK0oqezfddX1CKmCXa5AgG
FCwxr4W8LED4aUhE/nalF0O0sge9TcNMtL9E1Zn3H9YkeKW1odNDCv78r6pjUiVJ24xx8Jar4y3G
AjoHbkqUKXQTsSo+GzywiRlIdLlkTvcYkLM6s5j1PiysbY2Hz/sxbhkiXeiIuLbUwjnv9d/T65aC
BJZyw54+flb0/x6bViuBs7z8LWTFaa+DUxUZ6GT/v/qYXvL0jCx2ejIPntv7AI9SgaT5wr5tNeu/
LFjkwolDgBcT0kqKL7bRaVb0sJzg4SdukTpQkk0HgV2peMGQ2QUXkfgURzcXc90EH4O00y5Nvt0X
ivkTWOQ9MtE++jnOKAi0D4jK/e2EPX2Ct1aR+sbHnHnzKzwTRoXn2g7brP5FPWU3YyO2BSl8BKvi
Ewn0JVxrNieyBJV12IZdUjuLEw4W7naDL6zRIOSDZ1zQK+mhMqq9PFYWzjq28nFam9ftKK6jKxEY
tQrAGyPQP6HoBYZE6BYjNoo7QAph20I13N6OzFoN2e1kOx1xdoMG6KnmMOPUn4wNjHzagepbSvJE
CnlpNCbUHP+D+4PI1QUvJP0QA+SZfFwShI8Pmtdd+cOS/WM8uIAszZZSHIOSfjBUebhhn82ynUlM
7bSxAhZmQGkuj9gO6o16v1UqOPAnxduQzCIXPLUcIRARcaOIFiYkRtnLv+Y8bnqDLaIlAuRRu83h
WoED6rnqWN110YPq5d7otrbqLx84t674diAMHXCLGiDzaPDV+ogyqNb+/yAVby34IDj0pm+UEp/W
7GpPmstBrA1li0DljqSB1g0UYyaLinkqXFP1ntsAAaxVulzSygxsD3pXNr8hYCZ4TikmJH+hi3Vm
jq+eh//SZHSzEfrL72D/EeTyEhmdc7lI4SC4M9VILVYS7oGNlMlA6I7sNaIO8w+rk1PXLYpg8e9s
82VOz2mpqQeVBhc73bJ83ayCFS8NEchId7yhUAJA9x5/Vq06/nAH6na0NpVTuEgXJDF7vNy0MHL2
e6KmXN8SxQFwtaofI6yItuY/yfEZYIF9ngo1XkqFPFUKBn3U1vQu6cALpu7c/CVclpJtI2uhGS3F
HoGs/ztfRXPYJWFNVrEaGDPsfkBAVDK45SsbRg97y3yyAI/Gvhd1w8N4HQhglRP/qXVHodi3Efah
ml6yUDq2vbTwXFZ0DKvdW1EE+JB/UPo34S1zoOh6DW3ifZN63b+rW90RE/+GGjg7ZlRab0mRb9I5
DVTStg/m0NPGWH9WbqRiIM+OeVhjl9nYxOzGqzmCtxdy5zaqi3Fwqo0lJONwVF1YaVjfWqFea/Sz
aCsx1I2CoCOjVKWcItl7J+idyrEFFY0J+OvzqHGrTE8R0fttBMhrzuf+g52ZK9sZ3ov+8xEKc7jv
6Ku9wUGdIXTpW9Gee5hiLHWah988cIFO4hEE6ZOZtlZhX8PzBGJPzh1DnUQ1nnNFUUUL5y9orc+R
pMXKNPGJiV2Jqi0abpRiAFJ7Tt4I7uEnLQ6jzFCkl8dWb3P/+i9GbigibvT4/rERxJYuiTyGjUKp
bkABZ8ynW/eixFwQf95T3xWBfZQv3piGeS4S2LDlYQbHMg8yky77V13hG6KB53H/m3r5sVt7lwGg
G37dzuki2wGu0dyi4vc9TRS4wxMGpvaBUOZ6eo9dF5t8ANCuogutpSamf5oHPrHE2wcoznVkM6aj
sauz+d4ABYTvKInEszs5lqlz13FdDFpSREbH9bK/VkU4AEnCnP9bfCSZKsuCH6AOgDmRFf2+iPMI
vH1bsmZUp5Wc0W4MH65klUJZ5bRTfZqapfSgef+odLvBDOgXlTMXjMOoEcBLjDqOyOfAFd9NnnSr
uacVh4O6FOoDujTYMspCJ8+B+aYuuOiQ5wiyXCCZkHk9lxN2vH8cwrMm7sJFi8cPNPlXrQDVba8Q
XhssogE6Mmm3I6Axpnpx45Jy1OdxI2oNDjf2bJUtFJqFfW3MjCuCImW2Ry3gKDmc+aVrpiXoygui
RaW5gIQFfZe1PtF7TGq7XUyBewePOAK5leeD143lAEei99OkUvu7LqOVWctpH8p8an9/s09QXWax
QfnD3654jTYUvnD1ho9+iAB16B5CCBcUVKvbonTziakdnL3N016yGfbFPOV/02Jc0QflX8aq+SjY
rf6HBRJ5oLAgnuBjyBcmlJw8GFUCu38zwjtl5r8QGiJogapIwBbt3ayVwZJSmoRGscQuQJ2GTaVF
2aEv3VBiUpgG5MUWFZZvRQgh4cSGG9dgkwhIVdpPhMuOGWMOdAHliqnRgE1A+5SChVkZl2kp/OE3
pSc2ToeiVLyb2rfDMMPdi3EuGqUNZpte0/Kl0cJ7lFIYXnVJjo0FuRD+AKzoR4hMFMMZyiPn/f/d
Kmgs/vbqc+JrE4TRaAd8KqjFkCz/e3P4q9xn4Ml/ulcQZI4kbNGPlkslPHcU8ZImHd1m0yWsa8Fo
FyvxcCYNpc4Y/3sc9lLBdgTvM+s2i4GQZHSGJQzHp0eNkGnSvjtLbw3CqXfzOshWi4+Zi7K/+cGz
1whKFC8gGGI8IR7UWm7i+RjTQA7k3zITCmqv+5+1GjfMnPWNXVaOsal0d+UfqQ1WbQRN/zF6q/wk
JczAsXS11/SZA/P/bl2r42RdFijLqFPBRrSjvG9Bj50N37y/Qv7pk2chsQapnO3znvifbtZ9J9Ar
b/axUb1ZbKuUwlWaC38xL4f4Kb3YyPLfzmyUSouLnEsSDWzDmkO6PSVqNYs+uZNy/J0nLpYMPFjp
LrSN1h2mognDEIlFzB7L1ewZtm9w+eraexhklkL4CS4MyfOexzFh17E5d0Pd/9WJ92bNz1rqpMh2
kHOaOdftdMRBf8icuzO8z2/6VIbiTghz6pUolm4rWjYmIUp7jY2FvsfDSC59tfd7Jl6MAjXrn6NK
3owizOH7vYZ2v+7N7H6pDTAF+KXh8FHznbpwuUE47Y8ejE/BEFoc5c1q6ICN39jJE5JLja/bE5gx
erR70g72BBRSoB3zN+Unn8W+LokX18bCQWfVe5cf2NFzvsTG5tt5mpN3hF64NAgE3We2X85fSVTC
SvCCIpa+pFxMbm+R8ahduHzo8jgRKcpaPIkU8eCavETM5f3Fd5VFKHMNGmsdBDhO09y4tG7mTDmf
1YvH55W9ySFAvqsTJC4FApNCIR6M4lALTukbhsfUnJLo7OXzAZGrhkrIDl5mlSE5HJdRmcRVpMir
roKq9X2yr4C7B5GisnVKXYhn9gV907hZQwXa+Zil71MDjefwITMu1pkAoyE3Zeta/mPk2+yJNv46
qkO/aG6TeJlxEzL5Cwap65lVUeiW+VkRCr563TEubzbwPKLZRuwfVgic79GW9XUmJaUoAk+U1iaM
a00dGr/jCKVZxf/OmvlCoLo52RHpigBH9EVA98+Q0qoVHmiBDxlrpuyTVAckQgNOTvDADuumG1Cq
0xiSaVcU0hccZqslE1ws8ragZgkggvpmE85fbxkIS9DhbYHBj4Gd/X0GVkpqQLb04KJzOaWwwnog
kM+JgqpWK6eMIHMHb9HHmbApb9YU3XigwkU/gAUAmwd/4yJwy4eHBO5QURIHwaeSXadM9iopP5qZ
xmi++ofR/Ohxl4R1PEXLaIYl9u68Hhgfs+amqw9VIN1KLc/FXLQvKmd3DjEo+aREOLog17iTXztx
GFfqcjolrGjCULpXZhJ1oWH/0lXdbjY6IVeY1EjA91PjCkhLC0aCMv0tCaUA5Rjoyt9st1NZRL7r
xiWhfAkY64ykpmxoqAhQEMDQ5fu+t0BmelEu2hMllmdxw+02NQaX6X4K0oooQanZwZy9V5ZbCM2z
j/e/LkGuXK9ysgQh3Wl9uwcDkkv7p0CF0/7ULsg86W3w3LENGQZNp+mdajtlX34MuqcMpzB8Ov62
4HgV+aJSZVcDabvbdjQJQSUQDSLgfgrffJeKxjFzqr1b/VsFaa/INiikiY9g59pyDuulvrcmMk1G
1ILss6WFLmteJpRzG9F0RvXEnP9QqCs/Qw6rKVjinThfH3WjyqzUCpVSqEtBg2MPDn5Ij3Fzc2/s
YlBolOlEnvglxGDbfuTnWSIyXINhiBxUHOoYgoa4g4mvvekast7FbAgoE8/6UAoPWGCfVuhM/Lda
0dPc+KW+ZNbSihuNI4zg1MqKwze0tUn1bt+Qqg6pVRqUUC0blZ5/o2OgVBHQ5CaV41vRUAggDiMI
O1QVbwOhy7UOtGUJrwkVCHCeBeVZ/PVfSAZOSUmiJAmr+a0/t1Cr/MrPvUYSu/rzf6PKcl5FV6gO
Ngp/xPg+vet+5uHSigBXCENDK5+ZYc2IneYE99EXSOo8hczTNPQJwG9ji2PNzzENkO+BeNGv3Nym
zyKh2p5Ul78ogWIp6XsbyNSIeRFwauKedGjNgSLPTYGYUDRwkMLYtluWzn/EPlL49k5+Q1A6RvvX
a6oUOhuWkz54nwKJNHIMDTTSNvbWvl/Re9E1Vo1wZr3TupVyWNROs9F41p1RyLtiq90e7WTLaSix
40qPtkb62f95GvL/ML4eWXBZBGTYfU9EhNL3KsUKpnJ5MoTkAzpHHGISeBi5krWZgXj71ld99Z8w
gbb7Gm1Y4BfWrKuKR5lQh0Z6ld/Qx6FeW5L3VKcln/PpE/7Gpb3abA/aX6XDSOeZtRv+EuIwA1Eg
iJzV+4PuKtDnsDZmHOis6KuGRysufzaZRrU1C3rVFRQDavb78//Uje65bQDZiopqaDgbN/0GeOLD
j4hCjeXpKJNvk9Dy91tcYY+1PJeii4T9+OYNQhHUbOkC4TJdCdjIJDPSijHFvk0BMtv+cJed2BbL
YHTRePI3e9ew0x1JhxuY/cL3OUep2gHmV3QRAoRuUzTCwOrkQY5nU+4HNyy1zy5oQ9R7sUCtkugg
zIu+lwxjjEv3JrinxbVma0Kg52wtVj6u1w+JjYAYrXh1oQSlwt+AP0fk0JyAD6fVpn4wsVxqN0Zt
2OpM69Cob3h20RncD3yAmKxGftGRGDZQ4WAGWh9AR9gM6u095Foz2MXjlpdkC1pJf7AvK9vsYF+P
Rhx2LLLO+5YLsygpFEbGXIAL2MY7ztc2GHD6WIH9u3DXtHAJdUY3hqutIVpN5ZCd1AnV4gRk5qCf
K2baqkI4kN2NNJ9N44h5fDz2UmqzuSYveDIRIpbf421370X7x1fnI4Dt59pRlMTlaayAGb01nvK/
7+qq+ETbjfObOiiAzOSVYG1YJhsMF+YGOQseaGemB0fUk2XobMWnQd4PBva0t++Kqy3XLBZhH1IN
A3slYy51wMeP5u0xHRWGiuHm/N6eG89uUrlthYCq88VtddK96bprCYB0ii/8mTZtbnAaEu6ZWd3W
d2mi2OSUvIgF8coYHyHOMeNuU0pfszdg8tzN6WNczWZ3k37+ZsS1sIQUxyxVYHLBVNEL9ZrSZ3ym
wr1odbzkeOvGtackUwG6ye1Q+jcUnY4Fall0u9NbCM7+ggT66b/NhZnkd4yYAhxXn+ue93tL/DlD
dRf+ZhKTKCDu/bvXSMXCiCTBKsdiIWxZaLd3Ec0MQO/DlYs8BQrDNfPj5BIIkzS2HKxlCXURqFKj
dnhFBiYn4agCODRbQtJ2Wvc2CnZn55tOaHmuem0zD+1C68oV1sRNgoqRItjk/0B8Rj1Lt1efftnX
6jgl3kt3RCvMToWzg9AXCrgaYhIyPcecPxJHVTNO5M1PNt38hy9BzzwEhLptnoCyXFefezibjwlT
WdivDqDUkXxtwHobwNAPCtRijNSNFo4KU1VnQ1tkotsCrDR24cYDiwyHhuCuBweBgJwwgFk/g8mr
k3vFv2JxWhTMeJA5F7Oxc53sD8ptiwlmeWnZQW6X7XG67XrGeqMp5uQMOMOE8Qv2DO9ZXor/Q7L4
9zEEUEjhd1g96zhMQf/aYV2jC3SYDIoETNVF2D4XAe+G4weIqW7MRSEapKx95hAD27JFJ/iQOjun
kpZjKQRbkOZ3wSDK8M1hnRcwgMK//wz2IXbw/BGLuXniSPo5bZCXzRkuzPZ4AWkqdHUfA5CrvO9k
CtrCIXPD6plKbTBtUw7FV7/h9oTPu693KvyeTfXSZoez/FW81DWIbvnplU69Yzy1N93852cnF+mA
RWFy3pVLIf+75iBBmbThAebOuwCYdl6YKNKhZCdrIWFXS0g0McR6Riu6HzqXwzCBnPXHJirjA9W4
P49EKGRPOiidMreObv0e168gEFr0r56PFwWx2opNOsM5FbIL6be8X0titzmHJm7CqfCuzgB5OdqB
TaXuJzs1aHwOxkAM4jVcrrbCON4w7nIgf3kNPB074gnsFQDaBhivZJif9TV1JUv8QGqxOhu0w90N
2ztcdeus1lxvbZmAT0svwSr6rrhVXDVQIc6d9zpe5tYl+p4fcKrAUIqsJibJnObRlvECB/ggmooo
xSCrG+fp+KV8BxMHNga3SGQYsyRWb8qGsL7VWyasCgjcoHgCvLbI7Yr9+LFYL8xxceIonf0OIKu1
oWkiW9IHEfZwCUL3M/g845lZF00uPY4kTd3DSKxvmMz2s4djz9NFopxe7s/BZ5ZDEPlUpb/kaGNY
VILLGhTOQFDF8LrylUroERHCCIWqpvaYasPrrmm4TLeWQAYDgfnHpHJaAqFWYqgKPc/fpH9H1HIx
oU8g0aQG46vwMLmdNv3vnwGf7IZ8Z97vEiMiydspWv5FcMdv50ap4SvRUiIVxUmWs+YecCPkOUdz
eBflBAZ3XCxQ/TIvyS+EUpD2Txc7zJa3rw4VNsMh4yp5VVTZQt6EB4eOE0/wimLR93ur8Xb5+cT3
hcOGIJ+kJdmiObjnHbUA5PeM9+ZkTkzvksRY1/rnzpirxOoOfsZuTbbV3l2DWFGA9GfPW1CQ/W9a
JzFndT/v7MxbnK/fPs90kwYKle0LNVK1FQCdWDPCzywvuXBhxTEL+Dv56pzboNliKryYkAe/ioyG
W40qrAB7rYtfp47ccMxBSwfdv64+ZvHG//uzRGMamM/0MsAzizHD5z6HFWGojasauJaroI+cZY7M
a2+KQXP/sSC0yTUBoRW6gBT5q0f7ZEjBspMgK3xOAAssRe6e3sqnhgZm66oIq4XZmkwHcJNB3o8Y
1APaEWFjb5S9gpgPRtqNieALQhLPqjp4g4HYuF1eMrWvVwmJSYFM96J/XRhbBfegVYVKQFJrTFiS
fcTmb+8wW27RwMo9vaNys3UOm1WZ5XCJHdPtP4L7pF7uhxn49fiww6Ts4Mkvt9Zj6aGJDq+IwjuT
pG365EYaVZNY5bkJ9dUmIAt0nHg3ag5DA/mmyro7w0v2wuX/7YoG5SCZUWeYeDl3Gz4LTSSdVtC+
vyg10APjYI4nSRgYjstvSAmgM11Gz/yHhiVG+9pypjNIPoZpM4EjdQaj8cREfamFBtsTYnXASL+R
64pf9DSSNTYOZlyCcK6Nj7G5YDkGnQGELbbmYG6ozpCnZpzUxcICzz6lrcpNgps5CRukhalY9HvE
AqG5Z/VjE6SMLPqKdzmKAlJxqsG2jR2lRhESw1B912O+LgTyFVb0LNHEFmchYEaUdUwri6Agb+rD
ZUClQnw/k62YnJ9bEfTw3UmNZ07zO1YRG2NAAPiss2wzI7WCZSNkbzTW90n4aotGeJ5ffq2ZT/pH
PK5gMr5Z4gKfY0i7vxdKiH91SdkOeB88gH/1X+RsQy9OXb8dnlfT81sM5UCcGoRjJiIbxzWjR+Q7
NvXSeMOw5gTfhA/seS0QJWlUFUnWvvjGyv/VmHAOcRo4C20o3Cbbw9Mp9FMktiWjyP+hPhtFamIK
UrutZUmJr9vXvU/8RDm625oZ4VXDNHdDjvID71Ovmm5mrJK6FipxUracRY5OCkQPwMBIaq4DCO55
/tW/ZvF6C0l5Wu/whHWaUqOxRdBEKq+LFqJT+XZseH3zZUIlWc0w5YRTSldNlSoCrSICIi1AYAm2
n5pv4uHaUHYCKdzPcfsMnTSH2g7WntW7SumzMW0hFOgwfL8y+EFW4LQYsUxJhPmJVp8RQcE9PKEo
44OlhuZ2fK8rlKEvb2zkcnezQE8uDOLefbwgCc4QIAjsmAtKDXAUBPh9GHtqbR9QA1nwCqmG2tcM
sgjF0ToHsCAiA2Q67D5mQ8uIeaM2IrwWd4yXilVkDBGN3aqsqfqCgeBDtzNtIQi9WDLygf6udOe0
6UeH3QNxpgMYrYPtqmChr+6u0Xsk4bWjv2RJ9wFYsIySCqwhVo/tXYsREIQSAwjdjswBz/K3D0pF
eUtkq64o7eCQmaB3A9Ze3c0ySIeRmjalvZw6WEwa5/5TXdV47tQmLUglxqFCxkaBNAaCDhk3AiUJ
ySBvh511ZjxeCvqzynmbPhSSGIEUsP3BEdvSYqJ28B2tly1P9Ep3EsrJ172KX7wKpvNYW8NSBl1G
QMK52q0bPUL2iJVl2eZF5W+AuIkWDziRvPaPU4NWQL6vAtfiadJAq5asqvlBT36aFgA3jiFYTXn3
HmWDUXf4mrN5rBGqbfwgLBADELVFtUKURKcEBqIg/cEqJc1iQdh4euMD0CcfNhXhOzDvADKuB4+k
RowDA6HnCztIDEmZZ30CVboR6ZtnCW4MG9GPTUrX8EiFtlARcDHQcxoHDjUUrNlunij+2jEFEqrm
5/ahs08xm9c1Y/PIibOfmcsXORX2FFHiEZ1OfJoB2Gsl8dCtfVo/f1kF0RBL+TP3DjsfP6x1RGO7
Yd/T4EHmRUchdaPuKKEkGjKX9lSZG7hcmBXpnpQCClzBiZbf/rbRQ8EertCMm6162W2fb4lI0zuX
K4wBQhQhyLpEemg3gP7YeqrRkehc0OcNgRKUQE8sJUlvUTQMWQOs7F/JhZAKS0Exz2rTqSjlsywq
Ip+ppgfsAb713nSZwfRwXxuQ3NaGgfR0V9Rn4Z/bwBE07oT2IFa2ZOk6SEmH37sqKiliS/Te9rax
ziJcMgWgtJRH9U/aPzHa8X5VHdYf1pnOnOhuUiRs0nhRLpXNLIB4jzcY686kCY+gou67YK2fSxVu
v7rYP06oSuyT62sByB3fJNHg3QqkdYa92FveGg7iAYrMMCLA/2QzV0MoqLInaALVoNbu6fQqJuUX
s+Ga97fVfjmOR3Hi5SF406RqX1K+upFjZFxAIMDQttgAjXgQBGhVtcIly5v/BIQP+c/aASc+ZS0D
L4nYL3Y3I0LmKUYf/zYIBibawzBIT20sS7y8CA3jWQAZOG6aah93mdQgTCw6MHkjD7/C/kOGG7ye
Rx8umusxX1rKf/2VZWRIazjat8qpVJlSAdV4QZc+4lit5mwmMRJqapMPeY3cMZvzloMzzRHMDtgt
P86sBKL19KIsCK2iM4zN+KuPTRMMYsnT8vAu5I+1NLB7DYsXKPKBsKBcxnK1HQuXJwt3GTkB+UfC
dja9gNOrFmxY56hMfGP4aiCwsGJIz6EpvdEu1pxzYeZiLnmrB9bIPWpciSLEKzkmL4Hkj24qSn5S
1qYgo98iFBSnJKp2byb8s17PsWBvJzn8XNWOiLWp3/JFXmEKdXt2ce35OJN7bB3dWWWlDRp1E4l+
OCBOQ4vZYy3KWm4Mht7dOpv80pYjJFk6CMdCtsQcGhIJwsDhqnvxdjdQ9SFosBKm6DzgPBaJo4kL
cSCUEgMGAn/46IQjPHF2yWTOcJflC0ncOz9hZfJ4trnpD4cP1Zw/J9z+wWzdeTEfeijYrtn7x9Bp
lV5x3NZ5SkgM5JndbBSs1vyEYGevvj9S1LsPPAQ2IVck7JP6514+gX1MNg5kS5oBszIZT7sT/Lvb
bf4M3lwA48ehYeGwm054S/wj4l4GqD8tNsgTErWJ/XwN7qftHl1y7GLQ6ILkhdcEd7jCjcOEavCS
Dvicgv/RDm1qV/xejaqweRdbWAAkQsTjgDdJPqqhJIU14K/qE36rSYPaVTL/Cc7V+XLI5jrBQYTS
YQ60fKcFBV32PFP5bXdGpaJnDDa6/oJ/sbveI/I3COuj3i9rFw+r/3BhJIQ22vhxCYWt/UCItwSj
JtKfTIDhW95/bgMU22zVVUTgWKDjOcWXwkagMqzNOvEb/X5sBKG0xuoS9AwHmqNSAitRDZdmN/Em
i974YhiF6OJp5nK4dJAapal/00ApPUA8zl4fDt9wgYOmdrvU/tl4zTEFBCohgAS9Gb6/rV8Yvdim
0upTAswy608N+BFaTly62Z0ucHIvWZ889folxxgb7dVDsbFRqboOqDJjb9c/ZAWHcZ4ejG/OrWoZ
me9VI5kVrXBvV6u4MC36o4len3PpaXops0VyTUjRJ2CbJVw14mYOdr2kb1EAdgeAqyQmCkqhKB2y
iCnmHf7afDsozQ0y42K4fbdxclZqB29F0EPrnqwnXmLhpCLA/SrBrl5Y0lUZqMzy0CJw5W8d6VEv
TMniLl7YGQAVs81lXQwqhIoIYFCx5Zfu5tP4hxSMzcg++y9tzv6GZF0CqRE8+3yKErxGnwsDJPLw
+KhgbR99LPv6QDQB5gCyq75VZAQrbGpjJ4rE4QsMH9b4av836QIx2g+nxs32v9S4fTHY5h+bk4p2
SB0ig0yXrX3HQ38yVk4ocyy9t0lW9Lqxxj6rbZqxIs/+ACFAMEXfvNMduS+apseXFXP0Tdp+jopp
yBaw8oQmVQ8CA1ojsGm8KCkj+V/VcobtIGDLrhN6185aiKL3LrbeO+SKrWqQESg996V1eaf+KtJL
NlDxGhn9Ezxq0+RITrxF12Mfh7SKFyYf+MR7GqArzsqe3Pc4lqJ0mezzDeP8n5+vfxQ+wtAY8kHa
yhoI27wkqBSsRsnKb5b0kcuMqHshThZcwP3c5Ig/I01ccFhYrAydi6iXkgm/uTzQQkRCL+d5CwfV
XRf/t7/w1y6/vcakH3VPeiXxRcahBg0Ib63nGLpeIjwZo80MSf4LYXfo76pgIJxBlTDggkPB10JP
2q7BmGoQ2kjmEDeR6/ZBWy24ShJFQTWn3qwnMW8oAbtmWtf5t4oObmR6kIPp/pjobu+zOUOeGyJB
PecKb8EEfD+KFI97Rc3DEtihOnfn292zs3mf63EG9O3Cl+5sx0D50fUugTA5wvH5DZN0BxeGCU82
AGPRMG5p7p8F5MibPmLKjARpf5oecq9KXNLURoHBkrNKkCKtHo90A6ZHtkVVic06SJKH/EKxXvbJ
Ih3tWH/a/cHs804ff6nGSYuGIgiY8i79WGBhvkClJdghAvq8Bj+QEO3MYxIvscNv+i3FRwmJAV/W
O58QQ+WJ5QeJYC8qiLptTabKvBwnAlrfWNjX0leuBEGGkP9earCA6WXbRBQhgLnfn3NbPsqOIrZ2
yaolpj8qDHaR+fWw1HGyIOf6byGQ/r3lXxClosb/shABjRtBcyUUFZ+2fhrHfLFh7NUyqx7mT5tV
JvrNY6UWG8xSDkJUd0TpQ0W/6pRBZJP5Do7Dp5YZU2nbGZSMDX/RFl2gJ0v94fyaX5Q0nhWUXQPy
iRZQ6wdZjFiSzCQfnMspDGOh9SjBZsS8sOlnxcljYDTfBWV2Wl1V8GyDdeUopb5aANih2uvA2FRW
WlU1hLMyY1FeZsDvJV2naXPCRssPTxH2TCsSfUBAmh2nqc0TXXQmBeZBFExnkyyDl3E86u0CFXyU
GBjlXEEJuxNrjjsF6HaR+D2RRLO4FaVLPb/B4d7k90i2NSSrJr6DORjWykwoj55s6en3he4Kn/nH
Cr4ZNnhCIuiWqCQoqiFfb9JZFPIsQ6+Gs56Dr+Asf6dU7BYKARN8azvQD+jeT9t89wAaiNvwPt91
x4K9Z1s91eoR8f5J6AiHMl8dQAw9qhNDl0J7jUloxOwCBUczE7PdopZh9DHU9R3Y5REdhOB3FS3n
qQrJbHu4xGj14yUSDf68Up/JXdH/aruSnAFrgNtwFQVvCa/6z3E6GQ6S9EmADQTq7A7LE0lMn3tJ
k9yhrqIQ23VPjCQ3sCWICJJkXjASK2cFdxDdnWvZuDkW5+iDrz6JxIok2jWBQBk9u9yfCLI8OffY
ZbS0jWHddXTcIBtxpCigK1hcUz9FLzExO+CpETgTZ2zBJ6eyYsLLCMKofs3gLjOBCoAea82HDVgR
k5oIK1NB10tIGGWGUq8i+9I3BDkZt/Ob0WfXeeYTvE/o5XdjI3pkNnz3gJzIMdIZga/NLAnUAeq0
eULyUQR/GOuAuSj6yihj3RUuzwLhDHEJt34dIfNGvX83zE1FPapw7AK92Wka0tVt5nn9BLUoc7g1
67kLxDPhAfVlbN52fDi0QbN0D0wMRdiLTtGhPtarOoHCdEYLJ+EnbttAnQtjs10oxo6OE7hM4UFP
P4fo77MCVWN/9jkqITfJUoZMBBqScuElkE7kobWnS/p1bKeUWU9DFZPq/DApSl0WZKocv2lvMuUw
fsQonaXn1Z15vNcaatDvqciw+562WY47u0ItIsuXdauxB3FZFJkcXM3Rke95OILiqp5cQetpeaGS
0deIC5Ety9HXQ0+aWsyRZej7muIn2ALtieYeAtV7w3eaE78lPfn8ihConZHdB3q3jHTDPiZuwgFz
fiMoHp+ndxrJBOHA1cCxXpfdxKxXml9aFsYztgx+0QezFbTs2cWI3Wf7OwWFYqKg5ewqT3ePvNlN
7hSinDxSAI1YDqVOi6MtE2wQ7zVOIES1bSkuLKfCWVahUZfUvMs9Nn/Qi8qwW0Mf99raCOeZi+G6
7u+tpdst96tvN24nEL7w6DTCl6SoaWclxIZ7WHPJxxZsDwBGInhqgKHoN9Mo4281+/ucwjqkw9iB
smdh9Ch0/KyTll2h4Nf9oBCL8s/gdFfdrrN00UrfXlUysMwPNymW5d3DFXRhOXIVo4bjSjOoZEBr
P2ycFspEDQLgJN+DIus2e4v7Pwaz10diwWH+TeLAVr5a9uPL2Q4S+QxkHapnIoGqaZwFkhcuG6I+
FgCowCugcvK7lMjqg6q7zLk0Gm+FOrtT5RTTTCK2eypByl2sHtkVrX5+f5aqKkm0j+lbf3fLPq+m
mOAVFe2IH6HMRvSS+y7Q3D9/QV1VmQh70k1rs5E2rcfR7/kUoCTePH29GCn4A5IJU7cCvMiEMTt4
cIXcrHEUz4SI9+7LhUvQCroNw10hRiOuBiLV/8Pg0Va9scWFLSpGslmVFea+LthZG9Raeuk64prn
tivc3Y1gfr4kL0AxNeNDf4aD+QjhWQzanQrw04El5kIz6OcmKDIhVImtzM72fQ0/xYymML/cQCyy
XQRrCYP0JIYLaXgid3G/sBRlHzq5Tqvr5kxslvewLT/WK1sJjZPdnsIKiDrbgJKfq6awjnnx/tkY
Z+QyYKQUV7kRFj8qok72g98WyRWp3TuRDJZ4yUPnLgnfKgMt7k2qexTOn0N8IHpwGzFk4FcjXfXA
8IYrAev1dzogWy+Ws7kgfUX8VPwewsTOdziaH0AWkLzWEgzU+kLMfvPkXYlU+pMAEnfCHPHyB/eS
jymN/MQz6oLp+rDpcYoq2KoYKfGvQNaQAE9DNJpxsUr1JLRWAvGvV+8Hszq/JBRalm2Dr59inmvD
Vdov7SQ+PbIBzPEPENOtX/CXcMV/ZgjrJpTprJOAGj3Vt8uSndqS9OWLjDNMMWenaPipYCu++FuT
20wM+kBWDKDKcEB0BiGEliNZW3jyhvEWrj1PdCkg3zbqst4LML07oZ5hB7T5rd/mrMaTOG5uH+or
KwFJ600IaXfP3gVy0SOPLHa9tSEkqjpR6ND/7XsVFlj6NvyyHBWJh0JF0r5QItnCLZJ/SxeIPFK9
dlTokJMw9nmA27eUdzcOBKjfEJfWFdGErtLW8STBGfAe0J42JBMajIZbSck724MOPHQanXgyuVph
Yf0LdVyYIK5c3qTxfH3YA6BvSFRp0Uf88uMo/HZ2tyV1WOiF7RxUQbneKYB+OtEQUWISVq2YfG/V
nZRhJzefDMz9jIJMk7i749UGN873AWwhyvVXc+4pgoB+xADzac8LDrU3w3e68vG6OqFEGzJewj5l
F/hHpMSPAuaErQ0k6vVhXJJWCR8q/XRiQDs5iMbUtrVPCyoZ8G/Bm5+96e39gE/KklCoMARGFq/y
uXlHpJ8haY+3kSmxEKkXWeaXY2Rfywk30sqYgMZv4U+gbGdIUGyXUMDohnl4nhQtW+I0Rfn8cfbs
kTZ3bEzisnh9hViqvsPbGEzWIwqhBvx1hK3RNQKR2LPjk16AcRMlYAF7prdaJ+oFQSkuyxnqU2xF
vMGdeRQGXf5I8O9Cc2EtNBareYLEjLeup8pGpf350AlFlva6PKalqi251tAuNYz2GLdqNQajPUYh
QVQCImtR2kvE6aWphTOYeTp2qBAXcbsvQ6an770Liar2oZ0Wd5JY1efY1Ge058yOfG5Zz8hT0FNr
4GqcOAmJgrHC3g6SXgR/zW9ltsxUddURc5G5w0oMXioUs8mVi/krc1FHv3dTiRsA6ewgF2cqK5fc
VOlVHOEw7CsEE0qOb0y5w4F9UF6oacJDTbB15il11gUo63EEKz1sTP6l0nxPJX3bAulEFjCQsxPp
5AyIUBqJFmU8afonBd8/iAOflDhYpozi+pWB5P7mx7/EaEnUREWQWQLSFN6ib7LnYGOFXAyqSC4h
tG5wIIx8HtbeCwmd2hODQfBMnNtdWjnalIusQDNSr9YkQRqv+zCB3hecab2v4chPiG2nsn2GYXje
BvAYKhj6NeImjifHauRSIW46qS8NU2STmGprOP87gUUMuANgsTV6uHkd5Brhy3G1jY9ezMimtXCH
8DfQq8qRbvWBeEaDPxqj7qHsdG1oRuLksZXncxGIN85JO0O3rFpaUhO0G6G++nhboSYYCbfzDLiH
ccHp+EgEytaQuUNtJyjyDpMscVcni6YyYuR+9F7B6HX3xZpwmJyHJk7faehQMjhfjH6M2WtRwMX5
6KqWH4jGGdJQCMHIBak6CQuvAYN+FQgs9KE2fIUnclfPalHXLK4HMZngQQ0e3ARs37+ngHSoMW1W
jkVIzeWSfHE9MHAAA06LTuMW1JeYLCoi6lWwe5jU8i0/2s27InjwZYDILCrWNGdF1ilp8Q+4b9TY
6Oz0g0j2Clv76jVlwEEbiMrRs80Rwx0v6LFv3aGgbeN1kXO6kuT1lhPGIg9L3M+uTjgtO1ujZRLX
scJnfiGLbKQF7NEWd2wANYfv90JLYJ6zisHVfhAm4UJ7WTtuanJLbhpYsHUylLSsZjNgvq3y6Eaw
BMu+YjeslLGqVcYZuTUtORl1Yo91SX3aYaaf887FCtv4BGj+unZHFJNu4Tq56F+U177TgX2f6j93
3JIc7en69pVK+KCmr9b0CMh3NfwtjNxWzn9qWP8BHyfKeRHfKss59gEuV2ZGHXV6CO5ygM7Ly8e0
EZRzJWJ7/kla7FScgvSZ2N914qS+82yU1GKhySYdjx7b8HZQQmsnk6wm9SCHTU7QhSMvg/LcHFji
p6aJ5GzYx6e2thaY/cbi4Xk0Nq9oECE9ytfRGKnVGnzCFPN/UDEwF2aI2+We9fDg+J5qhwpAOon4
6k1V0eBFMZspqV7BNA3dbxzcno5KgNG0d2Ug7QV3Np1LWh/o9oU7b2Cl82x57luBpC4pPXWnxATv
962QdYAvneohwEIByTVS/ZVopwDyi5tyTQNCEgrzY9Yp0fJY9pP297Ry6g683KYkOrA4sM20wFhb
x1A/B/n8feHHqhjTlHNkdcErkntshOFqjaoMWZw9yY3iWN87IY8700MXB+YDKxJc5lsQ8ynWD4K2
CtwIuoyDH3dVmEjfyV5ZcSfF1WWYjotG1oBLOWsuB0hX2zcUZrbPQVuryEX7qRpnQdtid0zRmeXc
kg4Fju2TI5ZFrNx8piWsLq+vra8qYj+jsYBJfTHC1xwvACuR6YQcI7jjTqYjxb89SZvM6RjSwu6h
nbLhECaPV0BIbxSjc9yeksAVe4GyOnQFf870N4tLGXW1zbfKdH6DxL5vtQcE1SU1E8hIU032Iq2s
FG3U5DzyMp7kJpv7EHFTbZBrWiGfxuMLvYwBLfGxESA0aDDiEASnZf1kdbGA6mfv2LViBvOljOgu
Rv/f2da7VnIU7QOeGeuy+25aW2W/BrKhPxq1s2n6lUfng8HdBtrEBGWnPaXmjMFsS4E4Uorsw9Qy
QHqbn2dt8DbuZDOYedmf+fw82L4YyIHwXabJ4iZxK9GZrUMDw3xEBftFWT6G8NW+UWXCuWXhKaGG
7xwHXB6rhW6aRPMZrZt/0Ux7Zk8XdYfCjgG4COY1p61xFqyQdCDG5shsAAo521ntzMZs9nx6J668
p+tfQMOx1HywVcIx6ehht7xe52F5MjPfJ8R27RQlsDKF6TUIqS7uWoPtOTxiIbRpB6Vxu1AI+Y9z
GSEyfp9+HRFi7i2xn1MYsW/2bEoWqM81zexWYyqidmAgXcxHhA7q3F0nFy1DCbaSJ6BWImEgDh7D
zgMwAV1wHW4hgPSxhKyCHd5XIpyndcPs68kaZIaww/P3fjCgOM2Kfs+ZntrdKFsQeIRSzPuHfKnd
gXPH9qynDQxEjyVsA5qZyCshMf9pxrcK9XMc61qXdUve/jRkNKSHXCa3hUaBM92aSyRmHou9uQoi
U9Hy63NvNL/NOOY40mIrvFiCxS+UYUnnNjsadsnxVrjkWp7Nh/rGMdp1VOVbLRCGHeZWrfPTgzN0
MX+Ws8n3CLXOD6aqjWGcjX8ZHRSKqAgSlrRijJDRx39FD3zRHljkwTnB5/5b3xK3bi6nLNVsPPTh
+7bCm18t7k1WlCmrGvqk834BKyLp3aPJ2UN385oO1aC2fbPun16tLWzLzpPG7ME3/apfTvjSHlru
Ct5tZGLMA73hP7Qe848Ec5l8B6E/oUjeCqQSW+hAQ0jEULa/1TlYoTGgF2itymjccpCeyGHXcex2
y/uGyV4hVpzifdYKRU+SQnP/1yMOot0mmnENEowYVT22grhCIZFD0rTl/Q+1d0QOk4Nu3MFTdiLj
OW1ewRkqR7ou3Y9j2LpswhCGaBR9e2oax1g6WZU8PAD9odMgzPc3gW+AwcvkALRYPUqWPS8RQ+Fg
3KBtp5HNyjfV9kqnYfjKYLuaNrU9O1h0ustgIJX4Hk7Biu8ZsLeOC9psgR1nRyQj+n4+4rHRilIK
vdG/1hOptAbzwhsRIXRui/OVEYuCPX8luTZGrzlRGtjEGnLM8/43OZUDqU7jRo2yt8J24AGOGzUk
rcvtZPWhK8GJDT2Rfstx7uBHUMGFjbaVd7d6Yv2dryHGtBRPZ3RW32L+nw5GauC5gSo4BoqSxpv+
hEXFPNp3kg/YAZjKvXuTxqWS0Js+aBlcMSPaWcT4Si8m5cDEdyt+chMQrLIjINRiOmgchZUFKKv3
UxCRKnawE1W61t8J4omTdArSHj4CL/B1cZZxkoMvPHLlREq0A9Cbt3eQY5r1L69UPOqeN/+0BXp7
cw6WrNH9C+hXWmhqahX71ny/bvTZ4cb/QA8RRdybF+6lf7aUw3ct7GTavroH3EQHZqNIo4xC1RIU
xGvfV+cuiS/njrKMA1jT2VqTOdHRAFD9NcKJSD4/ezae4+5Q69ZJ4EqUlIWhoRkWZb/3w+sq6JP1
/6RHUEDRx+yst0akzxDSysZtY3YZLK4UDu2xkzOVDeOr6rK9ir+DIUHjzICnZ2tAbzr/aLXXV8CW
InGC45GKblTxm1E/s6Sk0t/Dcr539Z/jmYAa5N+sK8n4IxIQX+lm4Q4H+AvcXjDinYYvpR/oCYul
0OK8W8JK8YBEv6fvHbMMlTPCN5emrNqAApRJSZJF8AiSbFCyXMo8fyhUxzqUkg4zn65ry2TN9lx4
FWcGdB3gtbsfOVJvJBuIW3D/dAawscBwsDcSmlUNg0eWzkruMhVHu7OBCy6THntgwfMqxU4oxlKN
F1y9EhHkEo0gdaSvLtbceXAJqN91mJX9JQXuMw1fq+ecKiEXGOp344/ctHPHnQ9C94SwAU48qXRE
grqSR0XEDM7YFWEvNXrn6tiqNa9FH3739BS4rrB/r7qHk79pwRdHIWlmldw6bUR70sQCE8I1ZNGz
9X2nEYis06AJ6W83Gei2VnAyQkUaKd98AlhgPwHaKWImi+TMM8imYsXWyK9UPzi4V6mgMt4afkzI
FZk+SLJ3VGbLnJEvtXeJlXB0Oe1w31lTOERzQrPwRA/Z2EOKITREpeHititfk8B5ZeTzl5Cx5vlh
LCvkj/NO9UKSV8aG14mJQ2hSbsEx5cbZpt/QwM32FRZQCcrwZ0bKAaiIqEFGqNUYI2RVle1Ew2iV
//XZeYzTSuzGsggxJ9sU2vS7OXNmi4kCpzRBfjFhN44iFBnmWORzKUNoWhXNzgHjSkqzUH+6WNb7
kXAcgkEj4G0Khfyd8jN0wD1dowq5BsDmiSnGC0ofsH5XAYlCTlLzONqXtO1lkmCzZRu8JQfoxFtB
yi04FCl+W9wbIVpVWG7i9OEYdujulub7CeyxO7fUPRrcsLWF4FdmNJEcQcRRKt+mz8LGfxT9bdFT
V4UBwxYw1vdeCEpLgAodr50+1AqFNSifUtqrrgO6YLZ/czZKDt2uZ1Yw93seNRyU6vBQEEE+q0Ru
j7EUBjdzC8870OFash5qR/gfQ3Aw6UVZWn34cYZ4IUiM4J5HoJeFaI+YCWorkBmKDQQAWrJACTJn
6sVQ//hMX4BdDs5Q+2fshbATmUwCbOq4zCHU45Ef4pssAg4snIHl2Odi5wjFjVok/6Lp3mBOiLnK
S5qt4w4XY+qRUsf2LSGngCiVaa9wvQbiSwoFrzjFbDjKDJXc3XXeVy9S124qE6vM2eKdhdC09anT
8f1M07z2wC3cPM+dE5EhtmL3olWJFLKJrhlg/tjBOMPm3BEqCV1/fdeaXWvw/5rN0bWNWFQU3n4J
E0+Qg+fi1NObrbo8l3nHiI2Y91jl+p5Svr4+Up3/rNnlusJXFbbDjgCByb9t9JFik60QBKQ5sTeB
/52RBKs65Za4lcGBECN6qEMr+W6+9V1WinN5P2q5zi6znTvoJfavW6kKiOjzA51h0LWu/qBTHpmm
f1Tntat+5+nGhEd5JLd6IgZW5U+G0S/HBTZBoR2+ma39I7PIUhL78k1iiQ7BH0zULUO4Rbd0e2uJ
brooQiU/mr3VVyAHN0y4Ds6pU6g6pa03u/j0MgXvXnasN3X19K0pGroUkNzfYceaRzvH+P59ayuW
sIftJqGFQWeElBEmfWDFq7+tCxW2nDqF5Y+dJSDCBUJKz81nOI3GWJQBn/GoXyWGwvGa45/46jB9
V1W222EQDBp23sSJbNirVK7Swi5PYVuUmxeUFfGlqYpEYIj8VSwrAEWJFmtU4TMFyO6Uv339evwI
U3zkf2aKf9OO3DYbeb08xoZFe/lL2iNBe3OXxANAjh1q1js9X0VsAWJjtLovFSXPWhEcM/YI0xsM
OUXe7YQagaG/IuY8F9h+8fyQ6XraR7XJjJj23uZCt+6qqwrbWo1EWHOapImaarHYas0EC0dQgjoa
VYJRSkci88R2Jgr9WDR9SxfYFshMxkEJ4U/HXIG/TuzFEiOYjQG5zoM4XJhqzFrX2zNUWzvFqs8B
U8zqmgWSo90a8QDJs3nX3J5QWsk4Mv5PJ8LCz66edybVVBrcZ4QGIw2FiPoSlgs2GLKSgCeRuxcS
EVTZkfLwm2SpwXFjDeNu0kUmxEXjLDWQM2+/OyprhGZepWw7dsssNaYSYqUxojLF1MKkA2u6LRsw
OPz6M1TdcmV4Wbg9lG2XGPwIIq+DQeY/sP/oWsq08PAfPi+f+QSml05XQhLyQ0pZbHEYGXxGglUm
vt8xAbhSRmmanLI+JsKfbiboaE+Zrzn44isYZxXSH3UuAezBVpt7bjhu/sUWmsnmcKonzlGcT0YM
TWz6+F3sfMnpV4XF1AOZLmHw3ba4MrCSTkRX26rEq62q2fi9YZo8CjyZTAu/kM7Km3QJfLFVVTt+
CZMBmdZ8DSoAjs7EHK8+FB7m7lQrBlKLeFJOn2cYk5q1RZXhXxPBiCbMjOFTvTtnN6jpPkEhcP7z
34iCrnH94xep3NnUBGVRNGTdDoh2E3IKfhkPMuFqaFg8mYX4Edp+UyMoacFxARDwUaU2pr7Rq67o
CsR5yoD4K1GnP8+Kg7zyOEZjvmowK5MsUBHCSSw5y6X4xMy+95bwnT764OOk+7s1UMl4UOpAfmLL
iEuqDaLvDE3AWusmAhE1mR/uL1/r+K1bV7yeY7QQ3iy2a7l/Yznr34H+ztiP5ObJYFgTDVOPSopt
m9yvWKueOpygh8mwS7vWfm2cPaxxJE5HcZ28rvmU5J5NCGFMi/8gCQbxaH7rs4MqCs2B10cfk1TF
gOO6pPfEKRyclXHuAyLCrayPSlzBFcgj6H8o4OlwKlDct4PJjXbfz5YQf+f00MnC+caLnRQXNT0p
tJ791g2sWi9HycAgtHYM8GA482cQ0/m1ja3D6UipSP554oVJmqyD4oj6fZQDRVGfjs8QgxkiMm6o
1yVLpVDmdzWHfJupzjiTK0hxjb0vs8HLSWk0x2Eo0ta7MvkyaR2Tl2r70OpS8rX9YLGxJkJVwaR4
c8+zPF71e94xLEU23QQUftLHzz2A64zYpgGkKgV6ta6pU5OFxZVtZ8W2Nh3/zi+lqH5QF1Xd2/wZ
ntaLxTTKgTKWHlOlT399TjiCrPS+MvVruEqoVRkFb+8T9UMG0S6M6f1f7IAqdfxd/QPsDIRSSLT4
AycTWpfHeFL3LRlaMK8rhtNqBCmoyVAAyqs9F+MNGdg8tEckUKuXEtVIrzD4ibizRjeM9gjy0dS/
BPXkQ07aqZMCG0qw/5xnmR+QUT8S2frvEt3yizm+1agzAQyhQWbf1TXjrt3b3xsxYvoMpVY0ZI/O
KCRhWCoHUdyEcVG94TNcYQWNwbicZ9uLXa04ylP+fHWJL2wNYj0G1XlQQhWoH46fqKI5KjvVPjJ6
UslOonVng/cMTL324c9nvsOzfFcRWP65JxNU8VunRle1ckLJhLNM0ZtqBFtPMrreNQuehsqTuuq9
l8pNCibmDcZ84F9kpg3xxGVBHhI/L5w/1T0IadlQXUkfpR9MiB5xj8MC1LxFh6opLE9j4N/jfoVa
qeMFWx+ie/OcIecD9EDXmribvb7/Jzfft/Ifm10ERkfXAycrcM+hQBclkAVIfI1rk406gUXNQHYh
cez626JuJP2TxEBr6Ye+huz7Nqk5h5RS2RLBaPxLmsdZjZNX2zpNAF+0YMz0nzFmSshXLzwc3yzk
it5NHbb0yGtOQWvxF9Qtx6YVU+A25KYVv8rIOufjKUCkMRTu409Ky5q5c3uyk3wqOegJH82AcDKa
gbzUptT2aIG4X+QuRXv+FWt4SHrcf8ohaOgxx0ho0lpOVv5ShKfz6pt8Yg86jWvV1EK/Bpq4wQPX
al4TJAcSksHzYnyDwRKsd+rtXvZYQ4U3m5CmNLOfE6xx8nT3jV7vyJMT7jXowr7lTuGnLjHpAeoN
P488DonzoBgnFKX4nXnCKiiWJ87wGwcUsSfdDsvggiMf/bDUwWSnBdpJnOk6Z1wxFW0ZW8Z5jvR2
97pNURGsiZvBG2+SUdB9/nFSvq0dM8ubbbQM9H8ZBeOvfTsUIYtyA08FRXNbPXCi1QXSloba4lwO
H5SdYKZV/Zxugin3xrjPzlNMCf9FRmTvG/tMQ+HtzE9jm44qL6VP03iT6orMIeeN+PMMQWmjRpQh
mO6iKn/NOhEuPO1O6n3d9SqeUUjdeO+IMaFay9Ahe0PjOvb9Pr66R2lLh1fCNMxp0P4mpXSp1MZD
yRfNYtICAo76K0D8FRT3a7iBM+IrPceGCBfhv6kRseL7p2plrGv8dx+GPxxb2knNuA7Eoskdr8xI
AhJFotHl1imyWn6jF3CtgdXtryhDVmN9dNBnunfO5U1slq+SmIH8b0nrukRDj6LxdI0MAP9j+zvk
7Cw9H0UO/AARdekla+6nY/g6J+k+ukZR7dm4s9egSC2cwDWG2bLjDgbAVg0g8rjMbNGbGnatTaM8
+7ixL+hL7c3Cj0jK7pm6y0ZmiX3N2CoavKQyze+p3f0FmJCJ9M/H+aNy58BPdc8EM+AP8B2KbUBt
Biobemzaet2PLjyY/Tys7WklfoA+VVUncO8uKGkvDdbuYsfJZWrUknnCCdhNoLnzulXdqC8ltjHl
TvpvYxS/dZtaTan+B69RbCmFhZ65pG83FsqWEU2vSCOhh4E7JigOTHBkF1fbRETNkua8R21xp3D9
CzePzk0Hc7xvrMbvkRAzvJ/vsjtoX6BCw/DOmhWhB7FU2OyBvnkeOCGhjrW08Yv0yuYKbaDZvUw9
lFaDFolbgP2E3hLFRb50cjKD0z0gDy613IvAFCmWa2bxhlDXQiUHDLPeXJcCd9XqHqLH6nvgKIPa
HP9WsF3I3eVIRrO2Q7wCwO6RZHmcm8I4QyzlgL8Hk527IU0cf6gf6vkS6sH+vkBJOgYJnrwxjIW0
3cFGKu3/pYj5SOVVSxLPzGIw0DnTVKwmXhVImUam9Z3A5tOZLDNMnnHvv4gGjqzp+rP7jqk8m7tr
M1GSQRuA5ED5ptHGtz4uiFE97HzSwpiaFBVtlMErILuwFzTy/B+fZhkIzYwMvKk/2rfkt06JWzI+
PXE5C29wGrEdbC9c7hKCVCXNdZHujXBlQZ78WyU5Wu/zAo7V6PVZRZYTjniiw1UGTwQKjT85Wn3t
92gjLG665rpiwZxEXNHiFCI5J14cmxepkYMWdxGNtMPLeukHTzixL2FmRDo7D6o9xn066MvOGL6F
xEfixha3Qd3Fyphmisn65Y/F4Unh8hSKjnsmXWcsg1aW/tz3ce0mIo9Ld5rEI+4ps3PAhOdZorAW
kfRunnuiYoEOaAgrcg/bCcmcYPYlRGLci/ghk1Xs2gFhd8SfDt/denAWSsByNqK9x4YFCIeEVzlj
9wpihzbS+2SYSeN1JVEmhoj5TDOxTQ0sCrd6QOaI5tKYcgb29+vtcEPbL0CvpWeHksXDVeGDCjSJ
65xO0MTUbLuaLmD+xIPWQRGcIRvZs3fdUeJUtXuQx+yjg8ygL66XZ0Idq4j40hB0pvvpgSBdkJOK
YFkYX5FL3GR6wnrfXZI7bK5rv03LZxEbtE0YTFoKDvUdPLOAJQcZUXHV61BVf5OxA+GnpzJYaBw1
IcXLlZSKVazI8k3AkImTiw1ITs3yXrqwopRDA/LCXbwY8eJufOROXj0bGlkgdxuIVuC3ehAe2EEz
YO3Wcb1uM8W4bCCxFX9cbzii5TWf5l+PIdh9xTz1BaD2M30fWqdJy8HNjOQrzj/er8+SRbef2zFl
auD62wWr0zANh5DuBIAxJQ3HB3N5ZLYGOpSkFMX9qM1WrIYwDgFHbvK973cpDOOdh9KECi2x0co1
F137mVcrQK/rpP3OtQJ2OT/xaG3BZo2n47BSeBbc4NOswyhEoddnIIM3rpfFvYGzRnsWaUiCnXqE
HGkLj1GUU7FBiJIQ8HskhoZaVAq20MtGmBoPzozKfAVPSTlIMq5a9ZexKbcPeTyu9xK/S02TSCkM
V6kUNLCEhPHYqfk+75hnh46CVOZrSmTrn0WNaElkHBR4d9ru5K/XJ0aWihLX6bYzj7qxH1rc4eMK
0APOlpCrs5oj2TL4YHCUBbf4fMhxIhfoaFWKXI76b4nFsM5Gp8pnAcffURBhM8l/DyqKpruXMW3d
Mi2hm37r5/AfilHjY+BX+JvEPazTyvPnqe6tygQEB5XxJjVYYAL7LZOBEFl+EeBGrt8z6dzCH3za
6k0MSGrovb3xfumrmviMBe+JgMu8VZioKU9gWLJtVLuH3YL4xwZ0dvJVfPhVrB6dqnvkG5/IYOPG
d/Fv60qykPdubvK16copRFfG0pwXudoPcuHlYQZAU+c0OfMj9yFUcjysHQbN92nD+792GmmZu2YR
vv4sOi1Q6XctRJH1UmwZ71NBXQgmiI6j+3lajrye9puxXqTBIWqfQ0E6XXsIF3PL43xp4KpNpDEy
QgatXbdYOLTK0RHtVpR0zGWIuYaCB0r95KmCYPyW2ihNab7JCXz85eVzMjkt/tM95PVcTDiiXHRV
oGC9OnQ5ktJZcOhMu94bCmj23MdCcqJwb0kvGSFmlza5Fzai3dhCjsNDWrQR/vEinpYsdkYrKGh7
lOGww/4Qxlyx98p3kcMVR9VTbX51OhMJIw7TjyS15h7Pz58g1o/sFbK3BQQFv2tjrpcaByrAfXJq
gFwuuKHFeQ200zTeKqd40b/qumNfuHNrr1llL/UNiOJmE7DikD8Soq7vvA5TqKSTk7jeF+yyzZsi
spdrnWyD5Ik3kwoXpLheTMl0vwk5fNMPXxz5LCoNZywExDuGOGkRLi1Z///QQx8KDiT1ISgDYgao
EgU3oJioDLTkGxXMDkyoTbGezj7CYOmOdbfZVUlrqZ0S4FenMto86O2EpcFh7XTdP22H+xfesnCL
NrlcCsW63rtGRST79RLAP4CBLioxzQn9JEtROLoTkkhiRuCpENFW1o05EHMeImn8ciYQMU7fG/+o
ybbhGON2BDfMKpDi4vS70rmtpnj1NFOpSqJ9QffebGRe59VXVyiJhW9oPTzh1BDkqNszGydPHoir
LNFJbWxWKpgD1m8sFq+xASo9+2TYiTD6j43/RCYAwUpm10cPlELdumkTUZ4NoqKpqHuVAIy1Riik
VoU0U6Ii3Sywo3x/uW80uc6QpWbIB+9Sf3mYh7cx8vGtxeGXvohJq2euZz4LRGf9VelPxQfRBGno
ZpjJA+ZBoZ6xV3EcYtpCiV4Zo+DLkL20AZAshmtCG+S46JXw98ngfZIafeIf9Nj6p311uTGP8/eY
G9L+ULn2kZZFVoOTLqcdpAlYzl9RFISAF2WA3S95qxpnwTeonR0cOqeheY3pNSANTJlAGUspHXCD
l7xe7C8r3LziQwOEO+hgu2Cjg7fawtOM5xk3XTBNefxZqgSFozcwhO3oPQ0+RGmXSM3Ib+1168m0
m/LiYgjgS5V6Kp2gHHhnQRNvjEUhi49v7V3ZFTB32nD9x8gpVQr5gC7aUqdJGpXriGSNflaUMBoC
pA4quAUvyUm+EnIz24wbi5jNGrjuHSW0pFhhkugYzQ5OyHcRFm0SR7A2aMBgjUPFwYbKGmAVDKBx
K0X87xRkffzdgmMd6U155qypXyOY1649mynUcCzPyhMzb1cFuT6nV9aXuEzzVLIyqLDbiLgRhdpd
hyhPV2NIH50urJzv9NPfc8uMILi3WcykUFTPtwC0MRIMo+p7QTk0MuSNN370g65LNQ83vPJWnjPA
+B4wD6qY6tNklcnrmzVR+mggzz//hi4I9j+bPGbGpXb9OjSaajinrtDzsgt2G7k6az5I+hNo3y2c
KlPTMp3eaWpwQwmWwh+PImakS82paSM4Y7mgL6KR76zVtchEdl7wy/Ik5gzA8tGFRbKVUOc5/bFG
IdtdMPDtBXsgA8lVbCUVuddunQe5b2M22kGwLHmhx4CHTXbbCwpY3Du14ztbLXbeiDS9Jic0Xsob
aG8KHDxcGVhShrFWy8m7DDua1C/bnVDEDKJD34dLQHTC4NP5GgmjgwRhJHLwVZEWoD88uB6Kb/nT
3d9prll3r/8dV3UQAzOviz7Aw1mRneDCVXBjdwTDx9MiyWDhXSLOnupluvT1yNOVLR0G1vzGPOiR
Kf2LmxhUtFTeIYczQLUvo2gjtRVdrqLyW3vfskFG0fJBhOSKW024bNDe3HJAfDLteDIbU1ehkw+N
06kqypeX3+07r9KeRubxXsNaaATPYe1Hmz2AZ0KoEjV85a9IhoSD+eBWiTcpZCTF9GETFp+35WbS
0X7kV4YaqX0g04j8ZzZ+cWDTz0cL0ztpRO0JIKBaE7wm6maxpgR1Rv5xf9i3/KZjKPdlNIsHj146
9PLyq3xXY+PlbrM/gaYdin1rN5BwWGPqvQY9n8rPUXbgv75LKDNyPZLUvnD98UjVhh+HgvWwkID+
/sJ9TtFr5nVSxuchYWO976+iyGWj8AOFpH+xSsStYTx1CpB0m6OMGO9Mb7682gXFMSyRCFETXswq
pAwZUGvhBFDBoQ4w3sTgd2bm0Oi4bAe/83wPQm6P36Fsz3+GDQnTXpeUUIKUfzFb3y70HboLjbH/
4fiEXMuhvgrvSH//z8vVeDkiCoPwxoJG4s2BU7qHv9GwOKGyyRIN8qPnCAMXTHTh4drzRZ39Xjy3
T6Z2axbfsNbMi0KgPFgdhx9WRXC26YMn2DcDqfQ5Gk9EPDgTSATh4z313Pm07EjFC85n7Ke8rdV+
xkUDbj92x3GWhgshO/TJ8Y8WCTiv5eKRMCTYE9R8BAd+xqISQhRkN3M/J+CpowbNv/kiaR7DghYC
P34tnqhJhf/6zC7Kp3YRorTAZlKsTZ1xv5UyuDVsZdxgpsybbN7bU40SSG2hUsRcNhD5TBMfDqqO
wZNXQcTj2Q51dbuWu8G1bC1wevHElEkX4P+JzeNLaqrI5B2YyikTUeQ/TPHl78isKzAojgR1e/Uv
lkVITaOAmvjcRYmFWndXDIiXB9RV2vbDWLaSDtyHiioRqpn5rOlcrlzCmi74No39hAYfbDWAyYzt
17xlCUY92X/1hn8UDE1XGK8b1Q45/vgm9JUeUWY3HW+s+4MrlTLY8+fI/Tg/z6ZyzV4xOtg40DZb
kzbegdb9JYYVZ2Z9AgDa3GGCsnPm/5BS8KFb6nmRdQO1BfM3Rc68/dpZlP7DOFMPQt7kXDGjYDPm
jmfQiV0OiwvCEmluP/xLO3BF9TuqFS1cDfl73xU+r9ocXZaqakUHejjIVq0/4hveNWSqfgKCuN+G
ENxIgr9VNCRxD62WknTNIJNkq/OudOFG6sSi44iZ6aza1dQG9jpivk+AOEFHW0XndpWTrXFam24n
BPzpQROKfKg0HyCZwhpNmkV0V8ZLVVnmlllicQW+mh5USCprx0YAtiwvkzGxZ3O2ifsq1eLqhk+x
sHWQTUM7elCoQQvMDxPGa9kHiutud2uws9A3wyDPU8zsNdHSh/W+2NJgBQd0hfDW2KF8H6eanwfm
IY+Qfr9sjdIUWIH2RlM69wld/LGiR64LXzef0WfIhuQjBfm7bVdf1YVgWVniYqrP48IrWVcTdYUT
PXV8/r/zz0j8gOVN3t6Gc5aIG3ohCCo2avuz4CVZIRZzRrbD73o2pggMwj1ITq9zygKFd6rfygKb
Kr6Hc2mT1VDsGO2Ma6CTb5n69SIvuCkwfEUQnFVnE/pRqvekDO063O8Cx71LIlaSBRpXYN9sGMJz
uoeXlZyQwxHArfs+7XBBuQbCTWi8V2u2t98+z6X2sGuafODdgwkdV+F2GgCy8srEKCxbEthTAycy
fHfjfXfFb6k1ZhkTDO3QyWeYJS4kh86H3iV1lWJXX9f2nV7H/lbHaZgFef6FQZOaBiFyp0EsH8bl
9f4jrI1nRXizM1s+wVUt0KJz11BfHxJPKXmycAmraVjOThlzX1+Qbl2EnEHVVI6DO4is8ocoF47n
qeVaHZI8xgZe6OmE2dRR5Lkko2XogWA8ACdmNDlBrYCzZEoTMdEPQlvTIl1+2WpCki87LdRUb0dF
mnbCrdV7op7YqO8D5Yfpu2x7UYYIx9gahifRrkL5JDid64IaG9pSORLmTdx8XLS6AqvovNMJZwhl
SuInRABeG4F3LdFX3ww2cyIXekBtsVh5MK94IfwQ+5WbNuSBhnGsLk9UiOI/qEg+qjv7OSLNFKEx
tT9Lesap+lhhFLJMp5jchTyQ4J2SixfUQ50Wz3AxrMM420VoRWnFZHDahUHVJj9ilt+kyK2ebkWP
TsdaHrgOvBh2Ib+sqT/LOTi8Xi/ioeN1KR2G2mozEpw9SgqhuYVy6KEVXBB4YkjWGMIeiRGgmL0x
BpKVLwrfKxgoVd6WQwiwvTshWexNrRlJf/GmjZJ6cV34yZr9M+keWvrzgkKD2zHfp3NRMJec1FTM
t5CzIrEj07TAVJ6yApFTI06vRoIiiURcffOVV/9TPdV7r1nrJLrYUTIEOve3acw/yZoFUKCG50pq
9rotcxOAGayh47r0u8xal3XCJUwp4/Xcrt0R3RF1+z2j8eOatV3WKJougif72s5E4j5X//WQw5cu
uJbLhIQ3bLbQhwz855eOBD3RpeZU2cDwJjXPOSr1BZ85VeOG1zu1Rcs5duOE0GgPu9b+uSu4sh2t
pjwDh38A5kAAJMScexTNncx30FILGUM08DRQoHRsYolu9weq9TQQppROPPdkU46zCkO4oj9jpr1X
Lv17f9HLhjBy9V+gT6Aww9D5U9j/7MT5dkU8gEqmdLbJOKuHIMsqv8iWKnIjeqHWD1vHBJ1amoow
uycpI41gNz82z2CL5cdF6yhRegHPxI4S0qiGPSmGnSKG9pt5ifnwHiXj3Sovn061URe3CWFaH6rb
8XwcQtk4TxzdbdDEWrEqFHluWKR8wV2MWavoUV5Iouf38FC/pURDxtNI2IGnkL0XK3nuXYP26m2G
ysHSLiO/mVMpt91rquo5aslQxbMhN/fO2CIJPetDJ1JHfLrIqJ87zu9pOWmtecsSv+hX6OuM5GRw
VPOPEsUoBbkmaCcSPsVOsRubWfMh//ue8mmYXi+WDWk8ifd2Z5vv/ZCChMZ/fjC/K6jv4fj0dWpo
T/g+DXdsQQDvs++LJahgj24lTNSE8Eujh7BdJT3mGuv9rZ+nXpwoqMdmReK9TYsI+Kj36khlZ0aq
QC+rIF5m81EaG0FG4g3AHJFxqhBBPOeXkeY9ETOJh7nHUIisAzVu8ut5QhCzYKdNhsfK6mRxsTjC
kJUixHE3T+azJ5V35ufpYwpln3PbO8C8EplfXnkd+fm+ZC1GBXmebTuzZYkl5zsrb2cziq/eR0XC
D8COe2swkAHlIJwe9Tj9rUtVYg2PLgE/RT5+He7KeGDLiCdUONYs2F/Q717J2qH98cnz6AeG0L4P
Ohdm5QlIzmOYCMuohLzLLq8gaJmn8SAJsj6qMx5/YtfgtcpPy76ZV9e3bvU/ncoahli+2ejHRLEJ
EDE1O4kXjLcHqDk1cVoigji4aOGl7wj2NiTbWQ/WxL9yafOQRSrRONwIHSmXFbKVzXOvP9N4GFN9
LeKrTOK9vH6vhwZr+2t4id66CmW0xzqN32QzPuQ9rehbWJObtrwYRTHloxRVKoD2HYI5QkmtnjzO
MS3w4/ffLyHbc+ZEzUpQC+L6LddLa+V8pvjfsmABJsq/61YMbS6tqvIk+/lF7E540Ypd5bsEHc1K
hRLkg6s6J7Wbny3/FK6sw9YnzBbLTxMkCK+e4CHJgyc62v6s1NQiXC29W/C3qOvruQmGToAep2SI
Bn5gYiCxp2BeJGGbEtOm0TGWylaY/tiO3KsYnm4BLbh0Ql9IqYWPFn5TxsM+fVwjkuEyFue3jJ/f
6N8AC0ngJaciCYUars5MdqBIhK8EFvj5uA9MlRLtgU4cpt1NZ7VktsPhPTqPzxzR4TjM17Fzgi0V
v43BsRN4jiq6rErd0Igq3flPkONF18jHJsmLe25mlpgzCx2rnpPVtg1JbDJcsSe30+pYXRznXneM
iFXdAyuIfz2dpz6r8uQclxkcmMvRhrAbUWSYtEZwz2Gog+TU9uMDz1PgDf3auBJHbG1oXUITdZmB
jun3MDPUVekyJddC+el0TMZsOF8durv7dtNU3dcYSMt/tVW7ZbO7hiQIBxMt6D8DgTEiwpR4u6SB
Jxn/hKxidAop1FUtRQljwlxoj9FmO4YGRW9BhPZKnkXpQzgAyDOdpWl51k1jS0Gm84HejilTu4d6
RE9JwvM1t/RK/tvp/6Dk2xRSIOItn2Tt4DoQ+kKWke/dNoQYJey2cGN9gBIBe2KFg7d8V4o2ybhq
ssIq0wgh/UOnejDi0Qjs4L0meYf7oEe++D1tGeKl/PY1ycFlvW0Pm3DS8e2A5DiRnQHaF8t8lcEG
zptx5KQJ0EFOlgRU01CWcA49S03kW8Hi+mmSERIIXJBi50wkG9BGPcSo3jH/Vg5uYARaDMN/GqxD
urc9ZcNFDecbdZ3rk1DJmzrNZlzCfa0jI85z2splEFuGDStpdQSRp5nOCBYy+ZIqU7H4elDy5n42
hkWBFW2xV07e5KqP0Gtp50NryolyIgimE2QgLSGGzO5ESTpFp5sRsmS24BBgaJrEOYv0llT7zWUi
lNDUjm/geTe2e4yRVq6ULXyOXGQqHr9MeTDk455sJdux1SVhMvHny3dWy68hYpZkId/lANpNbxYv
RvnMfDbEgVlvl1oBUWDwAwDLm8L9bTEE6NJPVC6l/W5oDN0N8t7HWJyRcbBIlCdb172wmi00h8AW
QKhrWzJXKwQfPbTDGPn4J2O314zhy79FDH6GLVjJg/e3xc/7WC93djhDDOsJrK8xOWeAZ8NQzCSU
9R6PUz4B41V6SQOg+cr+HusR+O5R7+gBn2RJ0x090hWeFGmOmVq+7TltdPznqyHHBfwh4P5wMZsz
Pd51nDzCTowySo4vt61EdfIlaaTLyqSpljF/0kF815yKbdPPb7kBcUDJokKEWFEchOzjVCgSFwUP
u5WmZRcRHgDIebVZMZQ6K81TpkI41/B5kQ/2IYQTfuocy6NlXdVdGeamHEpEfk6wcw2F35n4cK4w
YFoAtZdThWdFa6/wp7qIUUQf20k5AkvplsFRtYCUgaORJIeDvESYMdxNDsyM2M/KxnW/r+zXY1GL
M/FyqCLBjoLlnFlvoY1kTame8kl6iax8e2oxmSJof8o5+t93p/EEGakwLwprWi15WUo3nFvKxSIG
OfwlA/X4lfHXhk3zib4+bmMVXDufF0x/1BP+UzX1aNlZ1jeJTelkv8rmZ0ZzToJv556ojI4trjcx
atcnVCK9CJQZoa/dfYIuIwU1q8UYxIxuqJectDTgqaJHE7UbT6eGSg0SF8rLArlVi0qylOKEWm/c
JUX+2UzJ6d9rs3rSdGzBSXeh4Ltg1aEIM/pQgCBIUJ1v+tem5j3Px2qSNys3k2Py003n89E47Qmk
U7mE1Tn+WFFNd/RN3Sb/O/kINUHYVbIvaGf3W68loUhnfSwdX+hYZb+owb9HUE0Jydh8bOJgfBA5
eELpiIJgAAi4LdjMiQ3aMgk9o/hyzjWT+XSrp71jXHTX5yJxR3JiM5/ADkeecYCxnf6yxDTmfWFU
YHvolhkBvitmRnJ9wN/J6ZJq/FcIp8HywsXPRAic1aJQ7FieSUiVjnSOM/DNumJIXtBR90D1eaWF
LJwXaT5Ou5ggGH0jVRkT+lz2xQBSshorawqJb/aN3hwvpRQDf93/7f72p2DkGHewFPdOIyBvP1Kv
SdBaUBQzHp1BEBOJvEOfxqqo1XiF1WgtJH1lh5fVQ+oXy9DnMOYOz1pYHcnwwqSAGEMsiSKLGt1O
rK1q3g+YtIPLk7PT83CbtlX0qQLTfL38anquZCtPr47abpwNF2pQ7Tf8a6lyFDikt7kWUy4xbXRa
QO6cwqnMu8KCkUWyUv8Lj3gTW8v321hoSHUXC3DwQAV+LlLCrT+PBhEJLYHtso7JNY08u+d2YLFH
O2g77w99jLuAoqbZlWBCBOwdmvW3MgRPidyo9m/40ui9k1Q+Up1qGDUwSFXEWglILJHX4s38EedY
yja8UsVNvPDQLgOdM8GULKK5f+1FkZ/sVVdQ4fI1/0Tx6yMYkH8KVa2dZhcN4Thpsf3fKDCFmQJm
m2E3YhDah1nw84qy05pZ/k8OAw9CtSdY9F1fOO4cALJQKfef9HMBlfz5ddq1G6O7eVbwx02j7WUA
lLvl6fuJDHjoxwxA5ZAP1B5lbd7IrZ2uKoEXOkuwRbISRtNeM9PzhURTXiGqV8Uwgkz9soFNkwVS
iIy3JOgVrE3eP1eZBQYULXhU0rS1gJ9Q6SYBZZRfTfUy7O8vzGtAAk25b7STd2SrfDunEwJye7El
yRlA5lVEzygOYa9KCrebDwja8QpD95HaDOhmQKJxD1H+tiPZKxmq0sVP2/3PG40u9xUxnAuD3Q5J
fHVCLLxewypn8EX/hN0Ctc7HWYRjSteBxaQglR/gu5ueFbMM3F5NaQTMoVFRFc8VkMmDu8EDS/tv
TtQ7jz90nyCl4kZ7S81bNtbGJiV4/eANhsZNeaINeyIHsXsZIeMS2/cUGFCX9iY0jpwPnTFrqLY+
3MKXcPN2vcm5k5IcRT2FkwDE5dhahCs5rvn90bYJqV+iprFmzGDWZKe94gHqaSWigIPW+kI/EhDV
2wxdVD49rXUpJ2flBQfz6hMxO8ZS2qcGNqf6zjwOFJ2YuFiUEV2zFNd9Prqp2AnP2hcZ6RxFKgWI
vS+780bmGiDPpI6g5QO8b8KY4n9RnIdav7YJz33ImcTldCy+IooFIP5q7P3mzO/yDyCvgV1berwz
97YgMjGOGhxiFGUxK4miurKzpxdqIK9s3Z1WiJK7M7BWwOWigGnfAFlgm9vqL58yp8Fn2cSKp1NB
Dziwhrity3jpLtH5Uy1sENBqtNIuH7Hww/wrirmHPLz3IB2PbtRJgDmqZ7aeqXuG4W0/QQ7iU27q
QNbpR9E+JkACyCqeoYNVponwstyROhSwOdaUmfiLd+uCiQ7MNe48nkRSlRYceajicRHK2GzpcdjJ
n0dZ+kDsFMamJqiJfWdfMFUFmhE8IzrFzcVXchYnVeLm9Wx06mpijnyRBMBJ9qVj6xvch3Q7Orvb
7CnxFR010wFHd+5eX13yv/FzhMMvFAlHIzQ/D0KXKZqVfoqqrmBaGMhRm6G+MvMz9TEVr6dELk7r
1hV/vrpfLXzC6btP8XdGyDu65zyQDpUMa8RiE5xok4D/MIkgDC5ROZSjzsHryiknkXWDJW5DEVIP
fccQs+nyqUKql3GIJ8w6YS5bdcFKJV2YLlwrNv4EqppF5L/ZgHT0Ga0CUy2LeiNiy+f6HmZazzUu
Ooe8CUGfsVfvYM7kEqA5EY55hCpaH+CSvuCD+oSC8rSu7VzZ+QtsM5av6P6CJb0mMAlefGIfnsYp
Y21y+APEEF191wEPd7Q5ABK4v5SBXM8Za5dZCyfp503h4ezzWFBnfjxeX5scomtv7szljTaFSVeO
N+/2vWumE65M/GcpjepJJmmBvbSqd8DDug7h7ne7/dCEj1BrtFKnEwy8WSSUjAWZPPUhcjXMl85A
wyDA7J7mcwD9Qa2ANGdTjsPkrJwg2jQPPwz7sq411rhTBo93p3dGnU5HT4VXYsp6O5YciMP+G1fp
fkXIpOT/GdHTceAD807QnFNvAEakZQzGrf+9iTeGtqCwSmfqSk4KWehMC/wQXJJ3G0jqQ2ZIf79t
ZYpar60yU1jBqBKDMGS1dNuEPmDLhwndOsnNnkYleg6j80CGO5LwjUbGOt0jC8ts0uKpCHw8VyCg
nt3SSxvU+Dw75wRFQrZ6cc2miwseb7W3m/4R5hq/QU4FN3NjysORPggBhq4W5XRbWxzUkpMdnf0M
WyDU05LussfF0pr9uCTFlOsBSp7NOU2/y3tAkG6hRUEgMljl3CoUsZEfVRdixrgFB83/CV5C19FP
zNn/J9nxUfXsb1AZwJcRkf+f75lsRy4ajfkIAQAyY2J5YPmzvNxp42DTot/4B6r5rq7FOcaJ6oKs
dDMA7tgcF+F6HNTbdqJaCxz80/RLprYyeLiSXHweBClX40DVWzuCBSl8EtCbi0v7qPTWpOHEio6Q
ZfNKg/I6/01Wjt92QeHVF8tG93VrrXKEa41NRhEf2iWQvKz41BTu3HY74zapOSkxNas+emYuEFSb
6gqGiEt+teM99uClmlYs6lfbXMJAzDCfUL3IhxEAvrlDJ465mPHmGh8xLYtmHuZ3NSitzg6QgoH/
/wWr98y9PcZUHiT3DnymmyXp5Tvm4jgNu7t58/iNWuikdujnmNE61abUVXOAEYcgSlHg+RYSf8CY
nXiRbLUG2HjC8P2/i9MLvaK0gKZreOSt3NRKiNVjU2Bw0dZpDKoMLglylNPSO1ulGMkDR2XxCBYy
ADmj1vXotunHMeDVvpZb0/X4roofW7hkIZTRu1yGWoeZCmAx/wUd0wOyosXugtaoz5Ko49yFkod/
myUTsqIKr27wtw6hvleLcNe6UXh4ue5E8JP0Ati+zq7CSF7nAK4zkAVFe4mS40CJu3fsKQ793q0T
s+dDrb+wR+ptN2uexs+jDeC6R0PQ6P0vYidvDkRzDGgBcojqN6qHtACFCtwTk0pqfGs+V0O/NznX
0aYKNxo00mIBEL/gdSlhSpkv4b7e5DK4Urb2/4c+jgs1iQKzEKFSk45keXkXzybHrGv4msFp9gF1
aQL26S/EE3DlpttxVRQrMqs0s/1a7w6z86kH5vy8gKAZy8R5gXbfe0OlvQ0zfArvHchvpnb1wXe7
lIw4nEyd3aNrK9Tr8EVasPi44PQr9JF71e4Gk027YoK/UQBXxqOAnfcWSBQOoy2FpTn605oWQ5GM
Gd1lFSkr3EEVDWgrs/qDZsGbxJEUsgBHNv1YG8FEcueoQzg7uJysHRkShZiXYvsBBD1aTeicJDJF
nA4SHdjn31SlEjOvC7iWRzOtEki1F/FnSchhSwmHcHpWoPG2/Vi4OnDaGlNwDI5FwT+22pwIE2jp
i6p5ErgtfTkGzH/Ox2//UEsubEKQrc3lAG3IkHIgsv5c/lpppt0sVN14nqWhNBx2aFibxkVuDOaB
oqcFHf2hWcRq/CpF7tJkPF2/+f9D70DlJdgvEi3VzyoRCRsmukYbrH1mZTTWW+PdGkkmD4ZQio6F
eUn1kLGkx40kIstEciB6WNXeWJ2UmnfWR0+Hm81khhnj7Nhw1kDRFRMityhBqt4EWQNBYcIs+C+R
8AI+2BMk/VR7XzPBcE5ttiGb5s3oFT9BtGytotsrf7Th7XJbmVcnrJCDKPCeHlFUEYshmLMR3/zY
rk43hj36R6rXMz4G0yG0KkPLndmgsrfZv3qOMnenF6XeBh+AySIq0QwL4s3lHASqNXoPgDWPE6Or
bbRFagd6yRdoBjsokwWpxgbd0+2smP2o8XI1XPCv/hggV/UiUiRgeKo0vZYyFfcK7GD4U4/pCJBw
BcSwYDHLbXSaGmkcsa1w1NlpOwMpu+/HhBCyHxfJ9oUwksdDvArGaDSgYrIOwDNwn0wo3YA22WkU
OZkMkSZosDM0o3YWP1WWHPszbM7QSuy8axu3Sbr5fFvA+h47vcm/V3Bwt4qSQCozj5ozf5wVBwBs
7NUOy7fU1tMVLWiGU3VdtuXUndc9d6xYFXqyMtIepVKHT3EjrRiITmYKDjbPeRlHVuFJBgwXEuoU
scT2sSg/sILpRN9PUvpm/MP/YCc06LyCkKRrX9VH4VmpfKIIQ+ERTbslRLOQyJQns4RXt97cf28J
PAZaxBk5bjMxA9G/nvj2RlJ3BmuKtg7I9RBh8brOCQJ9tcq+9wMhQEjQGlxzga97F8pyeFgE+bbw
WwMTX49BIi/DpJ0P0kKXgs8KWAvGsohyrYL5EfrKFh1eQK5vvutMs6hcGDoEQMxKU3kGFSJ2M1WP
iC3xa/ydGYj+qhFPmTLHZeuH4NkqJi0rAkK6gouqJprNQTiyTxv1i+FPvA8VgEV1UdoTBh1BGgCD
yumG1zn4KOArdoI4arl72fXTyHPyPQt75FxUr5IrSPKZ5SycD5+EemoN79/av2HtoIhHsEOgr1hB
6PTC2cakq9niVrRYBhIIziPGY7T3nW3ZHgL4hbNBFvtJ6S/tYgjxWi3vuTgCNfr5ncRRQpiy3ZtO
GCH8Ssvs7ipfvp9Uh75M/0hGiODGFYDndFfIqRYMLroIKAAW35i+JwQ2oKe7GXwdKYmaAa2Cj4Md
0i5klVqUu/uA9zVBed7YY/xpinVzY2k/5kQac437sEY+aNNUXuZp5KFPhM2TuL/SjVl/MK9huVt1
QcGG6qhltx0HxlEHoLFBNCvv07UF/2cHQAXFp+bYO2SoT1H0DQmTLOqPpIJ0h9tORKngIgH+ttM0
7NuTVKTO7MNakeJIwRuqHe6b2VAe41wTx73fHZ0s3SZT43BNWeJ2rDnBwfopmfoOsIS/apQ92TxM
smFZDZlp42qUp0yjBvKtXRByRiOG+x5wdUZMOnIwv6CW61NlUlaV5q0L7JX+kT1gxce7kybcrNJQ
3SrU4lEpqe1RHh5eGACzuEihopbxpKrdut+I6liJxhTzg/LmDZSdN3PSiUP1zavIW4eNS+Db6dM9
+0yb0c+/hSYnbKmwXBD9TgZjTID8Fli3E+e+Suw+FLRVgWbhTQ4rJFlZmYQZmGpAcQ0R6Zjbp1Ss
WSFtTS9PVwYdN9ysANqeuFtAHwlUU9bG8Mq/gzEBJ2B/7JYCgNZnXE0FJszjZdQBtc5y6jHzQ8s3
CWH3OHlEKjKebOd2tgUfK/vHC+h6WAXxQ+lCVOZhkwZHKEW7ezmbigAssuTLbeL0yKtfdVzX7aUb
HYAXBFik+L/T/AnfEaCdcSLs8foScaAMTwEaM7qp7kE6eqaMHax6R/s8mWYnLO/okhK5OjlHGUX2
3EzZoFq50TUJnb/Fg4tXhZ4Goywtzt7IAnV7YPzXFmbZF0PvgLjeIlVsKjohT1gYK4iMeD2O4JWC
8wQBUrflUiZRhew0JAPwcAo6AukOM6y5IJSLR7clTlcYQQ2dSyJkeQ1QDaGcAQW0/zSpphQ+yQyv
ah0LvlE/AN8Fxz62Ks8ss2PYDnPBctTEgvLx18paMHeHHv7Lp7/5qmhvZBQaC7nE86Gy44O6R/AX
/a6rQqfCWnrDO9sLjdct3PR2HvmT6mGP9y7rGnkXKHAPh1aIK3qcYRSYxpKoHQkJpDA0rm90pgNa
SreeovWl6U0JBIpknSHrDb1cCKinvN5TCaYbBVmez1GDnSuKVn3xqyM3cVSjwqsJ5JbJ4NKJqQS7
/szfL/TFtA9OJYEwzDS7p91dluizrKG0SQGqfYrp9M1NY81zX72mx9gHMu6J+k7uiZcv0+8AYcjB
0wH72u2TdbsHm0HhhZsyExvjKm/hMxZvFXzXEylR+P07dxua2aKqhtlhH/tt8PuG34TPQlBQjGp/
EJ/kf+FyCLgdpZR4o9bOoyhmUkdSMryLQ62r8pIxuf/NJdSnaak3rwTpQjj/iP5uy60D/EWrk/+p
2ijF1ikizTikOTPxu+8f6xzkavFQ0H6ZW/tnvl5cNIe/kbaCXqcBF1oLWCdJq1/l71YzyGsRvnf+
w0aCp7/Y9yUkyfPFI/V4M36w6C3WfulwQUpbJ6CgymFaPPfxBhO7R5g855Oz06/vn7mRp/YdvStN
vKRws0F1k/qdFX5F1bJ0TQae43BJDVn7Y9ch9UdUGPNdeaEuZcGjaDrmn6ws+MAgSGseQA3wF+c1
ip3kVASdUN9doKjQs3W9ouOgTsdMKJKdJKfA78p+tWKefy8yPH48q1bGr+wwFjcOKwUtlMpTZrG4
ghWwuvwoPB48xtMM7NHeQRvxjPbSwH3r8uXaMjgnM+Ybj02mt7LaHhX9IRTlv7uKVW3eARZrLyZq
gOm+xwS3ZvNk/I6a1f/mSkTXQ4OO4Z4gQNvhVVlSxNfdhq4LRctZIMQU9rPJ09N5BU52fhTm5jAM
VoEoX9mAAxBTPY0Sw6y1L170d/RJ95bIgpu+FhaCAJ5C3hVKITBbQlw+Dv1+kilWpynh85m/U2WH
VcaBn7x1ZNvY0C/n9Zaps9a4l+wlq/eY5067iWdQcpzvSUtuEGCecCois2HlyiPo+R4VY276+hhy
VLFqIVDvEICPRB2FBWzyqqPgweKUgtZ+xLHSzfDfcm3h/qrMPZoGzjoeY7Xh/T+YpiBTqLjQvIxZ
r/vkQFyiLvVkuJoKk6y1kzWE099Z6I1vOJdfB/GC/oVh2HlDnmJcGXgF/DHdQtXltU5AtOGZJZR0
JGD4ylptRctyWQ0DMUS0meCmLNQWNIanB6gPisQ4VWdpbpFmn2ExvEvuLatGnlAUIWw8QtuN/C5v
yYn6T5SpFTqH1j7ncSrFwmwcTX7syRcKHlfTkzCeArqYnkdGMY0RGEF0srO6HALYvU7fJIXEFvlH
fn5acpWyIBuyr6chnbUjqIAHVLXtwr6heObqw7DXfZyzht9OV8IuYxTvceSNhP6g1pL2snQZSr4J
hMWC6y0syZDCt1Nb8P8fYy94Tc93EE+iko0Te1QNKg9sBZVwO7XlxOTnkFQmSLHx/eCHKEWw9aro
PCIzFcrYFu2eAuMacpWRiAt5n7mbXTy6gOnlJG7ynLI5XG8X7AWNQ+H8BwbU6ORith9FBE9phrKv
+xA+tqEOWOpQQoouTIOHec7AMd7vkiHZY6bh54IdrlWRRgYFXSh7jGkvxNrdVIejlyDBbi9lljZ5
yp2UkFJKPQkxhpvYyPLoV97EEXosZ7CXTw2P1SfkJPtSTeCQG9nMzrKzxlktZ9Qf7bhNoBGa2QvA
LV6dZJ+EFU2ahOeESkWh32RLWCPhNEwA/QBwmawUWWaEZdpJUL2VxkoeC8y9TnNFUc68DMLsL6cM
Rhy5w4Z1yJmIYA8kZBH3Wzmg2qMZB7Gn/JmYh8cChu5OslO3lpu1B2x91TBDHatxdseSJusPr8fy
zaBP+7B+rgMhW21ZrptVFLqJFNJuGSTHCF0yKcA/ZIcm6V+PJ2ueyFCtxh/AJb5oYoXYbuFAA2hw
c4XLfVdsrr1ddOcVOS6o3HWm7UwNZWIat7oKljtyJf+JTM04KJrcznDX0Oq9YgEJWTl11sh99XHG
0DG7W7c3lnVVZatNFR/MbuXfXfwpzdpgL83JuWUV+k4Fto77Jf3fmTJ64GKUlJUsDGjaDrLOcr6A
5J4mA+C5m3JJ5GpCzxTLO/RW2FW+YQMxYcFBQ3c5T1ReBqXx/HfOEgDJap4ht1QWiy1iPyCzZuQH
he0vMxohfBXlug1QGOl8F7FvFTktzvRf38MXJZaO2mrmooE3IUeT9oUMYlrABpIzmozL29CGpGzy
CA5FY9mwwo2KtRp1uFi9ImExo0DUbw4PUDB/a43q0EPPa/ls2PXRvneMbRP2qbymizTSbeiM+2H3
1Z+DTmAdcIiOXQd0B4Hw0onbruewp2Bz3q/ms0AC3hX15q48IFnAmvVv02/pEXB9Ifitzt9zTW6f
Nwy5OTsf1mtI+vn7+sm+DoPnfQ62cML31g9X6dg8FAaVm0OSqcFD8x5wdvibRtRHcpXFKTmpBYdy
EX9eWswlimgTtvaRviBY6usgLeRTWon/5HqbyHgMnWUfjPh+kH+JZ7wL7eOfyeFa5Sk59VdP9dqk
U4Ia1a7cJl//t9JgHkkZBY02jQ2xSYqTXaHO0Ejdmuk+flZfeG6zLnos5KTvbknH6vZgUuD8vlu+
IRY1FBTySGz708mOdt1inma/PPhuka8xiO55vujpzj/6cHFMMweTopZhLr1KmPmPF0+Cxlii4/+O
+Ju4AjDiWJwEcgOdUT0C5v7aMLc8LHkRYzv16UE7tKA128hRi2HS/ZqDVIwyMZxJSlqbsdPV5kum
1NIpXBptZVcXo6TKkB5JPQHnsjLv7nE4ynuxPJGeiNKpx1G3QPsuTeluY55Qd0OJtGyQ6TphrZUr
uH5e/nYZiQ6IU+DwT1y5pzv4MeyKfO4u7rsvVtrn+evHY5CVW5SBAY0y8zNa9GWd5b79Uu54yfr1
QFQqJvpa0e7GtQU7sxcvtElJi311sbUedbDs1irkAJEkou01b2gjBtwS7AYks6yo4/eWGTdd1BwD
PB3w698+0fnfUqZyrtlemJhOrTi2v6Vn/UUN9fnW8IVZXz3F6Q+PVfHOn9Jy6Ybv+xMrT5x7VGNe
AhYlmXxAW3ZFtBQKpmiooliqkxwiNuKPkTlyuRXQCSyMuXGLyz5B95ATISCmMLIzQiATAUhVwiGe
WvI6nHTeuRI+yVkkQwF+/Vzy0TYxX/WOTbsp6CAiF6MtmzC+w+UWpYk2DkokI1NxN2VacCj3fCui
HRCLjagIGGdyKwylH8KFyxr62eEf7QKWGw6K+WVJD3VTkSfgbTGte2X0c+L+/ppMegNK7V+4N2RQ
gzcEZS7TOOwchbzwGmmeq+ct8JBGCIXTnv5IxU3z2GGAY0/DmRE0G87aZxlol6LP3pZcVRNvWZ8s
X1JdWgREfo3sWf5FGZq4jWDTUTyofgti5ebm2JmdXrPz1KU5SoVtmEYtiuACWr40+JeB0AbyakI2
wM3UZxVtXbuwev4wgQbRSWyDK7PbdbQcHPCgZSrjC43T586EoJi4kLbMTc2D8uLSQ1W1rOZSCnYl
gHGwce/87W+bv9mQG+5KB4XrCzaUNdCVcxDMSJh7Mhrwv/jkjGNIhjFjDtm6GQDfQIAilAk3dhHc
S7a9ISDiIq/URM+kANBWG5Qrg6gieqAMGGby6k0ACuDsWPWxHYqAMu4Nh8RfzUP53tdNfKa8HzUG
nAb3cw6J4WG62Zmg3U+0PG4ZI5YEJUScXc6nE3oT4L2gv82x6QcLRroTqga9PU2J7C6ZxeSBrRfY
Pc2y4kgF0kP40hzyLAiV+JO6wCf5+QEABXyBs5KVvgbALWb3kjuefKs37fSxeAIfXGH7RBvrw/kx
i8S/QvF9tgJXVEFYgY2z2n+UbyfFFTSnZ4/viJuKJSz3UzrkzqyD9gsbW1+DcXZFbJW3JoZJxnVl
gDMktuygC1PjKxjxe8hdRkh6Z7qv8hW2vhSYoLZ0q5AS1thuEQhc7ADA4f2oZomQHf+h+pHiepH+
7MfnlW1QxDZwkE+ZpUDKXndoFIpDRrQ2p52a0ErQB3SoNkQz1E3RP5CzOV8udHxyufqSm14YP94u
RJC8R9/mXFJRRgt3KCnhkDgc6xCHrXssZc/Jq4Mp80L2ayiOeuko52+G4phUNN7px01+3VjQAHxQ
EpwbFx501Ea+zAeRNPqL9rg9gvfzNdSKkx+be43W9Nus34smRmyjuZ4DnpjzQUui0niCeJ93ogkh
5ocztrqSA0pPJ3K2PlEYIKuJBSWTEtZOFavoxR2nf7O7AMk34XYiQcv5JQmNNsV2AO8iG9KD1alg
reTym3L/yaLR7nvowCD2W9xszM1z3NsTE6JV8jcVuQ3Y7HhS/BCovSZsanXaWRAIyCqcGIxe/Kr6
1BUan624ksy//CRabO83XjcvEyGcKy7j2hgNfykFiJFcsSTqZbEhBBh2U7N9w2bCIsY7VjMTO2L6
QgwFcUqGQ0v0MjqYqLkKe0LKQYxEprgqkR0xE2VQsD/QbsV3+MA66K2TUTEgPhqa7E3nDot4ymlp
QlPOiPdFUnoAfGdHSLLVgL6p9Pf/60RdcNaTPpEU4PbtTnQnvsKfIUFgBiB1cIykPmV9sp6S/K4Q
jMvg5/xjgo5IqGYP3qEiLGSRwlMp6cp2OcdAZa89fTy2jxaxdPVbwiBlRucKnqTxMG6xSsazEnq+
9mjKOlfxUbrTL413m3AvEABnc09IxbT203dXgqWzwcZOx8bFMqn6ib91SVvId3U5RlnsLEpqB4UZ
8jQm/ow0geeymn3LrhVxG1BQd+ciJI0CM9zhMCA8CgZHNkIQ420sC3t3Z3UZhnp3j1vElWhFKgbq
1UPQXYP1DpmavZkKDs8uka2xkIM+8L0IMAqftr6uy2jcbVd6Rqo8u0sCY9tLw2PDXv+hknA6498u
dhbGWh6gPlJwjQqr1JFpSDRY358HmNacpcR/YF8Kj7ZVqrxd4lc+763AlJaZOceoIUUeVj2lLPNJ
Ur6VIHFl/lSLxoxYFyRm0FHnUG+tAz+lhenWN/WWo7ijRpEenTm5Kf3T7kFSIKGai3QllAhd8nnc
30ybuiHCTsBequQugLknuJxGfXhJ0clg8u7tjm+axs04oXJ/yA9Rf31A7ypQYJ+1FFLom5URs57d
t2wWZU7/o9Y0qot+isCPzD5BomGslm+HuCfYvu92OzwtPHH7J88gpebNAeYDYUW9TZ0EZMwU8Aej
XESLj7LPtcLFr0+B2sfNsd7c2yC5SNll0Q8srWQyZqzFsl/B/7YbZ11NK2cxHrOe6cJgokyRnNX3
s3wvGMMdPK2aeskywydhjg+nwm0sMrrvX3aYdBtTT/rExTgiiMPQJgSuQLp7AwzEir7/Crmim87P
aEb0X4gjGACIpEEiVAs1HSlIF+y57DjR/SEwWefRk0+sYr5bK9etFWC7XsFJyilxb2xkE7tH91d1
IEPgW/+WqRL5M15XrfET/FxXJkEj+FKmhK3F9JXELoVvIE9KiqGVexNEJJ3tM1BALKvHItQySzJn
nRsUjDzJVQP66GBZkLvQmcxu+PAlcgzhI3X3cUfWsxdWklDYjpJjAroI8SAMEtsdlo8BYLD+PnPv
bg9l8YTYEMpAEFHDNB1/vOXdwQzqVdfYzHhfJBCf1iFF2eTKALTmlZnlZtweZMa0PlqH2Jydd5vs
urpXC0GTZIS90rOuf4EIabuNbOmOmEfapkfdOpDaUOoW0cYAx95qsCS0+8q4ZoLa+2QOJxtmQv0O
Yj0kSc5glBSEd8FyB3lkt2RGFD3Vjwj57/KbzL1bNf7rBprH4Ps/lF7PrBSNOmsZiO6MUzMCLig0
/yKQok3aRqGThc3l/usFtmb/vp2seZeoL4WlL/M5M96CCKRu3hsz1OBcwEZzldzqLJszHU61oUDI
0ak75kGTgLVBm1l0X17dmNp4LMP4p3rlYHjyritykeDuaCbgBXgGTVHccJU+gSfDJMZ1q2wxOomE
NjJJZqFn256eGwbht9kN8ap8g42kRPj8kXbet8YdftLVGXYn55qksFodKagpUo+zF+dipK8fdu6X
u4WBBIaPglDmx45fjETyD7xMfy2ZqMtAPybIG0jNGnayHCOfT6fddeGwYh7cM8bymcx5cBxQiFOZ
7AaqQbzE0KMXAVOLVLdme4mQtqiPbBpdYMhSOf+EkEOjfmd0D58AFau8HwSNo0/dGnP3MxbSBCo3
eHDOjRpgY3TOt8Qt2Qmvek3OoW44lnkWs3MkMtBseY6p4OAGTlQKKBoK/3/XNjdsAusmLQkVFp6k
t1tStuHIW4Whuak+39wmX5WJKQu+kWckU1ooH2WWlP3WfA6AqAWOjvc3+F8bEyrtE5IXdtZGa2ub
3BTgbTA1J/M/Cu9g4Gu7M4Lx42RXoc4NHDPxitsozq8UAWKx/b+XTeYRWBylEaTQ9yRJFaIqki1w
qRW/1M+glJaa0lHYHVsi6kJxc+Ae4n60g2FkTry2VP3Fi76I5mrVDC5Hd5i3NMkGMpl8I1LEZQiw
w2aQb9XJljgQQvKtUD3sd4nrGPQL7VTB1pNq7GdKnfNUuggHV2VtKWmCzTlD53n2eQYRgsZOg2m8
68e0wysIsDSNyF4C+6CdTQlNNK6p5eIhpXfRH0SazLsNAj2Ms6rTFMV7pEe9Gqri8l8e7TY06L3p
QIWBQbWbqxIVmB6AdfWeL9LpqcU356OcyBQZYfFNBRxTZnbhwFiH3pQrnPNUn/Hy+w6R8X1OFpVq
uizknf9KHpUqtO/cWpacQgwljfG0K2T7ERlElfP/cvbCRqvcHGjC/MIjM4WvMJyrEpsDp3DFmAFG
C0QJflfTHfFRz4tTD3O/duLLReq5NjBZXLztimkR48NfWQ732UEFOdxgu0PfWUGszLv3YWzhuLCr
i/PGJNBORFsULmr1N6NLg/i/tcVnYOh+ljC3OilitOJNIJLBXpy6tv8i+KR6SHRPwMu+uRE+uAo+
yCCunpCOQ4KqgkvVPeUNlVQXg9aKSdvOUJRaH0hiPIWGl1HU9wmhYUv8u7O8e/kFneudN3DvvmGu
+QoHpGZXBUlyhaaZ4P2yekwpOjtFIJ0xe8+qaZQaO3rMnB7DfxV+WBd5Ie35EATRvYwHeOCtSjRF
T87Ymloctzc2ZKOxuH4HvQpdSIt/M59FKUUvNZWuc6jK/sbs/r237gHVqkhAWLpKq3svc8WM1sMh
ZNqS6l9lRYTi/iL8OhC8SkF4ewSenb0HYXmtQEy0DIvrNT/RPsysrdSBfFRi+IFrSePmCrLgxejh
uNW/VuH3PC1UGREciYDk5splIjXVExzneFyrUfuvzr3ZiCMSjQtKKKgM6GBYRuP7oL+05A4QXEw/
VyDMKTx1o2J2vQKAxZ6QVBabTga8RIVZ3GlnbydOow3/Vfnl3iLKNJKgBc7lCP7H6cxwGqJMDLe7
FmrJ1h0XCI/u/bPk8ovU9AfdihRFbhnHwbik3fFewfe03VywUQNxp3y9TUWtiujyTg8egB9HjlfE
lIXPkkC72MOSP7XyiEJybeA/aLBDFxbp1X3sOXOgy84SKKzZxpH8w3k1lZIxTx2x+qr7qux7DKlF
YRHQ8OJ4kTHEgV/Hw73SjI8kzI3h0PUlmxVQJLJeACa6xTxbq6RjrZz9+JyeMfTLyzN7i2dSOZoJ
0V0qycCgVJtJdgmHrw9qv9LMtcm27uJIXGFGMssEHt+Dl33Xg5YOTB4J3DVXMUZOcQzpvrpLjziB
fh1te08Xsk/iCSv5RC4PDbvNZrJ8C2L6522WS/mJ1jpoHHNGYxsMsba5kx/A/428FW8ZTjutrzjc
Jj4FuB56zVgg9+DXxdcX+AK0TrqCczkeEOv7Pq23DapdQlcuX6/uLIXf20JFmXjnAXVDP0dITTLb
ac9R8UjgYf+cEHKlY9osO8lb1JgDZ1jpfqncgB6RIcTum6w3Qlyic6FioH4JKKLZATAI1FAzfs6W
E2f0ppYI2CBgwq4cc+HF2YhzaEdd+vEKBgjOgUoh6PCLNf4YE1lW3j53aX9bwyLg9Cby1B8Z81jI
uCTFEFVVhZy30BnBr1LaxmXfgjzAJmzJRbupzmoiV9AlyDy1+PEZDWi1tuyXoch9nESBJrYdpj4M
9Yism3tXCdyuGekVOdfP/AXH0jAlQ27sWQbsu8BfBW8276BDSWmtJ4HADdV0U8GurBRgnYFjvIBA
c4iGvOIZQZFI6+XsRnK5AUVMbCEWemTzjnye6rBASddjre8XhFfA+w8bxldSnSR5Rq+DIyQilWF0
WHTRYzKSaz7SvlX0NukjUlZsvAvfhVhKezlt1jNgqOGqBcEXjn0ML4sdCxp8t3Q7BMrq1EhdF/qE
mRKSHTddEkYzxwPazj2EmCh2X22doxDZI6f2gx+TlbTI2KKEJ3SLyyFNyGwbAotwNRL5CEmjCd8k
Wq9UZLobGlw93nZZWzql9FIIZemjA7ptGgz5mz6TL2rQ8iAR3Bzy+pK97bvBo2yBiPNKimyLJ/zO
A5aygmL3M+QcwfbHr3gTXK1HQ3VmjPmhKTlFGD3OayI3AbiPvH6krvgOGP2jM5DO0i+MBaE09aw+
Jrz08BEWDD29Crpi+HAIv4oA5pj+j2KoWTYlbyW+x0vvixY9tgXAYlPzHuc2Ql3glO0oN09fF94G
/+dxXmdZPGYw6Gc2pu1kOd/KwDdObNvXStaYRnoPegAnuLHRq8MygIuQ64nIvSHodQ8i7UfuQ4ek
x5WaPAA4yemkuNf2xD9JgjTPmEq6k+il+ZALomt/ubvxZ4nQIWfNYmSEzAzSiFnsf2XvhkWnWSml
CcrUhG5/qTp2bLBJxZMIW8oh1bBrpPxJkzuVMcQ6VEBKEnJV6lMK20CcR1gNQna0mxzxowIajRmW
JvKAFF5cx5Rz6ENsWTl/7gIpLlhW4/rH9GyOduIcijz/vUCIVDcQCyzYL/2aN+3olXImrZfSVDs0
hhIdvqCacrXaY2aTqrFb7ewB6qegMQqVe79dw4CFW8nuAedgglGVoxzL5gVp/1JEwcUzLDVQXWCt
QfIEieIpBVKCUSc+v+9Gtl4LuQp6taqHEQPrgz09+mvmuH7WhDSd0uUOx6W9jUE0/k8ZkOit8aWm
rM9VL1w7W5qP56WdkqoNQksTVDLFTYLUnYm5J6XH2REG8EvpNvt0ct9kLIaLdDZVhfiJ/gUhtOMy
AZvuTb+j4kItm0WOJ+66+Ix2yFJxWxq4+g/Bs13kH0JBWytqR6nrgQMuLGcveZFp8gyjXIeaQXNJ
zYVK8d16UtoJM7k10svdKPofpKSufsq5zs7o7G7MwQ0IQfBT05KeNm2OJHq8fqpgnExOZkDEaHos
YtChBVjeuenX+Gwr4hxsnRqiIR58I6h+Xklm/7ipdcTNvihULx+RB4+3HXRazbVS69revRgjbyVq
So8U1AsTKBSmribaDaZjWBbvrlT26ZDwI71L8FX2my8Do6KZ82b23gGWA1SAwnVtyfitX9TbBRw+
Iza6JCcqf0+MF+KRtFjn/Y7lzUeUlx3W/iFFyaNQQ9WR9jwaeV1iE5EwUExwDb10krn6C70KKoWF
S8iTx9fphHkVpz3Cyc+hHucDfVzYyrJlK1B1bzj0fXdKdzDkQwgRlBORbb/7n4hW4nm8gHy9xacJ
UMcLDau32aj1GXoUrOZAoj0e36tKAiegcHZ4gAbM3cvQeo76btxurv+BXi7I89iOA17TmeN77/ev
JvVai7UDLoaIn+lyPw8+khIMCa6w9X9NRGsvMGckCwUd+6ux03JfyHV9vlsS3GNs9AodL8p7tvlS
4joY7UFwyWQXK8Jv9LG0WX6AdwmSig25mT25BqntqcPUtZkip9yu6lUKnNGDhliOLTwHa2KquyU9
VK+QFGre8reg5nbVQytmBQPETj9tGCnqB9Yt2qOjeew9uNcDyXGyqYTrqkiPd1kKk4Zn2My92WAx
1t+atmAF0g9lfNeLfwEZOuezzJ8zxrCaydLmJgIIYuoNKOiOusbsK8ngS4YFe8u31DJiPq8teSsq
CbMiZo74rWzFUIfaZNsduyh5A3/0ZJfvRyckNgzJNVs+u1ObcOUcIDYwHW8y98rqlYtygNmHFMr2
P4qdxwIlQO3UqenqmxAA9At9Ks0x+A6t4e3xOEraE2YQDhYONRfxI3FOyK50SVMvhix9GlgRJnoY
ocW5x8G+4psr5dAWbM3XyOMMz+GgJ7sd6UsGGK+GyMtaV1REwtV7tcVbx9rt+2vUZJtvmYvRrC8x
lAwh2SX2eWgod7IybdBOaW6oc1uNdHg3lHW5ydQvLZSX1hnV6NBrMqDxKgIfUQ0TjYY8H5MKhhCt
WWpojZ4pxjmSIMC941vnJEIzm9FYtLHZAGjdx90mKjeo2O2Qxt71SfkfK02CKoVgVpCii2AQP+ug
cmxFYNMlNc7T3ZV9pq379CkCfIfHI6DG6uzp8B6p2DUvty1f55HNbXmYhc1gSA0DdYpEoxXiZs4o
pyakXJh2N8T4HjL1kc5wTqWEqTj1JUaLgVeY/oJE2usZ5q/WuqTupJ8PJifpLO1V6lKHTVhZ50oY
+lzvr1bA5Ylp6LegVaDfv8cSyluUvYnnHWUaASfu1ID/JcSygtxDZSVmRoK+dIQ8tPGKYFTQG+As
uHLiPEEWhw9KkPdye1tsfjCsDCskpM7zAcPh+Bowi+ZHdU9VBH++42LV34muq2odFJ7Zp3gLxRCT
u/AENCCzLuUpeLVuwXzs9w2sRdDXSw1X8QAf/VuG8/Ygm/9y9For1ntliJGS42YV+CZCaY+ZaFY7
gTAvhhUJxofj5nW/cinG7+WG82NbSEBgmcu4d/zFmG1kFSgs4QRWflbRj0NFDn9JrNRgpPwUnd2r
QMcjloO/7DCoCLeatPSqX5lGa/H5/XUHOKzdQSeutI+PnD4eLb2V+cC1rtcRb/s9yQAYyuLtQ5gk
UAgFl3OcuvsK8ZEC8Zu3zlzZUx9llu3zDyH34zQPoZAVxSs0tipDJMjH8n6tVmSeIJyUeqDa+kX7
AM5YfL1BEGKdhPaKqeXz04q2RXdIZAouKWHT45T0GAlbJZy3wfKZNfQixl6qULIsRTUgxx40Xggy
tUhtIXxiyRaRGYlqUC8/ebBBm1UqXZRANzBj5mlA74oFhP5BbN0h/3oUNRDoQ9WAKDylgWrjGqpE
e+dllCWzgEJ/EBWpJyKWkHHS8IxsUD1XFBa/cVy6ld4upqMMewC9l/Dj7jL3d7OlY/8MQ67dQF6F
U2iwlsIKVRxM44X6qt+jGYLGjdPcJ9eMYpVVGcZc9H6xmfUvN87H26/6Zj/A2QkmdiP2BfSOPFed
VAw0oEgmU1VmB7JZYdfjHwES8vD0iX5WdyeU2dEHYrXkeP/qsfN5l4qXDDth7VZ1sSeYFSuGimHx
yrsq0GHW4lnYW8RLRyL3TPowtblOX1ngdt/PzkINFnlxgt0qB2KZspeD/xFYihbYRtQvMrlLWttF
ojdrjfS2t91+Ihi3E6EIK3wBLgrmpoGY+bqW9TJqHg/+HHtvXqLl7wpvZSpW8JasQrr43gKNS8tE
zwfsW4hlxB93QbgINBYRlm3WeKjtQTTUNPH05/BhOxGnBUfYCNwwTZcx3W4ElOKB0rRxYsx4cTC2
9dITICT6W40ko8cwuzl+qm7ByMCjeM90z5KXrPS08FgRXK/ARsI1gEYuGJysudZR4g520ipsaX7Z
fngnc+G89Xq1z+rzZbQOie9Yj6S+XgCPDPP7kK5lWFk0jfKIVeMo8cy2Eu5Cx08/qgMJ58JoTd2b
yiGZwtaUvTngT98hJ80hTOIqZiEkVUniHQkm6+H9IvZ5GS9fJKsuOLywpC+CAyUUgpURf+F9GF2E
7mfLIlc0ef1JK5XXLUuhQOKQ0O7+PtmzvMVg7N9av5HeK5IA1EJbfX5hToZ4P59Avjqlk6TSet6S
evLGG04GsjrxqUuiWP2e88uuzO2VG5uTnrqVlU51+iTm7R6xUDt55mayPos5fvFiCBqVVUvxHH2e
CFZt0YVN/tNB9Tpgesy8utWl/294rgq33LF0N0eHQKPTO38pHeLseU36naHJLFzXUkaZMN6p3qMT
yXqm5hiRw+1F9T7xNQN1XRbHYNmUqFtGCp3GINihgTBpfnp5l0PIAowJ/m8X0HFJjouHkhpHOrO4
Kv8FfVOcaSIR0JHU08TZuyrEDyqCXMJCbydYrIl4dxhJ2M2CIu4ZmS3bUndIhJHrcVMK3BkLfdBy
ENyYt3oee4nIOPiNR+nbi0cV8DMpcqR/KCIhNjADVO/JcSh6nfTeOGr1OyIXSdBs0iEIiSDhwNrX
Tq9aO6DZNm5n/LqmcQwhGw1AusrARiZuEnxHEuT6+DJruJEwVLVPoNnqS04eKDg2jOjOA9zv8+DU
SklJvMtmElGEywYHFmSP9MCGDUNotOGmGIX7eYhYFMD4tDPrlhKRAwuGmQcHuLEY8jKvZUrVhnir
Mq/aF2pDZq9LRsPcmYEe8naJQ6ugD6WeTLBqFimKrQHHGIglm8FjwzhQQKMul6JGtmoApiRbaXtz
JkW9ElWJRod84cm52GzdBfFjC3EdS9ibX5NSRkpD9b9AHqjGbgLts7ORBCmT3VorGqOZyXzu0Bsl
LhDvkdsKfEYN6vVQVXxhSyAYMb0iIAgCUefGq3Fi5Bpzg4sjt6QnpK0yyomA72sfAPqCw6snbsIg
k00mLc76mzXoHx5RSW86etkxj9k2Q2ArJLwFlf7ZzVufm14Ctb6L3I2i/CQHmEX+PrHM2N3moU6F
vOxozi3w53cSr8YZkEkx+tRaRCfqz1gCsntK46z/LrTqXy8vhnlTT1lgigGgnSVon0UAfdDHIryf
+TJyh9CW1QMc3H9zbQgb3FihMgVYsnj2Gha+WE+r5MKEWf2TlBuFG2CBkSI5HTy8L+lRJcHVHJ75
qfEykoe7Sa/P7Sh9H6ckWuOak2J9IG8Fv96wdsdYbIo0RdH1iA4Ou4XzZoTU1UceYG9oFhU5OeEB
lRy6//VZLyC9Q4FsCJdbo56wUrNV/DX5X8cD1FcxDVhAt5zuzHjSkUj03fJPQ9TUAhL3sGqejEYk
egAn6PhuYV+xD1r2AtTlMG2HEbW6P0vDSdEaRaBNI6zpVWKJ5RRcnZ3HppSFKxlzU86/j3Bz1d1Q
n+j+to85LPCYf/1wvlD6Xi9mx5+39124ZI+KuoKGKM+ZLYiTNuwjc6qQapGkaCphTcIqjTU7UFvN
815eXR29nqTmXjuKjkw1dPeysuO2FzpCUOnfVpGxVVDNnXyNibv0l8EVmdYMz9BhXB796DWoBWhu
OueJqvgHymt5MTLENSIgrDJKnyFFhzzZcdotSThz5UZHw+iKJVCVanxh5VgOtYs/wCISZPmZOTa+
V31xT0/gBIIOQSAcRHLkTM+ipjhXp4RjBlEMiS4aWuMzAQtPugY0avoOGgpWUGTNh65bm7utVrPL
taxyAJUrVIcxRr/96aBYsrK1C+se1oWQhAl4hvQA4rM9fyZuR4waktUsuy6NOKz4pMBWINbXGRJS
b9/5V6DsW4J3vc7t1w60fRh9eL9mhypGlQo//O9I80RlEsqr9yo3u8qUNSqb4F7NW21j8SyZB3yl
3Yv2pQr0s+gcQCPxiKIVGQv73Cv5KI7IdnamrCRLwmeCK/4pmq0pFzU5rDHdXh8rsBwkO3uGtsBk
J0gvbZCXeB0muPT03cmMW1LBDBfMJv7ncls3rDe1di5h8mnydCbNEsJV9iIuzLGB/Ud0A3XYdLP0
6rD08jhDgPRU8r8rSOGG6hLo0b5iVSWPF+yji+ZBbH95LWeZt4/cf1bmlwVqsZDn8am2ArQVjOV6
nLtkvrYEOfbYRNTqdZ9gbl93MZSggf0Dz32DN3l4Z9Sk8hdP+nAT1xlIzaYQiw058bz7jv0KKIpI
82MDIia22rsRmE2LkC/QHdQoq+8nz4E+I5KErGacoe1wIjHYZCcmzCU5HCWH0cmwvC38PlJOubum
2/TXQh6hIui2NiahTXzMYE1jLZqTejPAUeyoxr86YzcUYe0R+rPd2f/OBwAsGWhiKd2ylzRTVdUQ
IsTBpdiaffNMTpLkP1kJ/LoMLLiRp88yua2g0XRfl/x7aiujWthARaZqUFnKdgXHKc366TtUMILH
rAs6YqI9/6jCzIModyIgG3hjHa0Ac+5EU0Fhg/KLosZHeadENK7RBfQuJ72s2q9TrqPn0fy8GxcZ
qK5jjPJocl8g28dnpEESwmkewGDiCjqxT8frUP3v9D/Itt8lIPBOxJmYZNrEM1CENMsmk4jsg8b3
Q/LZzkd+hz76F5pylPXwOwE0Qyls/+47lx+No4tYrJUaf1xfBmdA7EwIK9FFcbDM+9A/K8sKdFH6
v+8VH3HsnyUm0RhSB+f3BTajl9g/jl4FKvzunYWOzL+qvVpKoKhjYdHG5s1POwFRcYWxkH5030P5
TjGnHIY8HxMwNwAKdOsCM+uRWl6FkSXprxoyZYdzxABPORMfXQrTtbjmfCqj4QRWkR+9cF20KcG8
1RZzXyrVl7qDkW1trODUEzASQPWF5v68TlUvyhEI4etANXS6At7RBRbe7aIAcqMJ6yO8grduzMzz
n4E1jcyGEol8VnN6WfeZmNrenazJ3piXDfTddwiS4yEZ8OR7EgRyK2KM74G103ImjbUCwC7S3Rbd
BOUgNgCnd9mqutv4HVca3qNXPW9+TtYd2GbpZLHA9MrPZB/W0dxNJVO3xv+xT13RA9oPDs9ERSR9
4spj4xt4eRfXBW8xjLnXLRpY+/RzoZS6wsRMKoNgux4x8SOxO/wjqYvGYpAmFpqeWn/6ESpMHs/L
p2/3nhEpWMzf+CpjYW656nb+mlJyTHizUvnL9acza0Ae3u4WmrVv6Lge/SsI9n3vtlHqZ34usXja
oK0MJnJTOtsu06g4cnnzEurLwkZminFY0XZCd8MC0QQzlInxLjmMJfBy7b4BgeZPA+9nwIYTnYmL
sJteuwxnW3LIpKIaM5gqsdsk64Q19yM1h7EcpvafXt/Ov7SfkUvisVST/VNcNS7gmAJSiFoPUdv9
BycEuI7hnWntQxUjZkRby92IYr3/icEd3sJFnKMSdxcpWYObi2Xd+nuaS8FWg1GCFmKKb62ckICp
HyrEnkWv+0nzrpRxLkypB/GoVAso3SR00IbH9wA5bWgIUwwikyLHb4vipH4JRJAEgRU3jEVjqnU3
vN4Z3WiWGZI63bUSENoTJeJHKqUDmjplYNjWZukBgNbUmFGX2gm65n7ZYysUw0m0Q6f4mWjZlL2m
OyFukk/JCiB88SP5dmOIunxMVWv+Q3qtwd18jHqji0/fnQ4/Y9tjZGF4oEGWgRzfIChXwDsGcEPo
Na1DU+1z8QpG83hvDJqYqovAAbYP0jBOviQcwaQSUfRMfBbyoQqSkKQFJ8725ngm/5S5qbgEISc5
+1eh9c3TLAiI0jD/8PO9crDmReHgfjOGxctS+GOSTtQxJ/6PAcPa5WerB31riDtE0+6v97kkyEoE
GXa4bJxMlZBO5oK2jERfSzRDoXMJxAIyfKLh2XGuNFRQUVp4QoRhF2E+pU2Wa7r1gCRFhY6+YU0+
KF9My32fmMdJk6gbfj8b8DpGlhVTAV0bIlvzkwlzJWle7Xvlcso68Z+l18/XE2qNzy7FHMLFozA4
1RkE+zaojqQKDUVFFVFDBx8JkE2Z+JOk/pWS3+ncUFqyxq4NaEi1uPHOAa2L5PYDx5D5dGxhHFj2
hpFbuXhzG8M8SDPPBGmwivTt5mY6mMjRVOGh7Sr4LvFYLFSMxV7mbT9tF+5lrj6eQEFnWbeceg+N
Wzg26SfSSG+is7u9+rOobg4W4Yl1zOakdi28YhDhcwHFrnq6Be8SZWxSwuUPX3pQI+Fj6w88dhyS
371O5zqmpupU76cExPePqwhFMNDtUJJjhTAMH8femgeX4XRA15fvT4ikXHOnxYg+9OyJnvRbiFuW
biAHy9jcX9Z9FigRcXfc6dQjH7dAE3jcQH/izwBvwRHK+cFBekHWSYLaMAV7pAg0wrgx5b/Pvh94
+lVTnQ9bvAYvKWBNJqh9qZTW3uqZVc+Kpvvqqj7z0372Yz+O9JHim5smGMnL4wMm45mWsaURzjSx
BD2c7LujPzbafHifRVe68PbdK85e47aSxYfhMF9OdT1QZR258b9zTerpaDWUTBJm6dD8x3LqvK5t
S9SrS/jOWs7ZJX84WssqMcTB/pQ+JuTDtRMaH+SnLrnMKCZT3uKkydNN034cdKaB4fj1FHZLTrRq
prWEP0vJn762A+j2gisCv0fswKXbR1iKAOC7YR+AZXxRWqCp+anNFq6Roxy1Lk34GNXr6V+sD3Dc
oe6yrVvJtRjNkWZuJnmX9vKCLQ9EisJzyuCHdVjPSTbBNCk/eQBsNcaLp3eSgFRQS+sA5TM2WPnE
TN3LRxDe4nf38eENFJ6pLVYM4s//ZggJQcHJf/n2pcuFm5bwQ9sf200QVJdCohi7nExzzuwlEE2n
ohmBdVwasIJOhjRpJwgc+E75cYprZwnkzd5ExQHOC4BbqNqaAgG9Xe2Vt6m0wHyP7UyXDznEh3M3
7xmpUt/OKtpoFuyI8a+BeqNsR3FagBgNzvJr7tJaXvL4my35Wq9A5roS5NdlTtcZnJiazgVL6MVI
CHdAIEc9tQGPHa/Z86rKZxMIX2CNsyt5buK3wm2R54oGS+HLOBotjdB8KkHv93pl3FWK2m9ahs0f
wfH3VBDMSu7o3ULElvE7YqQlGt5zwICZJq1CdtpGhv4F9QY8LQ0Q2ASCXaKJGaIY4bZ+uzJX/XCb
rxaZrVu0ASuxzTC1TXg1aAllXD1FcseYbLGJxZXgphKBvKftaKGJxLeezKU8rtnPrFD4JuPOQ/5+
/Nif9KhSY2vbMnzD5S8O1NTslfLHNAPiACleC9P/5QEhpTYlTrevGlxv6z2tg7a/XCGY6OLt0+XQ
OWrUq/IDc9RmaI6uT4kzXieGlxpVw1/Q30gd2BL583r0n+u+hOC1Qw0lcx3mfyp2sH9IzHn+arUP
14rKOKICWPDUi+SGuSGvLTg7R2o7uIpZd90BxbuzS972N3GpHtCLvySvfBdqmbgCd2bxcJVmcmj9
h/aqHpp1gkjfrofcu/Qv27jOKs/OTFeXRVakVO03UXyYeUPJgmXeISG0v4iZjTOSODw5KrBKKWyK
cShMjP0pshNvkTav+o7Knrg5Gn2WojXR2p7zfWEaQeSz7/lHVy4wPmvewHPUdUc90Mhs0xFvEZQs
+tFiJW2YSuLQYGqluBpygGRjMPfXzo1TqsIL2voLmMDMbJgWk7BvH8mk+7O5DpkYlQifLEGlbx1Q
W6fPcBOtTOQT0qQBKVMTKvh9Z/ox8zATEACCn/yIlbS2ws6SHl0z5BiZ9Gfhm9EXOgph0JRUSLRo
pSbhpvYNospaOR15eETRU3UnFbLLgDJkR99ihkGdfkbGTNxD1rGvd2ocyRAfEK3dOho6/Pg+Xujt
XH4keLwuGJGVCgSj2CDS2bTG+k0UyMKPZUHEEMv5+RiCWDY2yqDjLYRm4eEqzBJIIxrs9Sf+vSRP
v3ckzyyDY/qunEN8CQU6ACxPOvgfjQwdvhTK/BI/gZ+lOGVzJGsnlDxH6bnnwX2WmwFUoWyKR3/G
+DcSp0VC8BcFef1LvOGzJYbshz3AuAnbXyA9pJ7h3R47fsHCHweTMX12fuMGejXJKMXkBKTkohUT
JzVT4XEJpzOrgfACnaXYWDiz8M70kwQA2dob3IHCf21yJSr+bY0G0ucitaZYCDJf+vOQLH2+wS78
FbkZiOBX8ect6YBpzOyjxBtzP+/7Ycx1qy0I1NOVQwr2S0iy8BIIWfLEwFI8mBqgwBOpwTJcrtWW
8nHO5cG/BPQ37djqb6soyJ+XVJieq79q3S5CU57rrLq2Bat7c726ZNI+dbx928JTGX06WHl3sMfL
4CGXgXhLBcYsXDWAg7MmV1U7xSkIDpzD+R83e9yZM6gezdKK/gGeSLsZs45AtB0iORbqO6Z0vQaz
w2awZSGDybFgMrrKTXogKs70AI9idI91vm4pFEehsvPtNVQe++kFVtmkg1c59k67DYFdHhvIXozD
EedA6+Ygp6d1IGuHLLrCAgm7XKruuPQ2KdJdIwfXd8QHHKneDwvpjmPHcuv30yh7lWjiivJvWLPn
WnxGhN/A2GGu/aRlxbl3pk33wwARABni6htuFIJyv6nJ6Jk6r9bEyFvgRo1Rr+0rrQjA9Hm17a2Z
Y9aM+i/TOdUe+DHxXQ1FCpcBmfEIuufMOLtHB3I9ZzVi6bayMa2Kt8TaMmgPZ420f2/xcfjWRv/7
Ig2dsfyUcxc+cqidSeF4OqJWWewoq2nPTWM1mA8mozcw2t1J8GNqRM9PaEPNZYgfZV1qvi0kK54D
B+f18pYyuyDszeXLVhMkouBvvQUSk9P/Uhfg5PRU9bakovflMcCRK5mFD/rqPRGdbe5BqUDTpH8H
G5I4kWxN0vn5FZB5G4GZ9hgBkQ6Q1PnoikRcD5EOoUJ/g3LfbSi44OGQO0m/i7yROc9hftvBQqBv
WBM6QixzBRLyHls36lfhK+8b1nfSTJ5nRGJ67YUr80/BM+R5btdvzFTHg1Hxiw1lzE4bJ9q6ki1X
7VyPSIbB4DQvhWeBHrJMmHhD/eqmYh+nHuARvQzSNrNLpeYQIpOErugCy7t7SBNy73D7ZXY7J3TB
N93UlyTNYFhUC578RuoYH9KMVgRXYi7AN3b27elyN4ZP+YrISG7gfL92WrsIfVa3pwlK8aqNtCvI
44vv5xpttn2CY/fmNu/UZ0z9xXBhFrsOx1yYlWlfVnYgpww73aO6Fc1djuJqeDSbnhAuF4b+7RsR
KZzU9k2/JpIL1D/3NDo01Phq4eC40q3Skj2XNS90dj/rBEhc4sH53vyDPGhiWK7w7wHakXYt5egS
3Sl73bK20/IB5fovbwWnZpgUxFQ0Qy0aDhHSO2Cr8gKtmQAsK1tLrfHYX65sTH04bZC5bDwz8QnU
tFZQ4iG3AEsjOmOoekN+39MVVR8/Q6uUONigYlLLvY0pW7qXc+3aQ1vWOQkPRS88z0N1vp25Wf5Z
IESO9HORLlJ1V1zhngpUbaTowG/INhGmYYS4nvggBugv8HFSuYAVnHAc8MoXajBoGjW8hmDR7/kd
kAhK5ch1qLxIBeDmaIuPhDQGoZL+srqrgpoqKGlZUilzw/NH9/JOYff6cSD3dx+yWrqCPkvKoL/F
Wc96KUQbAzF3EbRTwlqTpO2nThMYO5cHVMFry6QcRX+hWEaHezu4McT7FtdNcYitGKiteYNLhcu0
TkRPSrfABGU6hozZwSP56bX2FJtdk/c7UN+6yNGa7x2dtumk4EV3I+MwY4Ps9Sy9t7PMDpn869df
KA2pV3Q1MmGDJDKzlndpvWEKmT5V1Iwl5wWYWgVd3gMEH4RbnjjHHWu39XbHAowYSPa/85Xsn1BH
CvQyyW2qLb/WzxUJMo8K0C1Ml973oNc5PNLWZGDvSthKaRkFCDZ9+8eevuCDuznFVVbp9T7fHrY6
UTeeR4JDPB6YN+Yqv9GAr88uakHakSkf/b5uEDE17RAR4y9yeEVisFiInRvBhbJKdWoj7gtX24A6
MOl89O+6SwIivYjeAQ3cPnXhsOhfUbaB2b0FyT1bc2K1328jaMaFsz7ZTIdpKZSJJAu0ExG0AvY9
e6JHmPLXr6kjdGFDQGZTjqCPUD6oOJsISkugI+STzv9obulhDR/tSu37N7IbfKCO42If+yootLz2
YeroDX4PoURvFhr+wf8c3+Gg3w7O4VlTQ/SVxNY6Ecc43kI0fxQ3LnmrOVYofT0piOeBQ3WbCk5Z
D8swei4ri2MMh0+LfmQbuOxPmJTK9sofGKwpLNBFRpNLk0Pc+IAYbkU+mZ0q97sECqPJHUqLpLH/
JhRtPm0yycEhdhW/Fw/oKTn7UPh/jERxq0P4sQx0lJitULTsZStww+1eQB+67J3rvBbm5Us7uFwe
spX4JZJXnyJS/bDHepHK1Wg3vBVHgwdGB0/JyEVqZR86V2kl8slFuHYCxFOZpNweN45yANOjl7Iu
RNPFt1t73w3CYGfWxDFCqLF4UJt08QRhT+K2LC9TK/M3sfY/lzfMK9075/YZwmQN4CuJ18DlKhre
ZXT9jBSZYf6Rbni86afNuFDoWH59xOfZG+GJRORnnnYJS4u2kUl8bDpUXJ4C8Um1X5GJSQprDO06
w4TWOkZ5Kjb56l2eoDQbageehk2EmntYjDXhQm9sNWdSxXjW2VSY/ZloRGb1Esy3N7HJvQD0GnAG
ntHTfy+kKdIlT/qxHgG2onYkMccO2We8RSohCLaluF76dkItgjryXyT/aD80f4eZZysSQeTSjAvg
4r/J8lCiJ7glnilgovod/58dPrVVvUn9KuD0NxKuXI1bwt9thIizNPv/DUPogQlcyi5gNyOsiRU1
FiL9TXJVNmSX9yq/vx3e/YDByrSSoF0Nmsxo7oyPAIzyXXXJPBwzPM6sLu5Zm/5Pv/MW0kN0iAX9
6Zkq178lVBG6XWm7JdUrIGVfOLr1LWX15dD5U8Qh8m2CzK19Vorb3RC3VOWKD6oAjuSobjYw7S6n
NhQLu+b4hvrxTFzgAnYPg7YkXlaBEDdQhjJ9QOUdUJM39L9yC3AsFPBMLHHOq9cv5NEnj9RzgVBN
pW6aJQr4e725ZDdLour8tWFgZpWUsAwLNNxchnS++g+qauThwq7PoGg8TxjqlFzryYpHn+S94euk
vHQyJOe06A8Ap96grqv79iz2DEzfVTHjk1gTnnIaN1r918Yt17i5askkAuMEzlMwhUcQMMZjKqou
CvE7RKM6Ae6geZJL+bIUr4b0v9+jJfMaHKZVZS1Ro9T7KDfVS5WDu4Yu/81Yhu+G+3XHcs+fgZcg
j+qdJPi4914dNdrCDx2RXfi7FwwnjJL/T9eFYeMliyh1L8JJxb0CTjEPDlPAAYR4gY+XJI7bwYOj
kVlmsbv+2jcWBAO6q4xMr8Xgr+SMAW2dvslrP6ySie98vjdWtIgxfwpKjb+palKsit6fkx9C4zPb
XGSA6xi3m8W2wczGdxNnucoC79bR1VIX2ZXPPot7EAxVyBsbpGw0vcp3oUHSJi7sf/JfmOx3P06M
yqGdD0S0xvsARR9+tdo0RzCJwS56CffvKTPOyq1hMFjWMvbFM98VdntC8uWi+3iFU/2BHPIlnUM0
RgIoAr44FmTGckrx9e6iLSbr+OL4qZvYXG8/unpa+5Ovun3B5h3Ir9htNH5d9NepXU43iqjehdL0
FEuPBYpEV3hOEfYNuBhR0CCN6znOjw7RDBQ8PsMzOt7ILeIFKxrPeRbScqt8++pt5ll872/0UTL8
lixExYZvAYHDnsV7GvWVevWZGKqsY7+AZXYBgTCTZmjYkcC+twJGUex7OwiU85Eq7SJER36lpVbB
X0Tf8BBTh+b5D+zlh2+TDvQj00CqP8GLCaBu/0+Ytigy2E4LFErujbkwgAbRlYuxNvMssk6nuFa1
gZMchrNWtWYN8qIE5p38Vv2x4h+piqAhiD4z6b5kRjK1VzwZv/ifFL6gB1M3OxLRXnJ1fq+96dao
lbSUzshX55b6Aq5FEl3Y7e8nxkBzCrowZnMtlfwzNLRoURcPOXoklpRsfPfx28Q0VqcAeA2KgPtu
mEgYugqDz3cwpvnNWo8TNHCl7whLFPveNbdvgxnJsV7OkZdWiu5BV9UwN5x6IMZFvnDJ05hjgo+X
b7W0zZ0WkvW/mAIQz0NoAlWlYTyJX3+5uajrWy++EyQY34haDeAUvujHamAOj+AOwO3p+gdekVAL
uIbwFv/lNEclGho/Atl7sI/AJajEVtSyaGqv5WWve/Pq2BqAzW1HN4j5eRJuxWFMV4cFXhgzxBk3
bfpRxUTfFmRLGgAR7+TKwxX1c2gY3lHxHrJpdskouw0uBEJqmd+GFe93Tl6MMa5y2vtSeEPXr6jz
MSHteNaT3K11Ux8vJJ7/SW3Y/1zmr+ydncYEiKrHJam/fnjDOZRBm6LwgDHCs1Xf4weqAHaa1joP
0T5eG/M7A462vKXs82qsADustTpwqRKlFjlCJY8JgAao4FjAHpqVWCY9mdCIXgP0VWkBwxNhL8If
YqC0HiTD8iOH4wXo55WweF5yhFJosi1liJraDpkqjM0NWzA4jTkK4PzwW7qR86suJRBh8Hyh7j5e
WbtfaTahFvtbQMs/OMPZoc0rGRG99pwxxX1jpnRPeZ+1BppaOLt19WYNdT40emdD6mSobqsi17tf
hvVw15IWnzR3koTZMFuo1beTgp83Cht4QwTEVhQcYbGx7icLjl9wlZX6GTYKxuSog5u1e+hyRc10
8GO2wyk71j1w/GyEWaL2HjRMKMU+PhWG678oOkkhjLQCIQMG+r/EaTD1+TS++u6XiQvtVYvt4Erw
a36UGtquxBp9QRUVAUAzwmZUzdk4NhKsp/qHbsbYvbyiP29u0ks9Pc2XY5O9p9el1ZDm+SrQnCQR
V4iyPNhQ6Hj2gEnz71YWl+BlQYNru5yuovDabUnLk55/u3Ss4Ao2KtBwXl32XH4iTiUHW3tgY773
geD2/zGRhmxekKw2AKRBiK1Wb+WwhZcB7m5rIUIhDf50FP1dBvaYzX+UmTnkgL+vpGNW2qK8PZ22
C8ucCYUUJLy3lK5DINVvxWVgHr2pIzjGbs5W0i/1pHXc0e9OiQ5Ms2RLNbW+kHPEI717iLYjYxDZ
CvvKBpL83jyFc1CxNQsoP5P7E9RWcD15JgfVFkYw6pYG609RXiKMEjAN0wALC18JXKWFhuCM/uZp
zdTimEGRGZWf7tGhcVS8ERQqTR0XLFR/sGJ5yV8frdOy449zvBFoaF3jkPsLDJO3fxkMoFxwHNg0
eMjGxdykrld+KElf4C2dKREsf2RngJTRFimpLdTdbYPnQUPiqSe/cKeiLi16tlDo/uLhxfjo1Ohn
27ag6JZt9SeaiNxqeF7MK88tcwlHkCgB5p7EnHrEfTsctRcoIgudNXDzGahRlRRRobKJpOLDVsub
15zYIGEK7tJZQ82CZeFsSeoElcP6ZcyP+TLbNupi1vL4auclgwAPF9HK3UeVkXJs/pHwEFGA43Eq
HtItX3i05S404Ws634KVQaybR0NzueH3tFOJ3FBGtX/Opb1kaITnJsuUcHUPYcI9sCxtS+P6rC5U
EkNniHfsnVkIHUC1Jt8k2laQLTFigEAmL9wjtaoFl6VVVDwhXt2+J5LamExVe+IwMXmiu30K+bdb
V/iuMUHSu46vJ14SCtcbyw9OV9t2+mMZPPmIvnzgvK0cUaxXNSd4zl4slsF6K08YxR6+I/rpXRG7
WSuzzRFIMu9FNbybqberblhpVK5uxBLZAwy7WEdPsm6++/kzpc8Od7HWg2+WwwI1Dc2pERQrbP0Z
Xe0RhUmoGs9HTUQ9s9VtzZQzlicN8u4F4oPcT2fFN6icpuBLdF0/SpRK9i0zZakhwSPsKXUpWK5x
FeM+/Hwks17Rw1ks2lViuT5fuGpRRzfOeqUhcp4h+lZ9JGYOyu626vePdR5yOmmF5dMd7rNY2/qr
NL6wUIc/9aC35DXZwE9V98a/jKYCnbcAAIB+U5ZkmxNzgkEEfs07s4PJJ9duS0u1CN+gVoIBVNvc
x7ygadknOlwvNbPByIcNZpYReOeL82cWhI/23QYIDbOt+SW33+aIxTvdAslRa9Lpc0095KCT0CvX
VJUpKvkQKgoSRu8j3WUcvSZik12iOIOdxxpEE/nBR/YpE6Yg1Uz6sz9cEvIiLRcgjpHhUVe9mgIC
kMm+VzrXtoMoVG/ZeSy6Ss5p06KO8H0Aw4G0m+FH6nV52k1CDVKlMEAPG6wVzpsKdQ7DGYKGlL5Q
CBe6O1wF65hKw6BznlbgDCTEjaEcUTnKsDXzvYJkuQ7d1pDxH2YeznnoQ/DFwhSi41e9mb3esERH
WfvTqvt+IV1H1wDlFMHGax9Y31rsOoVWgk/NYbZ6q4UsLNxIwrojmV8aSzSzflLw2azb5GBqnKyk
d/w6mbg3dyNtg3SKWSMThO3yHzsxjc3Za4IUtLxSHCS1nD3xPvPfmaaeS4Eqkq7hXlqReb+1fPR5
D8Gu2berp84tJfgRhIQRTH6MFpiIRLBETTrMjKYvUZECU4keWnX4DFAwwWp+O4rLeVEpDJbQfp4G
Iwq73d/x+Tniq3dqn/Q7u+AT3nk4NbPW9J8ZpfC8py7Mi5BhutG5L7gEXUiH9vWv96ohMsqUOfpP
bBVER62pkqPd7sJ7MOQApqabs2MYUN6UJ1tMjIIPp84d0KYRORqfbzZI3aXuPQJ6msITaIpKw4yc
0bGwo2Ds2zGRSeNJc2UkCo0JkO2SljofOtzme5DFejORGkmW9Mn+G7otLmzKkkq/4jkDEoXLF48A
OKeor/mK0T2E2zXtR8zhu/GRnL3QTs2k6pAlbmtg2WFlntM4D2PtwTM5bCRaAKYkgY6TWvhRLzK0
52HFWN/vlCtGKuhDBAEt5RjKiZb5wCQTmScqvtO9xVUiNM9ynBv7/eT2s5Ftgk+sAaDycKsy9QO9
bY6pMoUAmBAnFC1m3SDUAcUXqzGq9DDgjDIkHF3m7ILftPY8EWZVpG3N/Nra3VR0k287cEuwg1wT
edWWArYs2yYZRwCczIHTXFu2C485qZtIVNa9CYi/DbYtXInq21jeJrBq9DHtpE7X0MDWg8Iyhjq6
iI1ZehRkhDlW6UXRl1L4yZ/oUqrCIx/Svl/F8Jb8Ow0wV/4vQ8PdnZNKIUlxKdKhK57qTi2bw2zy
BI0VFzjMJonx9SEN8CaMS4so/CbD5gsr0UR7SbCb69eclxBaV8Wkz9Rkh8LLBQSbXXmLkyoDoojW
vpmO85BwPrS50mbFjzoPm9EiPa36Rs8VQNZXK8JpB5nc0lGN+MqUEcjoZH6q3M29/Gk147/yP2RY
fgXg/qoAGZXnYfRnxHBOI4iQkUC6SyLP9mYuyjsTybwAu6XduABTFdLrJJVXpinIwGJwJlZgT6wP
sQSvuf2nMXiIxoF+KJhmwUpvm3YUzttCDXG85q5tLWE2/WGkdQszaIHS6+hK+dIx896NmPSW0ldk
TRk+1cU8UOrycasQmvrQvXwQ4dyJUtJbB68dh3iGO6BGYEk2+Lx6pARMMbJnOBNsvOWiw6VTWq4k
Xb/eUWxKwPq2ZODBI/eatk6pioXZZJOmEMYkrpNvdfSKdRWxMzP1IresCNojQps/nOw3pfglrMzx
Agu+9jf4SIcuKUAuw3ozk7OMA6qkDas8QV1JSJlMp8Se8e4J3W6VbtvC3RJ1t4MowsBtTmjCLB9+
ek3pvzunijiXP3LwImKWhtkzfxBnDipNx9YwYhbHuIpxLVqnZZHAot2j8+X/afU0mxC8xfZVeyhb
yizYsGQK4trF+HonxxZwFtPVszqodvfV5TkV8Aq2Z+J+9Ulu5Fgz1/4aQrxyo+6W9IZfMDKRDUJY
PZ533mdFMau9FAPCC4S4w1f1fuPMN8Ci3IZwIg2uzhpiE80Q3XATttFkxsqtvvk9xK5aYVMy0Pgg
yhUN2z8Htn+tKDH1+b/HwQHPQfZb5GqpjTb0VLOYmv5TQlcp+mHUAEX5F/rU4R24H55i76ZSkXOq
0gfg+/02u4UX4FjZ0Sm5ludapZUYU8dPvFtYY9uHX5UsRKJpDzi7uu2icC3i/fzITikf9NcdD4C6
h1jQ9OYSVzxvS+HP7Sj7kIiOUp6gJ1xxFzae5gNCPLz7K2ZngdkwTWrk4XXMsJMFq82hW2naPBlJ
QnzeoFkoDMax07gRocv3ldoCtjzqDMlZKrcuyh08E+1FFyOkmdXCx6k0mtqUhtWW/8paVbYu/EyK
gsX09xi43AJurcGiUeND2OobJ6smiA8i2qyyuiX/WteVPLkbRQtvxl8qzeUubr9mn7DL2wr8iqWX
tFeRYlaZKBZVPbwr3153p1V5lwj2CmQMECHuCXRnRafsEoGHtcSY6l+dOrQj3Ck+Qhrim5zJE/GN
P/L1jV0LKMjZw/bPvElKEIXb+ONd3PFhoHgnyRVrACYdeAbmK7Utw+o3EGnfUkp5Z2W9WVUx/MHo
6vSkMnFMae8IOadKZO9vuG4vCw+O5iYMCcU+zJB1XT6OGILHjUodhJSkrW2bIygX+EUxBZmvB/2o
He7JhQaf2mPKnRLgBTFKZxS946G6KaOLXW28szjP5DO6BVaa5WMdWQ+LlnLhxYlpbqMNEfTgZjs4
qDEostU5Z7nsChiYT2a1hqUFEKbtK7NUYmP/vwXm0lOmHfJPZWl048unM5YdrY62pFgFhp4prQm+
Af81LBWubNthJlCBRLpTRtXkeol7Om26s/IX2eY4jKt9oQXYzDqfa+q2RotY/N8+LmKngnOQ/bPR
K5mi1YGUiCzwhckLsoSJkteP8o3u44u6iircWa6IloQmbJdsBGRZ4pTQu9WQ/9V/vNbstp17we1d
2iw5HUB3LuKbALh/Hxo1szvAS+FQIaaOJ9AoIMXZdKqG1Ec4Dl9zLAeS/cjxsjf+Wfh/unXwN+gU
T5j7URoVwBHzu/xN2cTqLLYNVAQvmN0d+cHW1YT5mC3KYF6mxKiMqwYG3GyhuDmMt7jWZoRqK3c4
G2jNZN0WuupdFhWJPGnxlqmFz6yVPyf9fY02GrxTd1svkxLt2IcJ2dWViWSnOgOl5qmyLdWvQlF6
poKg571pSKeV49VVXtXo48pnRSqWnzdx8ntri7PPkdUgOjtYg2HWPcrzUUx/SZrEuWoLTOlWfG31
MIecpMmBpcXZk55oIudzfpPjsOL8LwW8Imk6e1UNP26FjdfSFq5rtilAMYmFkBPOuwAFwWpC/0jw
rn4HQW/EWdTbegDWarwYHAlsWHDEyqEzOgMeisWk2HmtbKepyqyS8+Zw7l96slsvHQ6RzM38xDiY
CKGI+QMtlFT0RpVTOhMroi3fa1ra/XD5DqMv5YwAgzDSgYSa5A5qKfB4fw9SyyIFKbnJ7v5U6X8p
EQbORUk5WcfdoCZMrf7q1quPGI1lSLKZVWWbxoD+eMTQkaYBnQwvX+EhMtrB4Dk/BtS7DBx/oLqo
UyzRGbI1Uf3qMrBPggJ9oNZVwgAw3N6dm8gric8RzdikR0nT5Cec2ZylPuvbwX8c5EB5iL69d6Jb
axbm5b5H8pIkW3NHkPMR5Op2DXyFqyfZN4Qt+3QiJZQif3IeI6e+oHcVec1FoG/gEl6NFGwsFCEY
wyaX7+4v8w7TMzCpoUrK6EmzgjDCxLvSot7xN3OoaoV2CbQrkj1p6QS6wzi/YDMTdylRmpdinvaL
nl6KeknJCagl9ygA+GdPr0a0AFZGF9/x8Xy+h7O1FgJs5hmpmSCD18bZJCkp63P7+l8Hq510xFeb
x3snKk0TtcebNPEV+Aa3kaiIclwXlq+hlehtQmNHnC+VVzakxDB8vmwUgvgG4oWPmdKpyrDlwxg6
Y4MKCWxxSyp5hswmXIRqee5YDRMtSo9KKLLcaK6S1KB75ft+sudF7Y+Q4IGhvgbCpjoEsiRmDd2f
UmcfiFPN9Z7GTQHZs/VaZoK0+Xf765KqprbkfZ8X1stIW+m/sdjV0m5TEHc69o/Ff7r0VQA+Jd0+
7KCPNBwNze8VtGjZUsd9IvdeokEb4GqEyhgaBkO3uYyBk8dW/iE/E4KS3VhUn/Inmji7qm8jIxo+
bw+z1y0JXDrXGrjSNYz+Z43wGpdXAi0x3PRvffR7vCDeLbaLruCwlwDZkijUy/R65DPKCdp35jUf
MoqLhFqLaZLovtT8wnJQHYx265AbdNoMN88PStcWDYyY8Lxvy5Y6VYcZ6uFuf2XDwBfcV4sGx+7U
hf0ktJuTXSflvS/3ZfSvIfKJ3isv2Ujv6fgfIYpbrxQeHKBwy69IKlVTbYRPiTShQ3odeCvAtEo1
Hs3QM3CMqivI5ODtZ7nVoB+UPXBbyprARVwG1rO4kMyS4gDZGj7MOdHH0s++uOKxQy6qpDbaSWbu
RCX81A+Qp6nNaywh83L0EcCTqqBwvAK0la5HMhV9Gt7g/y4bW4RNlkImqdX/m/l8Dl5tRSrpegoc
S4+DUqM0EDMB9ZpS94PY7Fg3cbq73B+qcjBC3WD/tKEBzaa+DcX86MuWXR4wHLBBhDSuXmaIJVrw
EGoIFphtE1iFkknGp7LCYIRz19Y3GIfYu4noqHp/PSFFmFmo44D6HUr/F5bEIQPtq7y+5gleaJ74
l08LQRtf1Y6q2s90xYOUDtnmLy1UQiaHjQe+lnH10qzKZttSj+dOWMkUZ72AqDH25+8pZQm+WOIY
MNwWp79hsDPDgXT39gQMWHHV0d4wFYKxz+FMg/SL7cBlD0Y5rreiiTneLpclSnjMCHTdwtdErFKJ
T9gCmA8bF24psZLzMN0siNZkAZ3CGFYdKPfcyMZVsqqwWqYo2bNAhmntfYGG62/xHBXD+kynuWBq
w3hPzax19dvKSr8yvIcGXePhWXaCgRyuLk1sUc2yiCpDdu+XqouUhEWujWA6ZEn5w6jr3TnlEwTw
WzE6btHdUZ++yGOhDCMptw2bPLrMUmH1Dhg9fZg42cBf4RBlGx5z7+18ep90I5TMQirB/UArvXNO
hwN5ZExQ6nE9jcGHgRmggl8JPqLBp3fKi3Il4OqQXqk9rqRw3Ykj2WzptGdaxNyoY/RrZiX88Cil
avu8OjQnJhLeBepzghhr0BDHe1vFIiyXWdEZ2mitKgBPBh82dKg53byoaUFRehjQ4HQFvITTOkgM
YYOGMqyd3q6qarwKmzUov+BgPE+jMDd7BxN6Ix7+gLcnFsL0jsxmLtKs2t7x78LF7ww3Ed2DS9oQ
NGOA2vO9VeBZtZRq0o0+SrUIrEN7Gq52nWLdYab3blO0h8iqD18bYp4qeNaVE8Py4SB9nGIDHhQt
ooIxxW6yP/XEgHYwW7Ry95Ry/cr4TOKzRG6RoYvh6N6/jZfmyS8z82Yp6k8S7ML+UOzOwylD1Mko
y8xSTxJ1IXRBmDqZHZYigb3ZP8EUyi0q1JUkzR3gHPUS+LFAU6cl+Lv8hz5JuvkbSDjlDaME1s7F
h0d3b2Cttsnz+n1ns4Ep/jJO/8qN3a6tsTCpP1RexPZmDpkdW2+li5ycbzUKs5ACntN9gl22wlDf
V5Mn6rvyQhJD8etVXxQf8wqhiJU7tzO61wT4MsKbWdilcdI9smJufzc9uPwlXnPUrpwBF6zwJfmf
Y4PeFs/eZ3+kY6vEILlUaHm+TAnUbo5oes8hPmRxopKgFs+5rtMJ3iyVV97g+Ho/ZGCqYj/+V0ku
QYAd+tBr4Bd4JSjAwCRaRVto0CdwZ7rA4c0a3+3duJg4HPMQcJG02uOvyO2bvvidfreEffLgDsb+
K29asZtEAYQfy7vNxWC4fF4QUYHesRlWoFGQZeN70GejCJt8vTkVsuarKV3S3usub/e5uclwT3xH
yPssTGgaLC18XuTXIIL6fiGL3ggrIXmbxYATfyn55QYM1fD1ePY/ihlGNB1zWXopjn5/KY4Cn+uG
gkPaAqcz9toojhnwHh/gPgQQiaqwoEg8b1FGVVCaa0IqF8O+IuYIZtt/QWMRX2C2hLUxlsF3hZ7m
aJAa2IQXomRv9yraKzkh/PBK0Cy4kTvkhCO7eLrumT2ljYfsxyXbs4a5c7g0tahkAVnAxd7VPh6a
gmE4bbSOFWgypBDyKV2bOaL7s+Bzg0x+LbEBlQyxMQJlmo/M2ORmIT92hRcItAU+ZDQWNYimnCfd
EG1WrCOSIn3Te/LSSDbcVai845oaubbR4b/NOThSYgJWbtxaQfPz1rHwQW0dI5D/7B2LU8i8h+DR
8FPH3lKqV1T2WGN3TrFYm7pf2MbUfkF+bb8eTt5511W9VuoPteRw0FozeSiS4qCj18FP06BOGN2C
hJuZn94wAZ/J6kkNprnhq0gVYCR2d6Lx4gRHplN9NzpCQXKqiyVElMKCDW31yygBqa0yBp1MYL6m
lRRrZCl47jruTBIA1/Jv5VlJBhQ89NV1cNs8iigUHHLNlWfnI8gS98DmZdVOqnVR0mlvxfIhOZHz
U4C1ncfLCS5eUufTciPlwb9mrGHFc+Fa/ZMW0kjU0mfSPfs08Kx0AsQ+aRXsngRdeZ1Iu1oEfAhd
IS37zkpVDX//pEfYQbG22/XiEvjo4buBaA2uFQ2ei6XV7g5ONOOlqO9CSe5nusa9TdJwL/VAAVyY
FQjK3qaJ3h/7O/ME79O1UfcebcBUUHbd46Zn1ODtoXw8mtCtEruDhOeXS46zTxR1lml1o1sfZ6si
pHrUDh3bznQkwtzTn+C1b3O6JGw5N+qiKo44p4OHOYKsPOT9g3r8Kjx6M0sFESwRVB70f3bYeEqC
C0A9nLX/ovCnbt8BXrVMhas0C68OhFNGHUUU0W5Rxxli6x/7d5vFbRsOqzhYCPBK2k/FTFEiwGyJ
f5GF1hrrgEaIBezklotm6WwEfejD1suQiPcHq44BIlpTb5TkzgLLU7nz+WzjZ+vg06zM+jkIEryz
Qh+jrjRCG7oKWegEH+4P4RF7vYzZiviJZ4BmsC2e5hKwMizDo3/sAZeXCf83e9zHpM9oNsYy/zba
YYc+NN3yD/7/pVeiZJEdNJdoRsHEeeHVcZ6flq1JMD/pVpAxDNY7GY1tWtGwJTLhDO8uXMWadWv+
GAurBwb7d7z0ZvszX5J70DDIh0gSGnF7cKtLAMxuksc0wEWS+1UJwHONvIYOUZQbAaG8jDTFUl/5
Vgv65ISLj3b5jIeFbd2BxDr+GGl/Qt3yB92TdE8gwiyYbmhWDtWrEk7Ew7wnx5YpkDgCVFBvXcWY
dMqJpoD48oLT4FT7Wnu4hjhAG0inCSLLXPHcGTgb3Poq/cBlC5roei2wAXEdhMG2/i3Nsx6P5yqi
u9RIX9P6gVAYmERwKjhZayB88pXFCZSzu/kDGPGMIQeJDKQ3mEmDw+PMn8CRclcBBXUisJ4zdm1j
qw3OzeMa70q2qkgKTOViXA/WahmpW75VTXTRxiNKXpbzAoK0GQw+aGHXydC+em84CqtAABijFPZp
La3abPpRXCQeWUT81usNF+/5cjwGGPBpsqOq6wllVli122tToJfreuON6fiuRCnsZE5NXbLQYrvj
qL/YcWM6PFy4gKbJnk3LAL2MtXPBV+qkWafLKypxzmLgJb3E50cLIIEz6StuF6cd3QOttNUtcZzu
4C1yXePhJNoj5zwmdkkFW5NdyfgmdKeIVFPn9XcVDlHoBB3LNet9NbX58yvjRfYJjbutynqkgDgc
DseEXDUdZuU34h4+JCKoJnTSSg9w0kNT6KiQLA4dq6QIx5uTTC9iMwMV4lQnJo41nNSmDoq0ZV6n
N8XrfOCjH48AouYBTDppP0TA5or/cVSBOsHZV2cyCGucWX5428jDp8BCeJXiiG80nrcUm4lnRqo9
v+AWlwfWeffB6P2tNpW9FqSlvLFFPvYkUacQaJKyrG9hIBtwt/tBZOnEAtBeiHfY+0pvfaqLHU3Z
/IN6pvMLET9NHu5b67ajENySak0cVcCFfYBw984CYhEvw6r2c6IqyzFxhSBT929nZAVpnUoqMjRb
4wNp2SrDMt75d4H/7bIkP/rYeDyIOSSknKVMVpyshkFHJW71fc6gY5Yq+3YuZFy9b6+pOVD1LcrM
CBSd4Y+ipTq6tKeA350e+huGkoTJ14YrqX5Qz5K4wf3OujC/lJzdlB8ated8rXfbeP314gCYMoiX
k6nbWH/d42+ptG3gfBZUudypffxjtkmGTe5s62c1f9ydecfEu0BS4SgFSwzAqcqlJK6jIS63ef2D
JzvnNpFlPuihVMfs8lVGPfrvH+adZUVIZBZL4t0ZqzY4jt9VtQM9mHBZl3czA5SDD1OIPqh/HZHl
Qh4qGVUH53qkCGxkjAngAW2utcTatRolBaAyPLwvKM9QX+b5014nySf6QvbP3Szk6+jJulBG209G
lKNICZ3cBysf2wHRTH3XJZ25hBE3L7P0VPOKuRYyQU7Aau+DnOCWP437tksV1Y8+7581Tzwt3yuT
RYDBIlUrPh9KzLRIDOF18xaNtoOKCwPbiwEi28Z3aSF4SxU56xIF8sLOT8PiXvrRTS/7Vf4hOaKi
HBaPNjEHogss/j9Ouw5OKsv+YxW2ehw4MTHAcn6tLxsM3WC7vPMO/aIpLclHj86aXR1UnmP+CrNW
HUMom67a67wYF1hl99f1MlLNZsg0J+l0z4Q9/CFU49Ch+M3ohEeKfgfA+zue4MIOeop6cgzi+6LQ
bndqVc1AlBaWUAYZvZJBUw6aia47X76tk70dfE8oOJoVcQ+WbNcIO6MJae5zzzfG9KVsCyZj5bOt
3hYJL7cyONV/egiM7yM0OhSNrR9RPpVWXNVCC0iiw490Lnr6IwGHw+pphWhaJGfR3ylyV0JyEMck
JpgmPzsi+1nj0pNQPfkMd5GEDzzCDrXIRncH3vIy+YIvwyzn+Q4dOyGgBoZUqAWYuwB8qYpPUrhJ
HJNHJbclRQbtuDbxHMiSZbnfllJh5gg8WAg49bhDNRIzvJCd5GBM7FxG5evg6CjnHH+1E9pZCwVj
d0dD28TDs2EuS6FZMezRc7zTsyOtkga/q6J1pBGPRwYhGreZgJEwc2gMbC66dloUzDynMYzpNN0P
coLtHL6sRTnzzLrdRKFNVE+EsIXQJCN6w5thPVi45VH7VeDVp79EpZSqFVK240N6Ec9bNr8OW4wx
GuWNftlQW6jBZYBvidpaMT3gy1LNGsPJKWkyOB4z53msITsArfDsKP8Ct8087y3SXt2SRJuxwMRv
qOBXYqWQHXjr1zll4AeX8BKI91vCkEu8xSrCSkwHrC6LEWC07knW9U0zJxNzIL5tBNcVTRUDmdkC
h368Z640jKZDzSKE89u7JhBVemrQ7RkftfdMNtSwsJ/J/3J4fY1rVqmkAR6I4N/sE9a8/e2/Cb2m
BMtTXH7l9i4ZXR1bOyFwRvSMIz/cEo6NeFlteGrtKdx5fZfDVloq1OTb+yESTOVrbZ+6QNmarLn3
KiN6UxZUxDkFzgALms/vIUNIZsLaOT2yTP15PtMVYZtZangg9bcSgUpWs1TyzovH/hz2s7Ufrcob
fWLT+Qp2OFTFUaqgiXA7XOrBKWc5cFspDqsoz+o3+M0BPR9sQVMiP7NnI57OcUuL+55cfYl7ZG0P
GCDRRvexaHA4mWJ9ZtLHcntoC4m+sH0LdsVYn/D1P0uRw8+k1JW2qvpAxIDi8x69xxEk1Zrrsu0B
/dWzlmo5DciK1vIa5/hbSoC7facyYFVJ+uTCt0pL6WruFiEB8jdKBEK9qlHRIjsO26EuOsylS4a2
hdKCDjcb7JgZoARFC5icr2wgqwxlh+0q8BKZ9TCitf8bACl5Usdoc2dy4FfyFGiXzEWqOG77ug+p
8Rmn+N87oQyt7H+o8Thh4JThfGcB5LxXd4bUtQyuoEhlIDSHwR2s7SqE11PjkxFKOeFprELvcyiD
RxXC9NDZSWRkJ8iE73GGCrDkJrmwyuWeAopGgR/0GHHsFegkDFxvSnnxPybPMJewnw0oSoOEwFzZ
g5msOtWzb3iJ4IB8CyjGc/ULOLzvtVasSze7o2uJKujDexrxG6zNnP3SG86XUYhBx4BGmXbdzLxZ
Z+X8vPj+vPZgUoz4kJ5xEP0k5NLSRlsV7BDbQF/v1JMJfaqF+REcsiHex7mKASicWHC5cBDt1S/p
6sKzkKPO/5yc/ZoAdLWwsMSbQGf/IUHca4krw33a8vROB9huQ7m7E0wAdI3uIy9d4LjgD02iXFv+
Aag7srAPg7rYxcZpgR6sOWhDnNNAvBvx4MXCCm5qaAHx4gggKaNgPWUbO3n2gkZDOtoIPSHiTB74
DBL1Pskovx8Lo0sJrpBunxh7Pxp0DQ4xct7UY+JAy/kvX1r5KmthvxI7kFk5h35bDfvueJsUlKo4
v/YBGyfyZW/qPOliyf8+RTNGvOVYi7cdHTa6dt4XOTEg5SR+E5FtPTAIYc74SGtespqB7NyEPrUG
TE/vJ8tNsf+arXHr31URJN4VkIPTI8LOf9eW1ocUyvU5hciRWT+Me49QS4HIedZIV3OAnt/W/1xZ
g6LHA184HZG77v5pIrm9UtRydkwqw2HvUN5gZ4y0BCgykwJRNxdNU/DcJ24yjx+kfA84cTSvLYNY
jMETVGMGQJLKxMqCv1kYlmsOHvD91j9r0hoDmDvgULe0j3HGbIggTDYuacePt5/om8HcfLUq6/lk
gAmYD5Or8+sVGIT7KB8ejLd6rwQaVIjWkkz/JrcPcYr2GDaNLlcsPRN+0g8xgUb6bA6E7JNQvwLO
sb5BEcNaDNNI8UX/nYQzoMtvnlb9DXg+0/PK7UUPDCFc/N+K4byVGENw7k1whDRUHSN11Qnz7TYR
95BeG6Xx+rPeU4hdwx6TBvym+OCsAGlIYifX+c5m/ZQpWeRqMP0BhoUVm2B5yK5XTFB6CMWGglsV
gxrLOPMAtdZ7o2Gnh0+PkYA8ulozFE2TSrB62skUEhyDyWvEFs1+LOKqG78hHiCGXZTotGgikEf8
WhdB1G8uuzRc6Z7TsnhKdh8Xc1svCGZ7VOa3r7WxlSgzulUdOCeGBU+BNv6oxTrNAZEcka1CMYtw
jsazYeGfS5Ovv+2BcY/MadTwsiIUzNYsZx/Amm6dncaR3c/T2/zKKHu8SI+aJmlKvuRbNBoe103v
e8XgDff+AhcvN/B1xgizPZ2fZhJRdmrdna53Xu5+H002gE+z401aop6CNyFIp7lSnrfXWgybFB6V
u9Ua3gXpxgMiQn/ttK1Tx/T7fQruX2J8+MH9hRjppHC1fF+wOQWhrXZpPatlq1VAio9qDPyNXp/4
K//KRPC6CZjQNVHAKeEWMgL3HoyZuwbsfLcpofIo4vS6yrThfIY5MAcB6r5yh5RRZlCJrd9vO8ux
NckxJeC8QbGSNNDnGWo98l6YiVJqwF5pbP+iUuAh0ovUnkgq7cf8vbThPnyzZDgTak5acclZMKpk
ql+yvO3xSgdWphG+VYDBzMIW1rROKrGQdioQ/nqWv5SceNR/UDU/yYEhrwcvfbrecaF4OfuKK0Tl
nVEvnS/odqQpY1hBKhyHs6unKPyMWJXU3Qg8OfOJ4TvsXksNhcpS/2kMiRw5no/02gp35S2c8GSC
z6L3wI2eQgCLTySPAemZOsyJdZJPUBk4dd23KP2AYsBLODZerMSY/jfbb7+2t+cXo2LsViH5TmyP
fG6uS4U1zftkX9EsuwQadH46IA1CNAPY0nVJuxlQbdhw+XgoXj3VIT+2nPC5w9IQpuj3oqQXbco6
19jaOocJFCwUxsPZZybHmiFdpXIgdZkoiYXoBCIVWLPLK/efdzrFewfvgDvxNnYEJzML/j8UbgR6
ohUhqnbLqVuFlir44K+14PMSHUVeLwWV+nZKlRZnRFIQNjP3PbUKDwHvchVdU5l8zMBT/vOeWmwT
Uy5ThiyV0nMyVsHgDKGikHv6IecXO/sdR8zN5uQNXqOJuSg5jL2F7DS1Vfo5nERMxNclJdEN3IXP
6bghuH7zXovaRAxrQ5QH6PMOp5FH7VApClF08XxNgoyGDwnR1Adx0GA46cL/fGJPjSLygFWp1i9p
0qbzQw4S1Fph66Wdj4JJYVZBRMZv7FcfjEWFetvCBfoBVEzzyyZ6YGp6fgyo67GZXKy9Wkr6cjMz
m0VuxkEyRLE0snomiyWZQCEM5Skl/ksPYa7XIvszz9H2CuZH8yckO0DUquHAL1x5tS/tJyHmaCHF
mWJR0KK3/sdQMIVaLuXG1TvBmoY6xpceffYRKi5OMXfUUqtLEDfJEhMcLESFpKCQpXzH06hEwOX0
F+kPwlZSH2Y7rttg1F0JYX35kkHgRl/rL142IiACajiwTD1bCaMlHKdPD9lCXcAiM6qHSPb1+iDH
H80eqOU9NgDZEuQG88T+HL0c2ALC4/yRv7ii+GcLBFUHK0t3mkLZDOhlsKtFgS0xhpv0x8InSLBq
gPX24jPlsz/DBwI4b2QFMDYtvwEy19w4WPArxpvG0pKkRil4jq3f/S20zYBSvKM4zFnlVf4E3dMf
+zd6aPnmr2B08Cx0GOys9ZFnuFs+97SvZSUb7A8elv2yRRTJZwTomWE+aPD97agU3AaOMeZ+Jup5
RhimziWtpzGAv/pmb72hh/T3XcGwgthtdYBVkKBagK/kUlL3z2xXNbBWH29bZ2BLzFD2yePbM+RK
V0B0LMmqT2M70hk0FUdV+zVdTq5R9iKrl3DH7/kvA3TZBEufu0tFCbB3ifhXuEQ4qvi08UP35OGm
kfEwPeltMxFVqJNsNnpxPHhtSlZDDAgALjziYRSQokqDJw16Wh+arx3VTS6y58K8TeFR2D0B9VV4
9yxljEIbgRWoMufKfTcS7t7CJ8wv8cfo+dsnhltTHA5qiBrB/Vgj6YOPZbxVgBJDXoGtPMshNluR
45VNVHokX4sSbcKC830cEqC8q23vC2Iigz17t8rTRyzJbNRsVq8hs8WExjjZmYiTrq5cCHMccYpQ
TnINbGOb5ExyBp+HEwKygmkHnntSLfkSyO1UYfQmz520vSR2L/x6Ah85bRSvyqndpAvNjkghGjlz
m1521YgmEutAn44PTvv00lMDtS9cDL2OeQX6gPoe117H96KE2gckILTJNp7K4HImo7nCNDkP+W+T
Q0u9PhVCeD3ZXt3tde5hsT395NbJSpZM5AlZHv/tCVSTUCWlO2m2IXloc0SzY8G2oIR+HpzuFCqU
su19lVEMOIQQSyEaifE9RqSIvf0ozZNs2L3jXB5S+M82dkloWBBGnEtVYsybo1dJpWbSc/B1u3If
gvmoawhbo/L6W39pB2iw4bo4obeh0LsSbvsGENXZ4kunPbzPypI3wuAO+SnMLDLYD1jpgSC0hDUd
MDMckEEtPwgFySOfsMXR3DBrOb1LSNQyZqeX46XEsI6BaVKgsWMISx2wZIGFPFnL2YkulSahfcd+
0TfLuP06lfotSv9VA3U5JsHtnv3VdWX0Ln9w8ECm/MvAa/L/SO1JnXTYKQGPEPvHE2e+nYE9K1kH
2aKP0VVMOcJDhAUeros6dDGbl4Dsu0FFlK6oiuilYDWpRAIX0s0S1a8rdw44L91grAY88LqRWtD9
0b8KV0NGIKnmAJcrnzCr3rG3+1dYpHwitJ3rtwdMKo8imNMg8DISSqxoGp2sT/PIyfh5qkIhZqux
BsFcrr02ysigxD5Bfmc9q7aMtetl3haNNZnlGe81r88u4ehMzWo6fOuc+4k7ldjFkhLKqCLzu/IT
ozTgvB91WmY2I+QtK2UnDkOKFQ7TavqzOvYYO8hZUxRb8zLVlZHQp/aoB3CLey+ckEpoFO0QZtyA
aha37YANtzOlR0kpHFEKxunUyhwYT4q3cfaDALEw2hvY3j5AXjSysywPl69pkSuNMX0ac8UfrOox
mjhODoBzNVjMqLpC5bUJqSd51YBRM2YnPYusCFHPJI1bURBDdu2hMd28CmImpH3imZAHxPwbFDUO
F7JrUZL5ERiHDIUrMTMuJqQTLEBjUhnfOITR60meX7DokxddZU1fO0YUC/6Ts2JRifEadU2xnZa3
fzXF1TIyN3ugZmQZLKIdryQG3zVi36FMulhoI1aLfoRTZsyx5yK5C+/05vFZR+z+IXtTEhz8hAJd
5evs7OdMAOr+yMiJzao9BPxw0Kt+rAI8XGFJVl10/obozt1foB63QG73QkBlfXE3/wemTHPbkbRA
bW56uL9aGHbbc1dLPK2KdFxNpvBiIb05XDrm1OXbAIVRuPH6d29OaiORtB6DdjJOjbNHEgvtVInp
ifmtBdifZcIXj8lAuMy6H1YZQQ7vb82GNhy+QK9Mh5f3CRzCjo/QzJO7MRNY/iOnOn8ubCDzmTC9
AyXKsrOUUpocmxC+1d3oaCvRh4jn54wTLa6wYQy1qybnIhbnE89mtHfjL2H37lL2XWd7caIjWsqA
+hwAs70Nn19BlkBzpnScOe5SbHcSLzxLiqiFgzrXHEIMUqt3MjOiHTmwdAyWc3XBIAX8TnffWo5S
uppemaxkUor4lusXE9+Y46DSps7ZEgjvuR95ou5dejszdW9IRuUQak/+vWdHndH4WCXFPAMKpKW+
m0AX3PoK5KmA3fUhNEpyXROMT4QwP5TMiRAfuJ2Mh1eLPvDCc/txaQausVJgFPaNIDiQD50WOqtF
804cQj8lu3az+z2Gu9zP4fUyYyxubtgmKkAToPv/Xo/aIyHMcO/n7DjCloRLIkUw1YBZa/OZnWwM
SBkPI5QwMSXki4vPRKV0qvHOCpND36tvt56rglmCeGBIaxEUnTZeAUqD/reKCVOAcFyqxks8xRJ9
9hVZHU1ueOhqhZb/EUkR1CQZ4yi2jsCEEat+aT7+OzTUkZo71e8O0fzLt8uZjp20RzfAkAvxZPV2
0ezXBerEpztnbw1OsX8vdzaDO5QbXNzWBzU48V7rwQ0fXjVgcD4nlGmQEBaeGjCTQA+na5buQxyc
xnaLTTYDq0P4zoZ5JyMOmfS14fQOfOqBAp301t1NiwYOAY+tXzAsfDVI2ECpZ5ZSElCR25ffXbfh
TBd3YRw9+8qjYg9FqgzoNcjO4aLvSUu0xtMTc1tEZmod36xQZV6N1SL+iGk68lJcg1eGXeVLoZJm
WFvng6hh+qpYprDXuJ+ZoXa/7FnLc46Br/Ym0Bz5X31lZuNKDNSzR1Qwb7ncHdqTRp9k4/WYmvHb
EkueBi+97HtvvfFqhdmd0ODvvOBftmWkkG8/TnHhlC6fzaqVA2ZmvTDXJzhQJ/SbpWgnuEEe56Uc
kapIAPVL3h0jdFELFzOcPOLGJdAyds+exI2RpAEArsZacmsyIeANGRJGghwmAbu+IHb6Eg1S61G9
kpr3Vu9h5nwxQirGdfgGVcgBf1TGaN8kVRFWGDt0Ay5XOpYJI5vGvjMh59i2qp5t6/Z0ig77HiG0
aKezG2WatzrNfXSuzYDahX6YjScqZnjHfOmJ7OqKKjeZDvEQxpzoLcFTQsXu+ju3t6zI8b8wtxsT
nJqeToXNAWc9YtN0EWhWAJNVRTYVAalFxSNxWYIGykWNO/1EGw1eXdNBzYMid9b8YVIMV2Hzdk0I
kmlOLclYKRM7HoUfP2ehHvrCYF8rtf742kj2KBRyJ4CHeRUtLnyBWinQIZOMjPsCgfh+S7p/kmsP
GSmv01WDgQkaAR5RVNX7NMIUy8RRNyYlnLKl+gAP7MKUIwdsppAyAfS64A9UAz6B5OauyqzgQ26M
WNnthfHgT9spJOlZ/sKPatCnuToqj3XJQRuiWuvcmfaRGdCWzXjz7jwb8jM3FgHindb/LC795Jhi
ltUlq1jLO9YktzEyXBYanrvqJMhOfLy1ErIDxS2pail3ue7XU1M0kyk83mYhRTSLZnDVJHqTPIlZ
EEZD2GcR/K9PdPCQLGMjSnJodmzedbdMr88byNctTSHgh7zMDQMPeAOfXfQ37MnsWuYIuKuLZqnQ
KHb5j0HysEbpTLA94jU74vBVHNhXQ49crI8lw98LIWxMbpfm/Y8epVwno5wT9wQzmM/I9w76czSD
GFNjyyMcaNly7Couhu6XSun1cRDbKT82mdidbAmjUAcdQsakh/v/F3kbdkI39OkvCP2ypaqphOEu
4RQL7i+mkfXDOHxcD5zlSyOMWnnhvS/tARKe9vU3gEBpUNkd+rMGHU0Hkhp52qE3fE1kJdC4QaIh
MKqGnd/SyXaMY8ZpkCMMyss8byJ9JsuTBf76WcN3IRAH+3eZmsop/SZovkIIqg8FSdR68AwRaT9s
xT5095kHibE9o+heHB0I/mGoV6GXPX6u8unbmBKlJa5PS59Bq3TN+879FTKbwoEKvTXe6BkGGjOY
odMIuIGXhjPzTRx5PWT/SGvwwN9djnBUHiVCnT5h3OMwL0Y8BoQ5JhjAAB4gZORCCTI3URDrxSY+
+Vd+9LZQkHwbkn1HzXWEawsHGN8zJdKD5bEE5lB9KyewrRZYzg0LDpmKRl+s0JoTBLOcx6OQnryM
oONZoMYwYWQJVmgf1zrd60sR9XlFS9l4Ssq1+GS/G4RyVSQSEuhxSNBcADoIo6wx4anxxoe1HlzO
Uj57zjLP4UgBUWL9EC1/LWggF1K63g1qEurqwvOwN2wwjAXBK3cVn7XKYzjGlltwuxkIl9T1sJ93
AIjxR0K5VghImW6a/rvBeVNDmLdpaqQz7yGe2c1rHT5HJEfOoXnD1W3Nvj99xl+hEVXAc8YXylI6
83cVEA8OACWJZ2Rj8dHleSMKpMyRGUltfapnWqsfxcVoeM9tOJmUvEZlR81TCNP6mWjEs61iSAsO
sw6z4sZips8aabkc4cejoCi7Bi57/tpusqO53wh/tkdJAcr2xW6Sp3BTUQXadZaGp0ncsg5mC/8w
LrsS9Yk5LgbQT32h/nEV2x8zVhjTRaZIOz+riLegeJjbvYya15NOdzq07peO8WX2Oj6BZQcJXVw1
yCrqS90E/6qWBbSFSDk0fz47o0vLTp0rVdIPayRe/Ji3vkjw8ooz9kJ+MzDrIMeYPayldpoys3lX
KQM16o0584/x9IV2Jx3Qo3wVsTvqUcvx6168U29iFfW0P6dPkyHuQIS2ED5Ie9k0r0+uoCXyfGUq
VWTlSVovt+c1LVB379T/6z/eVKISP9fNgq6R9MsJwDqemTyC6oOh7sDAluhwkd7eQPwSs0zYhFe7
huFX8a1ZC8kHClUHKp0fnba0KHKxPFmJfaVsuUhIk8VA+YHwYQDu5WMsPrPa5evgWaCv0obHM3oS
HwoK9tyN0h/6NaLRKVYPxFk9Gy4EpHpuyO/LZwwu5tCQzBtJHsw6zZn7YpFgWKw0LOqSC8K5D+dI
2rp57e1cXD4vq1dwcB6LNYd/9Z8nnoCc0pDue0gepx/swZhfwNM12pogqKyyXhjY51J3iIWFtZBC
yMd/rCl+FQ0iUncCFkaEOzTU8x9+QFEwOvYaI0qPEswFKEub81Ub4zQ/DcXiWNuquF+X3xmCLE4k
IJW2KcDAVQBS2VrB28D4rACdz8iVzP/oNLUulz09dL9RKqMd4b1mtvhriDqvCpZBCZFOVplQuomD
GNMTvX0A4cMZ62j+AxHw+MuS4f6uT9jmWzfLv7uPcATF3ySpjwxa9HU486hjiyXvKWgWEzNqByoi
8RfOYNbAnu+vpk5amUbABHb08RYR0NwMltDysQ1anJ83NqtnCPP0Y4qO2JiVVz+FNzFEebfGmQyZ
SCvT9NdQvfRO1DEbtrYw22TOva0TAlweevmoFCrERdIdByTcroiWEnVdzEDbv7m4ehNFxpm+fEyA
T96nvtuf8lEF0xK6P3Cen+cYBGiPjj4jYrKtURDLA/8xz3KYG72DPKLZo0RywTBPXBjE/Zp24Sz7
WDLueYVFLheThAoPH//wIv9q5iAKLixH/AKsjpBjvwDyZg5uDylC+7LnQt3HhsANtDbv3+nInmzG
EE9HXewIg8552rEKmWT1pniwz58RN6bHUOZRtUMutZpM399TQMovQq4li3QRY90Ok5ITn1xbJaMT
BRtYteLdco8m7Ng3QSArXCrkh6lX8/Wa4w7oh15ucOi5LZLo9n7eu4Tirg3A/O/X3Yqtjy8OLG6M
8npQquIYPCBMc/lJJl2Xnmxb9RLUtr0AxO6y8AF6nKuvwSjsEZcQ7gwnr6w7ZwX8auom3Ge9EspG
+TWULORpOyKs4G0SQj7ZN8cGzeDwZDFIvrleozSRlVG3luu3vgt0cQ8oLakFJHc3qt21ORdjy1j7
Ot2fDQU9Fi1aVf90pnxC3TW+GKwKqFSWl1FwEuaqt10n0dk++LLelQkMwmweaTVfqe6T8t3bNC+Y
+1V9nGpmEmq/wrpL3MYyuzWcEd1rf5tMCh0dSCTvAb+HemA3eoPHfDx9WqMDtOOlHbmtzS5Snwc3
qpHVJhFGw24lr0XOWLwkxX8NN+jzX3MI1l6aosbuyxvP8XrP4kYGwv63wTNrcUuO1rsKvSfGew+u
V6h0wmpIUZMcCEnSZg7q/w5gPVWgDCqsWhy3PhRJROGUNfz61984nKUEmlNtsLJn59qp4ZPxMa7O
8N7VhfbAFusdjeuFb3EyoGpDhQRulShCiN8YbSskFEqld++fN3CD9+HmA4An74iDr1XOqROHtuHa
EWQVeTvGorCI5hvsNxZ/z+8OHf1EIsPkEfD6yESLdurKaZcbuVq/VpIQXwReb5HQDvBjVV0pJ5uc
CX28JJrL6mFMNj0R0ZB7xJ6x2N0HmbsiCmo87OUTJiQ3fEoAQKg5V9sDW6xaCxkkz6vgW9apuAlU
B4DpFBfJj/x+f0zy5ustFwPW1M7yP6GWzlB93PVb8HUPqZyQRl0LqY4Ug6XkNORLiAlAAJhOKc8R
yU/t2YO1xEJejsfaMjaYjpsXXfPATp0oeqW5u5TBAkx4eSc8dABA4W4hifJK13F+U5oOrfPmoxJ4
pij9WbNLnls7027uAnCJsz77sVQfxJE2Yni+XIBKLMVef7ah3jcYKkGQ0I/JZsEeY7rlQUuJNgPz
dRguXsgzra7FvTL0SJ2JsQSrYib3wckHHKmqBaDwx2RBaQpRnQ7V5+XE9/2+/RYHmgGU7l0wxYCA
If5Ei9w4/4v9KUOz+nYzLRtWadu7tTuYsM1/SuaZJ0D2sMlGcI8V+SXp51Lve4qtwqRm5DTKEShM
13hIlujqHnEzQY04+1LS5XVw27qyzTSnrIcOuuyefN6xnQ+PPaxbyfh4ss57FF2VsQw+CcZIpNdq
P3wSqUwERT4METfny9W/7Ydlym6CLWPChyuTKnTPzYzXUVFfFQQBbFTpg7k5DMwIWNP4620PWKHV
/yGXd+d4ZTEtUR+GjeHPGO4ZGoJn1CX1sQPTFqfp25iIzHUosu03KFNe4ycBHmpgq2nrgj2PEx7G
JcyWodIIX+55GcKFQfrpsoRt42+Q6Bx3bkDIc3qkkQCKbASMMmRqhsdyZLjfv16GCdkm0yFZkqy8
Bawewd3Cxp+mTEbx8DmDr52hUZVq69+coAm9sh9SEj41P8y7EDJ01swqDODilNl9vNQsco5UknxX
ctL/DMAvJ3kCxF5DytiJLMNBI6bSEOaSnfRTuGX5yuGQXUKpHLrxtHZVLHOXchwDWsXIxoxk5GKv
tIwnGjT5BqCzveFaIMHQgs3xL4k22XI9gIKAdcugF7XGqiEveXIotpSK47hQg+uRH9dkGVYBDVGb
9OAoF6jWoEq/tz5C+DLcaK5puaCgv4AA5gO3imLaXhmcwyQQ19pcixj8uThsU54mns8lcplmIIKr
ZGgDW+UfDf0glmGZcc6fLvOwmpe3AlaoeWWplPvZQ9dJ6Ldpm+845n4y1twcmwQqV5E+0k1nUISc
dnajJqh/d1g+pVF7/t6SItpAUGRRueTEVNU88ZAYAskLqkFVAcp4RoqdyvrcFRe11AAnP8eQ9SeR
kfgh931K/SupzfjPtz8cb0bCLJizfCyXLsNo4r9X8QkwBN8v4RYgcYuInJq+/br8pCN/q95AgtZm
EBrAWWbPdKc28d0embgudJk6ImvzixqE4aS0ksrsylklRwrVFnugHyAWyt7V28fGuYyXHC71n2Mb
VB2/YS/uEppltVkLrxv0kaZMzDbMz31oP2Jnx/eaI5m0b26BQiTIgkeR8ad+6wKIR1nmGfFfCqaL
Om8SB9bmLJt5DNNCUS5UiNVXooGLzVSN7RAPb0WJTbDwpMzQg6l2x3Kp/DVbyiakJykJ5lNU8uW5
0P8Mg+G32B1hpCkUE1R5bo/7O1MSr6yKAiwQ2ZmCv3sFnW/E4zSAVRJw4sjYMxoqMfQ1XOR+hJse
DJ9axr8jQzuazLXQizP91zlrEe3d/8uTRffKjzstldQTYosT81FP1pJS8VzaRnPjdp3trQewoP5R
2Qwcgtpzio36iPTr9n3CGbPb8TNpzxqlLRRmVkpV3L4JWzBwf/7uXkqt8n7ykv4Hy9BuMXxmrtcE
sMh3M9pcFWGMwO5pMT8KDhE+vL1L4DuuKs6DGw2HMFM8DtZoaDN5ykNbrGeYXjNcU9bQYRE7Rn8+
LInqJCHQqJmIUGdKsFLt3IuExpkLLscjH2z9yQsNg6kz8sCc/EkIZzKScAl7G/NEVDuCwmowAaOo
dFUjU1ZRPVcah4JtCbkVuFueGNk/G8RUFLj/N3dNcqqXIb8/0knga/Iht2K+1tRsrVlv7hqJRnx9
Shc0ZmbSSP5QU039Pt0k3gQSPz/1NoZZHBu2n/oaR1IWQi2fILqHORxEKEc7GeJL9IRTjll76Y9w
hgc5ju7fUL8W3ds8Dhv1e///z/5Tw5FK9013cVuG1fF1z60wa96pAw+5iQi5cUtQn8f1wvDiT1Qv
irPULo/QeLRacS62XqUGUGq1RUYutbo7ZbPpONlDoykd0tQL+Mi23mXIP9tKrdU1hKCVlYPB+CKp
FE8wUWu5tj2Qn1iQMvR16zQCK39k+u1m0B4YfogImsNGKobIu+niQ3O9X4/kOg/+pUMo3jAl3yIp
Jp6yIMkM7P6fLYI38HHWYlhRxipUr/7yV5NNIIblOsM723S+08uq6XhVGUo4livC83RHxNGmhnNn
46mSqu8zbVO3HOk1zfwEPuTCTpVnDVekAFX7c4ZTF/N9mOh6pA/pKty+gcLVsFbF1XgT7lxOduFl
TbWV0PpYvhMTiy3RzKPPVCk0aG71bWwksBjJY+ePFJNtWfmHBuvAgJufMuadj6BqXQXZjMvTJjdv
SbwSwuEd8tupJVrD0y7u+yfI8UlRIE8ftCykONv7wrCzmOXDECOOCFuwpAaZUQmALTqZoZyfZV5+
QTTVLfbnqxJvsLE0T2hoisXNdnjAjjf3ZmNZWjZWGrhI2MZIL59oQPHP+1QmID9SvIEBahQWN2ew
I7EdUpeevWkGP7qhNH8FV+L9kLqpaSBiGAmwHXe4cmwHf9frzHKRRU8G9WiGUuJdm1n5WqaVbEDN
/VPiuzWQot1qNFscTTiWtbbS9uFXH9C5Z+XHnNDvGgnbPQNqcoX6/uqaKo1oATBhB8K1EipXuYJc
OGWlWSRKOJZTkKZjc+v9B7i0wYEmUxCRwIHkSWGKyzxEsbgU5itytV7i7G+1MdTfR7025Gq8Z3j8
Q/DVnMBH9CXEvXlfIP+ygUvF/OwPLaEIDGSxMDGeh+/US1XAkvJuGq0mt2mB8KremuUxbVPSm/cn
K5RT2wcnZO+cmTXaKamIGcuy+Mr3/ifmSLQuwb8bhjR+3B0TNFQr8bDRZBThqkQSG/gMlAI26TVO
zKiRKNcSyOLAA3PhrYLnGjUcJx4EUL+U7eaoDx1hvohB79zZjCks9zIvX546g/N4B6vx6EFas4Tl
SDSKrQhBIalQxH8bAHOdFpYgmzUWnS60vzs03TK0I8ljdBeYCt61BRolmVjrQfdYf66X7jPvUA7L
bcgpM+t9Jdvbc3oRFGqdqoopjk/fkAwc44aqnTbL2a2AHIfpW7Kd5rlkmJHtXskuZP9Omlsqzvu5
5rSQON7U0a6zKiBFM8KzwvXwu+a3yMJbs4g1q8fgn7pZuXoj9MX+CvmLtuz3LOQNkT2YsOrkk5Nz
mjVV+IcgkKlQ9GF42T2EYatMwJZMmT3/rIIfNh8qUl91/NOSf8yXSLRLOK7rU63ZrNMXZB0t8aUU
/LNeb0fTouddy4YwEuZOzdiUVIZY2asyO/X7FP90lRTdU8hYmeZ0gXV1O54BZqnZeFPtvQC1r1pO
X7DJWKjsnXlYkPKSwORBCFHpAyw53yETlCQIxTfSVKxJ0eL7zspw8nfcrycAcIT+w9DUzyHMPmDM
BuqXXTFO4uCC6HjagZ8+UgXC9jHIorhfPfNwjctt2DtfPvaDhWwxWrgTJVyooQtSCwLzv/W0I3Ay
uTa/mWqDXIKHDmAGpKV554bMCUjWs4a/ClJy495DAJ1k1R2bgnLXHD6T+RRxDwTJYpGfCq8gT7/K
8L2/6XmxdYNbrWfk1sQg8+NShCIf3JfSynVB+0mOragqj4yqHzaSntBrgrQ2XYIPikRmMX/QiutA
VH1UtfE8H1UB53mXFo5nSTuC0Ait8ugPS9ovl+X40v59/rXsibtw4v4CcfLHCF3qfvfiML3r08vT
E29DimgdwZQO4KWwBENBieeao9sbakpvmWjVvcdHFvksPElbGEabWMHp7EtNL5O2HxhkN3o1859q
T09YimvwI4czAF0HK4tNr+qQInOutr8XPre/tU0PsHlsAr0WSqSv2vCppTgGOA6ypmyBaJb1aKx2
hbQrOA6f1pi4o42wHVrmLe4lTfDiBIi0YGFlGIinz+1bkLE/VJaW5g3w8YJQ4hf9BNbL9Fmt0S0t
vbj0S1E5rdatCsaRot+eLabBKBubTKHINZRX5VbvfpUx6o3hZsmu6QfSn7GnO881h5UK+7npPOpD
NwlMNAETZdHKmfvc7XjHo5m6lKfTRxQX2HlgwzT7t30hxThy5AvBE9T6aMxd9WN+OAYfKc5D4ULc
dAyWPhBkzQY1+IZZAXU7p2C7FlB7oxDr1EsHs+W/IdLIvOGGkZC3ZJDokwYZipnBowmwC3U61euW
eiiN8wtc6KcQXHuBcg/4lu9+xGo9YZQFC2DyW8/KXd6s4PZUdtp/oNTBotmdG/kui8czR8+huO2+
nbhD0liZwGAK7bO9YYwuL0Em+dFz6akQ5rOyzkeOrF0lwOqaaKwPRVHICAT54sJwXW4oxMNYDfyz
Al4jcRPtgQ8xWMpmlfsylZNWuOzL98N8dxroCfIyc7pMcGgBWne90ea6n1dfTufFZ02x1sFacLEx
19sgAgfvHfqWm9V/UrPvUXaHKcX2FPMseTreINx4CHBA2drhVX5t3niOD81Erev/lMoN5efLTaZM
ZZuFtlePzaM291XMfx2Goyq0xI9OfuIkiolr61Z4geCJ7rVRPCuvnHbRiP/dyOHwpoUUDVizkqbg
Hr4SUp0d4vrOea4tkNGOfJyyLvxi87817F84DQ5cOrEL3TYIrPKI8vQjQVOetXKIy5yXb0Otc+bV
j2ly06gmQaqrbMutBpU0+9hn+xbzJJPDfEgJNxKlIgw3XsL1m/sUU3lJmxGkkwhvUsRkH5CiLjOj
1l+mcJIymL6djZMn5mypa9/NYxP8/VMQRJK42FPD13vsGBGJckDl9FfQAyrMdHLY0gBs3WmlwehG
OnjxWmQRzS12T4+oy6cr6v9cbAQecG/cCwYlrTsuLr4RZUBUPlhPHgHFx/CrU0buFTA3kkH3gI5a
su43YLI2LMd+99TJ5Q3kZGLSrlDWb7BCtfI02arWy80y426vid/XhuvE6enl2g5zsM/egzvply8e
4rOJBbB0D9RkeBDJ3bpHqtOnCcxoxY7egyDyn7UnBhD70c7AO1TOWGSGiNZCABPrhKzGF9GPXq6/
UvkA1JUmy7Iq3mj5to5Fla7IZwNuXdkp7R+2ltzOyoEtAKilZ3QUlN3VBkqur/GwaGak/zjpLswm
1GVOeXgIj40qGlGyhuMEqD9fOSKOe4vzbbyvHN3kCKN4xy3/XaDAfbk7TsAoRhL9dFM0tJzjZC+f
zyAUS1ofyfCPd9sEPbE5drQe51bVHfd2bgUBDbRiXkY6qhdsR6gmwXDZpD1WxTDwdD2RNRR27dIG
eAwdjJScPAmTZtOUWNqjakYkTx5kspWimepnj80pbEDfh2K9fk0NZjPhtPpskGlsFDFu1fiZnliG
eeJfMV35vpsj7Q+Jt1erAzCVPiX381+Yd7XKMG52Yq1YTJZfHYllDQT62wmprs9fEXiD3rcI4m9h
lcS6kQHqlZ0oRns6HBBF0+suflHtN6efpneNhoFMZsCFDzfJX0SWdlI+czZiVoMh2WdB6j5AQtGA
D9zuKwkCXZYDgew489Vt7iWXpGEF+gDfU4kCIVb95WISf+kAaI3kRXmkP2/LGsM+YjqMg4/kbOFs
nGHgwuGCx5CHjVPfHksluBVkL5XVpzOTFLZiq5a1n47smPWilPGJY9K7BQakPLc79nfABjrZNmlC
Rf1cE+YYi8sKFcfSLDdTJ9epAajVuekbbupVi2269ltp3Et38ZefG5Y7ugdstXtdIglr2SYUiV4H
v0ckzLtOcWV9qzBT+ohby8w8vPvotTw0BfyMv+4wdYFvfUcAdsKoobKf3809Q2nZMXthRRGZ6B4M
V3pIXY2BiGBo5gf8P9xaMVau2x6frHNLDbeCnaFrVPci3sNXPMYxVp1muj5dwi1T4dMj7Z92i0sW
Tg+lkQVnz6Jm1fccGhqpDUHpy2OHdx6CpvKRogQeXGGz0dHAqgpEqt+6MpM8rbe6WfuHTE/g8FO3
/wCJz7VDx3JhthDwbvTDTkcG3c6hTimpHDLz8wUvPX5Jxv36fqFj3ORX6MoAqAFY3SqZrLAu3Ybd
DPppvPOscMPgSAymnsv30Dp461M8emJodNkO4UecTS6zDryjTzz8pWyZ5o/xtklvCGvQXLVYy+h9
02aF8rcdn4InkiAfcl1v3r2JsVK2IrdF5KcHyELKJP6YG+M7ss+K/7Y9NiSrBrlLfzp26FUB5dVn
7zlvJ9cceYU49GRCJrqwSfSjcPMxgqsyttVCemu+XYaYLPZvWzhue8P9PXN1IR7NBt4UfWomhgNH
vLnS50gA/S12TIU7XxHBnvVn1Qe9VwiuVJYDYBFxu4GEgfNOR4J6wVJt3fbgUfXcx82mmrOmzcSM
QDfnvgoQ8XX/lUnF4X+gKsQzparVh7vx2OIPw1+xKIStltAoelZ8PTXqrVgfGT/l5sFenLCH6fCm
iOznhoPlYoMrcdqsR3JCsrS09XNjF2sAhJGbq+uwWpuVo6rNCIYR3N0HQYc5n6pYrUKAeYOFI+6P
8xYtWEFJoAS+90U9gDJ8Zb6qmynCAN38+HommlWcsIZ8KSslnM9hZ+A3ATW1tt+diIhZft45MAVb
XqNhThdWlTClJTsCgCjhYUTBPD6kk7zUdOP63rC9JDdYa3dWrZUwp6bFlF3v0OFjBYqQRXZOpkfN
NWnanyCqLSQiMHJTe/Nx/6lwGd8ANel6oKqdHAnwXQWmbRkmymnW6Nm4z02DTEgmYksTQxdtUPUz
wBOlWOI8fqFw70l59tA3/xwdo1gHoGgzTsMVxYZlfsD8YzBQOQMZCmkieg2CkjKwA2arQ655D0/R
d4VbggRmPy558vCKI4ZBSitZw6/dCxwXc+Tchyum9xMv0FXFFTs55YKQtu86nBX1LVgUm8mOfftY
Z0a+VD1I5fj8lEFp7RgygznNHYfzrgZHpz4y1z6CORK4h1034TabqW/KvRSk+uKCR2yOqJ2FrZCF
xciptpmhac0dF9QCGJQFGb96MN1rjpk5htEozk+E2aFelRQB4pq0Iymx5gFMp5hne4B3YJRwIF9m
nnvvZwxWcA6TId0GipaOM2kNCUjNXsp/2iGADzlxgqAT4YHSLImXzD8YpOQe0hzIzihZUfortXKn
0toLmiV+qtVlKBo7tdPut1DRcF+uOZMRE037WGhSTZC2MJDcvuMWU8QnlVJt+qiR7GtS0rWh8NMx
+u0N/DquCds0bSjjuUmJLgYB3qm8JXzvZ6kthigOJqEjPQSLDN8bD+yH5bzyAJD2mBxj+Agd0QM/
hf04q1j2CHPeG15HYoeII6qRF/RFJ5F5z0adHP5DzSNsBKafdICatO3I964cGVPXiCkvqKfXtfE7
31r7Ltlyal20GvrzhkGG1cpz6RczkD+0uoWf/t8QawntyN2LMssbcW7VxKQbcJU1vWDLD+NqeUFw
o+VJFt3GZ/9UAJiZh0ixSvieduU1PcOKO0KyZ2E12Hpp1jZvFAFBWwRTtmJyeytV8DxZn6L/3AkS
7LkcbP/s2WpSSqEPAVDq4qRCJLLKV0HKaRbLds3VumV1eovrQO1PjSfeXjOtvyghTb2vYfz5nOOR
kaLa3WIHg+hE1aK1DmmXkGarLWs+xBjQBCDX2Tml8NVqQe3Q8f+7mwDdHDhPGOH1sBGH8je81eL0
Ng9J04iRj9kLCnb1lz93tJLS6sku0rcTwrcLoPiO4wiCQPz7YdhH7sBEjPnRbuVd82wJz8gyNN3r
tpnmnYPeqVKuB7eTmSNlIjqTqQbvx9Ie5T5YIoZ5omyt5gJDbPvbMBjSYhy6D1fSHlnwHT8WMgkF
4uj/b2tdleurUDOX60g8nubEziS54fv7a7kj7v21pC9IUkItE6a8RIpDgZLnDyidOA6sglqnJpQ1
TXtAiIeXJLJVxOcMRd+yXKhig7srC7z+x47w9dR8BELLNMkPG/G7LilJvgtzhGjzDDth4oLp60r4
HHT9/fugeyWgHxfe5E+KL94zuFGrHLqj6pQ1m4U8AxUjMUTlwc2S9o6AzgfP/4Gx3wDGvsQiXbne
mD+u1SgB9hNOLYxh0G5oNcFsfSeIV24McSAWRb6BqVmi/uRijp22SorbNyYPWn19Y8c56bu5DFZy
AYjXat5zfeoxavlp/njQ2KpujqJd12vlK2ZCch/NszSRyn8vnQQmSv5bINg0sCSXZaPV8K7a2SiC
/hRsyOLYdHy7jjm0MLGC8Z0HNOKGoKQoIzWSFZ+TZP+rG1G7QYqacUkOhHhzPWJN0xt0o4OkekJg
BNm0svD8L81Xpef2SJadGyUFKiKWDKI61Opb09jpOdwx0hh2vmekUQOBNrEgaR+PCLWePfTTfNSh
gsFO5pPt5CkUIEYi5J+9efi01ZjKWvZaXilFb5uHEyuf7FMJRVFixjZDcy+xLwYiuTF86EaYP3Dd
L3/D/tdy24ltF/TBFXoe00AMiaHSwOocQ1OaaAtSDj+OK4yX6DUv21wG0OFT9rMOehPw8YvH4IR2
X4D00k2GanE9Q9yjXLkHB1P/fi9GWkpMCT/5DtrYkQQWWZO5K4OB3MIMruXrOzQ1X+lLZu+WQv8F
Y0HFVnltqrmHgbbA2dtQA9Gtqs1vuTcfFHrl4URSfRCgPiRVCZf0f9Vi2AETUTKOA3sqPpbUxuqN
o28TAv8VdtG66/Cg5sGLM0Q3kdkearPNc3Mm1QN9/KCSorEIRUt5dUMT/gFxCDKatwK8UNhy2GrW
zA1STbZsavH9z1c4taiTgiTSPR/hbHf+b0lHkXiwveM6+47znrxOPDjQh6ttz1gd9uFTPLhqSPyp
GY/ixc6lsQI07GZikCYQx75iFi9cnGkZJLZZ44leMG7FBV2mY52sb8MH3umtb1r/VnIGBF6qDeXu
qEs1yI3/aCePxmlsjddWaM6MrmEhSiCJ/RlAx0iCpCmv5H//mqjdrdTfLRsTaHupLghQgz7ok8Gt
LydAOhFixk1N40FijUr0hxGv0lRM9W0ndZvtEO0ni785XmgjF1rUqSD2QHnuMx6jCVS7TnbBwBqX
lZG0HgYY2W18eLx+GsGxuT6q/CbXYfKgAE2lDS9BdtV8XvAwLU28iaIkpninYxCXqIF5heE4RhSz
YsUIOUWKirJq3kQsSohJ6Ert5H4mpmldCqYQ8iPdy9xxSRt/Rhpj9/opb6od1Ztv3CAu3Jmjy18w
DzL57+u+8i/ihIgNq1aAtTR4rgMYsRfBF4Q3tOj/ORCnzPO5DeZt9U0UA2HJkC0MFKqgC8bpkMHP
HuFvSOL7aPF8SysNM1XdhhQtcs3WGjSCfbnbccdVEH05qxHiu1x38N7OmStby+ZESAgxPyg0EE7r
osCm5R2wiGEfPyGWO8ptLP/JyQS+qPfia6lwgvXMCxW4CfnOYS2jsV+SePOF4gIFdbqhGmMdHPuU
hdLbGwA9Ty934Fb8nA+a4BI20wcZ1XGiH3uhPa2L933v/hUMlProwyLOO+l84o6AI5o6ED/YlXsx
zgTRJPnUgV/iqfxdTjg45RdjE3yPT+cNO/fx6GiAEUhj488i+nX4oYPzxi7AszdtkcNH793s79Bh
+xEmB7QMup0swTl/5KWnk9jfU54aXrw+gJzbVM4UQlAXIygPwAsx9mzvxDbIPzb9ucKSMeGLUqCp
bzLbQsNfiMWvGYNQqQO4Pvcuq10xYVFWpWOTAiW5T3zJlLVM2cdDAIOhkyqsYUJ8g2eG0CAavDHq
+yVy6+ckE2TfKqWGBIwilj6MhJpeZ75o7vdZh9AClzN7hRblhzSHY0zx9QL9xyTvX9h+DyFylYD6
eHf3OWlUZ6FVvhh1dM20veZc1ZTaQkhICgu+7b9ruEuHKh7C+rs24Q8C67r8FJoszs/nJVICGDRk
+YKgTdCkOJyDsY8rXXYpwNXRBUieqDo13Ddz6Y5+JMaR97Z0KNCoxo5KQoqrVlNX/dCCxVwCbKjd
tJnBf+BcrO8ok3elIPhfwFF4NaBhmORc7JrqkkQywkaXEUwf8UZk7D3TDkY306Yj6OXNtp8cUhay
oZqYpduLecfrHic7NHk3BO7lBWqMeXMPWBOKOkiSbYYkEUvi5ip9eBQvfr99tTQdd9zlx7F6V3I/
P14y0xJrkGZ7ugN3jKAGGWNrBXm/XnXrzqIpPuRTzcE3VTn5RsODje/ODCy50HduM0IsFs30wSDq
/z+W4SyaQ6mBKPgHV2M/9S3SAq3l0NXNEvFndqN5sZtKnpPPK7DR2fp9AL8r9NI1OOUf3qsVLkVX
0atqVt9nv5cTCn4VP5qlgxS2XeEPXTPiomqwoPv6RJUHjRFLKNlELBkJumXdwmnAxdR8GviwT4Yj
nM8MYqgMBBtiY6/XIPMvCkLCkddXwRzgI1qzCqLA9k1Uz9eYGVmlks7fnkY4pg2Yku4SCV4Saz8I
hr/Vfk05GwHES0IEaUj3Dmz7x6KF1pWNCzkS+Nf5VfD51gwB277QoxXAjyYU12dSqULgPnMtFO9u
mm2FWUPwLnPwSWmtVRBaDNk7atSlBxqRfaKLz7PpHRRXZn88HbZUKBHRUYh+DE4PT2IIqgG7+d6j
zYZ/5W9JJmbSS405WUUowCoAqjbnUgSJqSvvqeLxZvfe+IWnmI5oa5lUAvf8yEdN8jSiFcrr8HJX
2oUaLKAXCs2GaGasqkFZvbC9D8jaQ+xUy7RU/OY5IkA+QFd7RbgpgQeBZU1Q9EFbjmBaYcLBR0zw
J6opHUk926vAvK6tjl57zmavk6Ict0vCnBArnqDKOm2XiFDmEHswxc3eBloA7CXeUbz0+ysz/WJ3
EnIMpGI453Go6OEv0VZZLm2tF6RxoGbb8l+if26iYk82WqKDV0SO5zxzXjw0/bV9hvO7iRmkVRZY
uZE1GlVaID0ZwfscA6sqhMqgUUOOlwqH4b5QSYUNr8U+X6j7NNmLVFoEHNIGhvfc75CjVzM90lD7
WzeM1Zfb/pPOm2c55F3vFyYCPfFBZPSXvSWfaZQh7BoMfJkHtF47CGq7BZDcE4a60SJg4VaA7T2k
i6pY9dd6AkZy243sKk+LcwIBK17FUXyLr2jB+2vPcLAvBjw8rmXqh1byiW8jNuUc6jQwlQRCq8N0
DFxS1NEnFzXsaPzJPpyu4R6w81TjHer22kg0CzhF7aXXwrXQbQdAWg7FEvfdDoCm8krtbePx8QWK
PrM7iXHwdn2FeCgQLmtJ9J/6LSGiAGQfWBm5FfKBTNirHi2RGwS2bvqLlzi7+xMLXwJ09L0snp43
bw9JnAsVYjEwmSEbOAZdew3kZh2kpOZA/te4kbVvHsXLMutwJrSrJZ1zN8JNhCALrJY5iu9tNZQa
3Njj0qcKUo5jNecvrmSCzA7Q9KEQ6+tGcuFnfrME03YJ1fF9Ts1bmev9BtL5/SLbBaXZGCTXsInd
6P9HBaD5e+7NiIGpXQztSUyf3s8lG4znLAIwEb6aPJjgLVJbHM+bdUjm4xbAAfSAx2VmOuNmILZx
VXbQp4r/bM2VX48oMx4qosBvP4bPxGr/C99aQYVoUjGAZhEBCIlJD8Cw0SiAP81zInBvG2b8WYyM
gDqaj0V66jm8H4ZT0khfGbk8vrtTwmajPUDHfBK4uRSw91Cx4bz5cShdEocKZX4KqUdwE303A0rK
7stE81jZmokuGfCAI9EOEJStHt21Jv0UhEHDYfKTAoO1tQ0aOYie3yP0mSLDZmOKioYXsc8rrmrJ
L9A1/uOopXoaXX8iGKZHZF5mfr3V4PKUG/j9w9nq35V+uLb7iCev9q/QSIokKQbnwBfu39etFcbq
38IVE3UZiXMCokUHo3J3VcMGLKCp6ynB4xR8idGuLeml6Jpw3pOIitxcP7XH3lDWeh85GHJrEmRw
lk9+Iiz5z6QXBjtPgVBTtAIRkv94KJ/22AomgdyznQaToRG9KkEMMFHG+597siDYhJFLkCfNzkt9
38L1AIM3d++l7hN+3qY6oP2J3F4fENaM0G37hRL8iNt2GqNWO1UT21pHWwdQCdGdyy+Pi176XLYo
qLGQtDTG+ptK60OZQNOj13dWQNl1G0+kluFGOyzPfWC+4DU271vtJ4Xkm9mEuphyyKDFnaiHm3rm
pmuypqFAvcgtP8WiIS4hC+GLmrBJEtaJjBek6mID2WTteBqQcwRsY0GgyjxHCfzyP+QlvASHDMcJ
+yA9ROhFDgItyI2wlen67/7vJKRK4t6oFrYk9GARRJi5c8aNcJO+7Y6cJaL8BlLLLil2qOhhyQeP
uKPG4KB6pc9GgEff7MnG3uodqpszxvWhbfQbB3fBy8TYXfDmgOQP9EjZg9EO2kPRMnTms7anruZH
EFz8Mxx+e8MKjvUL8Cwgx1TYzeRcw+0qGO78ZT3No81HAJAfSyiUjQWoPclurAZIMkltT8oS51nY
Qud2yGpIrLF/bkYk9C77aJsyTeYSgYWfYxGhkj16LyXtWSXr72JihGd3ZeJeCWsSyKYfjQSEA4w8
fMjncjXOFvbE1qE64tYKudiPvYrRtyayDnDDh9PtwGlhMxOZecXA0D5JMFHV54tdk4uxgB2q9gpu
3NYjQbcSy3ZnjvGbLj/dgD+lQwJYKHPm/WEShe8C8VShW3GkJDX30nfSefs+7/R18Hz1ok4OVet2
G0AACyXFddRu/IJfhlPwArEsddXNeZA28HWqsdOme/JsfDVHPT6kFnKdw9Yfr6HHCp1t9PLTdXF6
nPkUz2rMLJu7l4nT/0q2u9RloGJKIWc40aho78QazhaVAEjP6D9x2GC3QDhz0f4Iwl16BdrVTf72
89xe63CvWUX69xjtU8OHP/Tyd2PeaeVCS53MOPnn4P4TNUtkasXGZsGgV0I0DYE1KS8ELJdaLC/d
g7OJKl+UvELLkS7nNzIhiiYbAFDrx8a/Rxycj2Pv55+5cy/xq8GgwgTCotkhKjeIcTv5Agk3eXtu
QLC+nc2K3w0r0r26HoWGbVfDpMiSGxIOih2uzKw/F4CV5CgXlSJExpvMGM44+c8IWCAL6974uuro
tnOvlfUl8S7EQQeAXrtu9la0ZPcw1Mxqo/SScp9y/82XT4EkiAsa6bmYYIN/E8YXkOFCuFBkEkZ+
tfyOyPbdCt0RbJtuuwPKlo/m4mm6hWdCP61WtgJdINhjS5BVpHv+bQfJqat0ZbtDMD9PGwa89Fpt
gSEL625TuBXX3X/eGdi37jSnzmLQRU8cxdYQ8HBdVQKjIvkdg4mxCuRXqISdGcsXX9neYBDdV38u
dfeBkJRR2K5BFM7zpruk1dOc/diI2niuvaTe3YiatWoU9MulBgfGcXZY1TIDrcLH+ssDGmWh3a1D
afE5H/sUFTABofumujGOt0zwIgJR8BSSd2M5Hl4EXtfeVseFWJMeH2GtkxAx0TAaqRYN9UVjg7Nd
svct/tgc+SdfF2PHxoXjxrldTgaZ/bqwJLO2PMmLMIy3PtnPKnoPpNDfogReWI2Z0x6HQ9wb1jXj
2VOTuJZ4DhG6c+hixJYSY/BD/VlJFcC5RVFS1uuhhQDC8cEB8mlAZK6tHaYNZm4ctMY5jjIjKnZd
mJ3ngAGnKcDkwSmJD4DHsucw+CZdH8AbSAT7C/p8MePOpwu9ZMFxyFVedt9ItvfaMXi+4AFonHHU
rL4kYTdLC91w82n2U4Tmwm4t/BGVbdlhFKybUu2ODsc41prD1kRZMyRWGVCvri5y4DdScb9PB2QJ
g7KeOBDDnbMNCEjSqQOaFxIptf8k34UbYkOI6lv99ByviubX3m7iMZo0Sw1PpfDzkqVBMH9nYlr5
tWve/BAEMDXAtlQT6h3BI99lOMxrGGKVqNp0WI3j/ULpbFPc42Wc3SNI9SSk++adNyNuyYH7UQwy
o8GDTwW8lcDcpL7c+AAiclgGOnWqSDYyXvYmiHBkLLuD0pWnLlE0+DaYfbyMsH8ON9HHbbZ9u/8c
fHt/0Gs4jV75Zt31o1FYAEQbjEItaaLKN5hUactw83ZsLhXl/mOzQLTbA8geh+jFVA9nsrISprKU
n7LFHGopShkbSoHv5PK+4yYbJF10Lx4xj3XC0zzq7Rv76aIIMD/QvYaRcxKWNMtbxKPiKhSxKCJ2
rowtMG5VFHIsBjUz+QbIDKozhcec25DhV5Oe9Z8xRAm1T51FAz/JT3rp5w8cI6xC5uAS/k9DQgUH
kwVZrDYo5bT/PTkql5KaDyt2Wrcvb3Jsh3CiXdr4gTcZuYDjrbfV2HYuY8MqY3yc/A3QywGsgZxR
vYQUpgAMA/S+Bz6bEnibDckxc4jG/0f9gYd0bcwNW0gY0620vFxEYbGkTbfjQCQcYpHB+8XNz3ZQ
2CggRLRxm3yktetxRcQw52SYExgKYkI5hYjqsK5Ad0EbZfektm7Ru+TgHWd1oP1TX2JjPe4NmEvJ
vlLt+VCXQyWhbJEQMKrOqOWuryuxq1hqI/QXEldglw+S6GB7eXgUuW0eodSrx5/kHChMWq8iFlY6
TIEfj9XFHHs921i6vD30Go3mkjR/dF6PIohGdgp7p4AxRdIjg6gQUXe0kVrblrM/85p+Xf2wMS94
mJGlgUx5Kw2/0yfRP8qQv/QkSLbaifKI9de/58zrvXGyegVfv+3mwZez03emDKfSNKJt3lACO7WD
jkQK4X0hXuM6rolJwbHmPlJ15GcVMc3HReiVSkLRqMkqZx33OLCOh2qo4fOfgGRupagkX6ex3eET
GXe6Yr2Z4LqnJFe/O+TtGXnNBswGIlz+A4pgH4GSle3VxUtVtxBAoVQfJd5KUZWC25UL8ddo8Eke
DAbEMZu+yMsxhopodwMjBZcIUevuNmli3l+coBH5R6xsKqb/bemJnE6sOGhChPtIlaSVib1qGEqC
gZNc9WnbP8KTrrCyLlcLI/RchkKXb/dtBXE0+YrfJ7ER5qCyRM33eOEWQ5vRa4G2uUrKBHGxPIzN
4Gk0dfNwSM911CnC6aDV3y6blcMsnBlCAqWDSmlygvikroy1SqA2iZkvvziotCOZz/q1ODcLm9Hq
Gwwm64SYTHOQ2bu8JQYRkpXXbpngIrEn4VOUMNJcGHXweeElaShyPmsqncOjAIHEw8KzMqvCmY69
NtmPh4h23wth4EBYtACYICt+fYxH8oATACiYScIGogEe7zQhu14Re/RKV2Oua367As2m+giv5MO4
DH4OJXhLYkbYaMchnXn5VE935fo82BReHkq1/foB2PuAgYwfbhNJcvMGa2RjnHIaprpFOOIFznC/
4Xk+cq2MnMMLx/iclYHaNcERaZ+svYjCe8B4JTP9FRLLzDspw+quuCATej9AvgKQRWMSSgVMdUQG
4pTueXuohmGUiXpmM4W5uH12HPAtOP0x0sFAoIWgkQEz92HhBGI9vZCQattxlIcLpY5uIn/yMT2w
WyY5a+8jBwDWPyzm0mIza1jfhpjmNVMG9cm6/omZ3SFcG0/4V3iRulz0gF2D9eCcTKoikzuY2UlB
5hAY7pEQ5N1WKizSjsSohRJIvsbbtMC8qLWC/r0ubCdDMj1BMDX+LKo4SXPCk+ezNWXe+DDDRkg9
7uIFmAJWO1CY19mOrRNYbPGAYwQ/gEf3hxYDRMat4sXg8dDo9XHrVOtNP2Wb/H8SKzeJP0JhdaF+
9rG3m+NDmuVSkkIrK+qlHSLSIjgWcBbrvGDaQ3005fIIcyg6RQlQ9nF4CSMHiGKY8sotvlytWivT
eptQuAP4WTRbWNM83ybnq08L1G9P+OkZzzmNDCSBJg1h5McjVsMPfDz2csG8q7gRfErMwlG9bFxF
pbYdnTRszW+yKZoR+ag30npNMxmHj+3Mpg0jBbo4/CyuO/Fh79mylAWZJJhXAZej7LrgV6KmKlf4
8qBWyGhUh1pkD90sTWy4OhE03/ZbDkoeoDKriSEWZ3LO71MqU7Fi6C2wWgOAELiAHngmmgujzJvB
G3Yh4FjW+3V5crpg5HlqZdI+fqxx3leWihTXpArF+jnFDGrjZGZgRi3PmKFC/vyj9cU36hfjsTc/
f1RRG3tGa23t+SjZTE4+j6c0mPAxNiJWQh+SOKMlSJodefoT/dI2AuLzmRhknFZfRcV/2JC+ekXf
GZtfJde3cp+1XdxkZ7NF/7xpa0GUAEADqQy2Dd+MgBVgyKcLA8GWlNLxu+kdz+0AlLOTbGKZHH5+
9m6kJbsu0IXhdqqI9Lk3k/FpObtsi12uZ2aZbxShxxw5ovzCZHFY7RoJ3KuEGIJtQ7z/CuRdcXie
qhvAzobrERc+n7inNAs8V89bKTHvd1voiRlzpyn8g5ogVlR8iPUsrQOSKVKj5v1XgVkl+4ph3q9s
PRRiXQ08DZCKbqmy/rcpZ+lLNcJtK10XwhVHHFFFdMKyKnDlp5YJkVeaUTImHM3pzViRAT6w/2a/
CYsBweHBtSyUsg6RWr3lsmpJ3xQ7oB/KPm53linWKEKTFMipmP6H1THJPD6YGzabNw/FjxJgkwsr
qQoU4UVKPqVuYnCUn1CEDfPLLa7eXbhjOETHV36AZstMxMckz3tquX8xvgDc21aGVGSOHpuFCaaf
WvLEWzFwD1w3FGrlnbrkPvVfFxC5uOse8LfodBAhJOyX5SnCCIx0SuNoXEwBbwNZmIt7TSBVeKrO
mM8jr2l35MNA1Rb6+h/HqD7Svuf2O3+yJ5pGAgW4+K0YlrcmqbSCxxu3kSWvD6Q+HfHAkGsraV1l
5LqGPkQcmlnMO+McjiexWPCdCbSQSScKmb0yukRxvTIgOq1renBpUYgDS4X63Hq7MDuBKbJOxhwD
GeFguJNJM6QqpCcMo+Yynp26yy0F/XR/rYWI/a0UZrNar3AvxwN90ycoDZetapriUJCCQwtGjV+A
Jo/9e0SgRQonc5MjEiinEHfvBiqk1X6x4gfBQoPWAWWY5CZ5NVmUT8sXbTLVnJrzf+lFyQxuCcft
OpqbLT95ttB1+MBDsbsBjsNhsaJ/yGTDOgCTiSgLN3pXFN7XKOwlBNvT1tAbztnwXnWOQRJajoxC
QbmNlJHzbvgEwMR812iO93CS/4b3xSysjkYbq0vOu1gVjVqEVW3MU71OOA/uJUYDsaXEhFy07qoC
ErpH8tKhj6Uo0tvNcd1qlC61FaqvJD0FlL7pg3ffwW+1flka1TOz2oiAX0iEZce+HNa0w96l8RlB
EsMu0rn+ZeHlqcNyMBYZtVCRhiAWCnI5GYm76Fr3mQX4h9QKaEaSUHIU2nG1zpounsyqzpBF8wIU
a10FNB7GbhvleL68mxG27P+XS0jnTHXPtAbHE8acRTth54Sv5fh6fuwdRZ1DJ8My+83WuJi+uqN/
md1U8RfH2/xj930QjpbGRpOIzzfA9PWi1k3jo3nciju0jlLy5AL47BlRfpH9mtiAyVLA6guVdysh
FHdQ1upB4x94TXAeNruSC58w5M76l+fZsKCVct3qWo5B2oi5EsGBIijk3DxKqsXpkcqIN4Udk4of
Siax6LzrEBGHunGhvunh1nvcYut55ROsGQ7tL8S9DNOQPqQR45UAc0To3w479G2Cya3sp4W4PvRZ
2SqcnRnKKvyi+oyFBbSVreYlbrR/6N8ldNjamFUp+LIsUb3vB4Uxd88TFo7B7mZdUtRTSgKxKmaV
V5akpVItrvRJcVFm7rIA+xl5+8ooaorxh4DQeRArQIOKctkv9MVOb9E5w8Y28yTHTlvZQ6I7l28h
XUsfm2cM8sxypTuBZRQuhHFR0wUVc1ySxDqNCvT21U99Zup1iG6Tgyd5X0J/vmqmilBV63a01KwE
dv/gDZ15fZenB0h3/o6VCTbnEyb3GX5B5TkayyEJ2V+K1VBbd2ZQIEw25nGCtbbONbHyJSNq8C9n
pIArxzc5MAOtbpbAVfJjVuh424F4OFnE5spl5ZAYyHi0JV6nczI/eZIkubz0lJBan24CMsU6dXw+
5PRgC32xpn8+tXLEusUaFGgmyihHY9c53ukGwyQrJtibAyVaHx28SjlrdHgsNzmeckrhJDXc1nlt
3JjdZi4ftab14jHfG1m8YcLbWLlrXX5N/QcCnOlSyA7W9XXz8D0HiQ1K9X27sjJOmTbgY3B1ygbm
cgf4B7JE7fLawNL4z9lo0UI/UffXrORNLc38kJNGyxpZ/gJ0/aFI8WyeLHnU526fTWCN2ZqaTSl7
VCx3PxMTmt01nuCedssuGBt9jX5oWt9S31rdhoK64mPx0LW3lZFzg130Yjut6z1FdEZ4vHnbR9vv
41O4chXuiiBsT41TSYD31pBNh8Po0Z2Ci8CkbQLSAVaU6GXeDk3wstY6qxghv4atw/s6EErQnxxI
7uDRf4Fwdccfz3KHvMflUkMES7bqekiAxqoD8ojfah90rwf6s1nTAheqaB9LiM9VwooDO1gb1ei0
kdxgfGdlUwuJsXxr7WPT1LtKfhL6H04qZzWW35v9vr/8iIrEFXhoOdnxzTNGgWlSEzUlkohi07Vb
1igtZplVtnmpfmENk+vNXpo2wIxLxc13ABD4e4PWsVMA4TV8baBtcg1qaNGjHh/K+fbe/cL33N9T
xssZSmYFuckJUqWaVFmlottmzA2Aw2AQnVjrALnV55i1Gfr2WKS99JWRaY9s3TQORiYrDXtgxFwa
Sx3MSMLgMDHEi2LxHRevfKLy6/50oXRv4yVCbZ5KBHVeWWocmLEjsDmw4ZDe/SQ1LE3qUnoa8zJz
zmzKWwjKEsoQ0F4KH/NcSPOVuRSqfheVUvkysjVMFiWgqEeB8KOVf/rcJrUErFlX+vu9/nlmZvSj
R58Oja4kSBfmncwQ7wDmwtVKpzI9vfBiQAd4LW135uK+3IJh7sa212iLLMnG11IQrz3MBWIDtULv
bTl53psjHc3E9TH0SNdYmOjr+nm64TpXk8hVHFAXJgJBIdGIfu4nf/dhFDFlGSgwpYm3Ob7IkEHP
wWAGvzrNbq6inR7kDqSpdARIKaYB0unCLk2YW1qYg49zdUYJuTcYWCvJuukBTO9eWds7KTH5pv1e
5gvw9cAmE/71Rz3VdWM/I1Mz/xnJ1oeUWVREazTtUoI9iccjk+8Hp6UTHS9kEcj3KQsd97MfoOp0
myttdmzH5/w5eAXPOt9RvjxrKOIa1LELNvSixcHwMLiWbdX55gfHxEsqnpGxuOqFW3InxVrckxht
BGnrGu5ulEkwsuEQlfLU1G0Xk2svcAxiYdyfIvZKaeuRYtKsWxZBqSH6+52uyhUGm3GvFf+I94HK
zJD5JpN98JzME+3J6r63+J4/OCg4xRyfH8OXL3/nfRBEYdiMm6jnOziCTXnNoI1OQb8XMHXEG2CN
omlTsCv17av5rS9ZPKybBcI6JgQzbT3A+LaQuQd8huvv4YUTXYmNFZqUU/OPijl3wGl35Jd3wgxA
v6RED0DOJWb93rFe8O+CveXF49TH6wlqDTvXtcKnBDKeq3XVZVM8rCAF9ZLUxX3PXs2ABDT/rz7r
tl1DmcbT3GdZHibBLMhhQWzYG+dOM+keaDZsTvZOE3V6qk4X/AGizB/E4kHVpv+oeJN/Wi82fQxp
SQx28++OWy3HqPBRSvEpedfw0MbBkcNJ67jmpdIsiIPWjURuSRzr1pT1SiZL3wxB0pCW2iFdyQXy
q10Ci4wmhSNpyAplbcTa4EKpGYfAb2p8fMuMB6j1x/CxHxPBjeTCwLKngpo8bspUzcNSuVWqchd1
uW7qVcZInqDQVo91m++k3dm58jGVyPvY3a31BeDpAAiHbq/GSGXPZ6AURewdvNIzkulgGo6bvWzJ
VjmdGaNZtId2u04awUDM55zq3vsGUwZ35W63ksYrg871/nuar0GbcOm5GvPHQe9TSKiaLfG85LFa
gzj625KlQBoeeG6P+62dPJPGhLQD6JdNPLqxH6+5XKw0MXNS9IUymXWhsiZ1S//PtbZLktXr73Pq
mpcZKfovhiG1vS6bbBi9RleRnakqtiOL9PUU+nk276ADTIlJf4DAEX2jIKOikgiaiR+GheixSO7d
K0APrm27InqI+ANE4aH39bFoHFvTqz92jMMY1VhXcIvm1uF6nEypst5CZuX4AE0Y3jt6G6GJHpc8
t5yFpNgMPrORjRvWb6CsCo9eYlK7VLl8OnLP8GDWD5kI6wgKBXP7ZTdGqypNRfpMkeisdBl29Osy
D9uXRdR4Lv6FatmOGBP9xLncI6z2+o67ABhVEkvouTieELBoMYgs+GNiMDJOcznStcnTjcEJDt/T
Uvhmms0+0xVIKlcwMhrIFXX1lMuNze//s60YeawajJl692E7hduwKFNWH/DIbZmgPSaOvhj+GRuf
RlFcI3ax0GPMlQO+I5tAkn5wHcxG68EPPPwFqXBxXh2hLcXwT7VYGjTFBDf3I0raYKVcXqMGJxJz
rLG45/WR4p92tzJA0QQVzLl3MhSPusGacVikjT+6pymROhkwrtQJWJWufnflVy5Jj9aMkV3cckOa
1VygmkRDRE8kQBaXCIhpmYOH4hy44wm+DXvwALyk78fENu7+ZvAEy+xnJh5luXHdjvVLnjkUTPkF
0BzVqOHX+KQhp96MC/3nW/b8teWTMvGfSc9sKh5M0dI3Gv5Dkk3PzdFC6HaSehPRrzd7NkfbHd1B
GkP1ZHFElqvyvV3yOfXi32NiMMYz3r1f5f8rPyJPY5AdWVzj1+WO3Mmn8xy06NDv+PKI9kieVuFo
/XTLxP2LtTYpP/ME/wpc0C1NvkRdJOoHj68ih2Kx+z6h9saee3Evxwq+uoMtd0fFZuaxtCPLvZVP
EIRBvCpo5u5uk1zM9GRAUQ+PK0DEfXPme3Z9xyYNs2p5+4swDW8BD5ED2CaXQHj881AteNdwCCBA
E2iltuBRhdjkUlm08qbgiAP+2e2CkIdP0/sfOje7FTlzk1gMw+9DEFd2oluqMUG7nXYr7qnc8IBE
pS8dX0A3WBr4GJ1VyIJjFa4NEpXC5zHDTHbpnkZs/gXJJ8dsUg2IdbVPaY2oLzLs7GNLWL8hHJLY
0jiTJHM0nlgSYeZTyQjrvENOnhOl6xg/qs0kpmoAylUW79c1i+A7WTxKjWvmCfOHRARWPu+50cV0
qXg6qXvUFlij5+LvteEFrDkGMlK4vRylAsEWtZFy+aRPht1D0u83+eHRSDN7QP3MyB9Ck0yvhkLF
/6DLn7ky7EWtmIJvYO7Iek+1xPsAE0vQKT8UYr8ZAQOobIoBDBIIlS1bO/C2o5TXNCo5/u/T6xNj
Dr/cgmngDfFZXzfyD95IY51j/DFMHIuSrsyNCjdLno7rwzBebBX38AbLo8sWorQ/4JUyLcgzT+/J
LO7Is4OaqjsdrgVKovo2Jo9bwnT5/OWxLCMoH9vtAfhFH7jJV/urGJutFPc/Z9L/h77WFu0h4FHd
F5nmj7pxtKikr14HEIT6fbLzYugMfW7SCl92nBw7rql1JXSXwHeV5+GEX+i22Dn7eTfS0BjCUbuH
IBGvA2AI+AVkvFULuXEPkdi3ZLGl9wml4MCLIDkhab67CCdm4MdiAVyyTWowpa7gWlihAy9B7W67
rd9GffDs0TXhUkz/owahu8BRnrhLQP0liASAPE2qPq7T5eJJX/otkDXRkyMyqg21dh4BcR1rYXdF
+I3ddLL9q5cRP2m795aguYGdI5e6mM1kWfVAWEBKuOHyUq+UhKzs0J3FcnkhdJ/MyhsuCNq8n0GV
C1VrgIM1IP0bI/Q19Y7cxFwMEToc1cFNQGcRhBSqPgt9nq4dqvyFdTdWkUIt213W9/mXnbKTBXz2
sTsQ6kNxtmytxILDYn9qWgdzN7owpr7MW4pJH5qOPsXNZV2PtlLaHuKhox4TpKtDvyaDeRVedHKS
MR+jxOjIQ8KgkdxQhK7fM0jlINvlnJeMrqsZjUSXjhyFioiHcnbYgndGOXAtrucybhogaacERdbL
mT8esk7flWEBTn7cpySWJQ1I8BcF9ylckgcPp4p2Ti5g5niZxgYX48JTTSxnNpUfklzIrLdocxdm
GxaCzjHf/S+/az7asaUBjgiiQcao/g+KK1uuU8ZeQjbm/u/Rvn9WCNZZedLvwHzZc2SVkFE/sOHk
MS1BnGvfLmAmQBqIFZqMcvL4UGrVdJwQkbqUd6L7IVlYZcy7cC1nTc02pTHgP2f5rXqFCoDgjxN2
qYcpAmo+KFTKE1ywWm4kYoD6MEnDwbuQkt0voGEu+ddY5jT2J6+VLpJBE7aW5eRTZgY3YL1ElrHu
02Q4tkJwsfUmsYEd0rfK7xsvEj/lLjZrEzvUycHy6FxeGwZbyu7cSlb+91aH1kiqPKMJRysvUt+h
6TTzhp6pAHNWFswq3P7LDCpb5KbiI0VMu3J8gB06tMU581jOsoBjiFvbKKk3adHUJ4A2AyZ0skvr
OJ6dmCYezklDPdVU/EKMNtRSByi4C5ijg2fxIx+EqeecIpziujU3J4EnKB6ur5+t0hos8B1T5Cv7
U0d7lt7lX3+Pn08LQExH56m2kn20ns0ItmjntZpXaJ4R4BR53+M0M5agHtIb935DgDaPs7Mf/VcK
W3lTVLqzMP5eOySf26iricQQ9ztnpAYH6nCAxPavJwHJ51+9gP2gsrFYXEPsdSdh0soUiTLXLt30
ePE5tSBiXmQ+gdXmCuSHg/PGBe7Z5iTCom+GnmfyCD6pcRAyiQihTiPAgyNkyfRbBS5mB7FRzBnH
tal4DGnRisRDAVZJ8Qz19yiFGT+JKCng8p2VS36ymR8iNFwxxDXiKioqJq3R5qJByVR+WrwWMtIf
6EDj/Vgs1ukq3psb9zRGsWmInFlN7ZEQ2Img6Qcnl/X0FI2ttxQPH9/7Wg6aU2xi4u9qna0a/RrZ
zWtFYdCkHARM4HUtK3TlXkQm0qY8GLuI0yT/8EqGX5OrZXED8bm7n5EZJc8PN6zewK7QwGAvHH2R
zN8ZVlgQ73LSLgr/LxPX7mjr7GmhEXR6Ff+bWeYwc0QNeMa3K/b63AN+zuvFy44TmKnC1BEsOg1H
hB+WPT6bt5v/pb73TIVQ4N+e+xwelprM4X4fWv0HmLLLdIqE+he48dkO8gOB3sunsw4AhIYa1HY2
9az7d712sjwscI7L7oiHNfQuFGFCV6vrE+6jeVXUtTy/85SmaW3aBNGRJHlTaHsgeaH4Eh2IYqb/
mHam2ysndPaWuyVgyY1DEx2GyGdbz0JkUWyLMYkxmW8+pjsSidEBl8iW0JWzlpCfVoOYwJsOF/A2
qq5pZT2nK/Itnwp+0nr2VoLMQKPT+Ac//4WHNy3riRw2WpWGXNRNxPQNsM1Ej/3Omovx+iL0hcYh
eonDtFZnARq32UE410PU/TjElsE8MFXLfvBJ6893xfF3lpbNFY7lUBuTSdCRebchrU5DeOHX4Fo2
GzXpo6xjDyMfufiAQg/rdoONaDTWIZlZlMtqf4S/zQ4FucvPijT9CVto0FJXGYsTR+G50W/NZQfh
+YlLqAYQ3yS8wuWcL291hJM2aQBjUuaQlNMiCIz8rjM8XX7ET6wIqi2lS4Y6rxgxFIYKvW10olSU
f5vJ+PnBRuKNT7n4A78Ewr2xvkjrBmUWpPNnEWOMUd2LUaj6LxjNK8BTM/rlWYFKqRlUz+VsvaLw
0mhL1Rx5VXU5dNLCGt75IlbiamwN4A+YkLV9TaSyXkiCZQjsXifgfeMONfs2yfGnLv7hvZ1QBsEI
c3yFfBOI/13g5+7Q72PjfBswXevDzPv1nxo674eBqoWup17kEzldwrTpqx7NHJhRO9BkFilui3IT
CPQ+GaO9ewOy+Bp8wEtvjGJXzzIU0o0BWqxm+sMvUmFBdhP9TvN7shnKoGwSTUvnYR3UI58XgfOG
yGz+oevte0h3reObtw4aKpsHfqpL7DmqOi02EN2qvpl/FhxU7GAqMj3u9z9XjFJ43VKuRa3NPuNz
mIP7ItoRETE3b8j1o0ZsyYw55MET4FWTsyPRssuf/MIl0UminURCDofGw86108zMUAaBlSHJV4lY
j2PYm6pc9+g31GTe2+3Wa5wVTTJ0ZJR26HXzauZx+KTCnUPAZc+ztW6nOFutpHOteNF4yfefarpk
n1nSLEPrOI5eYgGCr887MrZ0GNDfjV/febhaVkbfqF1coiUgWcU/rthhi+YU4sDT/Fr2Nzqhb7h6
gctDBbMvJo3OMVdvOpW870MS4b5uT43cCiw1HwkhcM2wHf+v9Qd3aQL4twDnEzmSpBUEbhHFbRdu
BMId1kPMDPsG/jJQV78H0dx4uap5sth5V9i4NJI4dOCTr6lw9ieAYgYgwRKqIjPzuXeCAU3Xx/kd
5TA2wL4bscU4ZyoGMw6EGUR8dz/Ytvno5h5asGlqWvGxHkPQehfVvOczdLshx/3iTiDqw64qpANQ
FwnCzUlgKPhyrD78FZKueyWW6GCD2iwgs6xQzlgneQ7WEXnx8cy0zjTZIYyk/kIE+cibLoEV66eF
7D/fWpu0LfSPW5mFCT7ubkt1a9+ZEPY0yEbWnOiOOhjjK/f2a6BuWVLpu+w9woBO/80tvl6vgw7r
f8Cm2GshYxV2kYF5fJmRvjNlmigBbYotjeTm5recjUG2MIzn1gQeD4Y6Rl4yQkTSNs70dKRetdLg
uXliSQuQfbx4QnJuZ9MTa7/5jAeTosyLoLDklRppcqbVNQ9Qd7Cht4ZKZSSI7r+5xB4ZI6bG/Osi
oGh17QGQ8e2+kcUYsIhNrWpke/j3Mgu3EFqIiHlUbBuTloQoxuv3i3Os+he3gl7utiRcrsAqflxa
m23n0OUvpUm5N4+5xTpQObVCEEp0NGENeRBdKltKhkqDkVFuO1jv17IQms9fhIaKt7eEmUqER/ih
D/KY6b/Fwz6o+UO/PO7jVPyPF+gFFEO6InC8jB7RhZsdZ1SM0E5RtGdvPWYUnvSutNmKCHbhNh/p
dif/K7TZCIsoPnb3TkPTA/mxI8WesrzGgZkOWZw2xcVxF76cVMma5QP21SFquYivWvmC3irP1HHp
kvr5ZFgz8Ooke3D/Xr7ZVDwJCV6iUMBe0VXLC3TsrVlaPIY7nsa3uoqcSjPUEf5JFNkrQ9qJYK6W
oFGLXDsyzvCGbVWyw6f9mjKocJ5B2nCHRMnU1mE6IOTQTGHAbXArTG6Uwdr3Q6WNsXRnCMIcbdWy
Y7oFJCy0c75AYA72wPgeVRHFyoUmxOeAK6Il9HfPawrSSbwsmPdzcPAm6PtzYbzASHHeVuCge0ar
1I2WL3NZSTzuKJbUdX3he/kPmOS5DDtH4FrJR6S20o+Ad4t3u0SI2MDwPra6a6QCYIFTkPewTTHe
yKKUhaVX8sgwAXGP5H3po7FUZv5i6Tl4czjUY/KAGDmpycnFdkWAZm7H/wFhTjqqyWkU6tbhcPyu
x4a6uV9su6qUQl6AkM6lK+lLXesiOJYWzBt4yW7RUAI7uX39pMJioruW3I0gnYQL8zyHQ/r2u4VB
Hx5y7Y42J+v78d0Wx7J/Quyy0Gl7ypdRJOopCw3ido2aYd0monVBswl+NM3cWKnZXb/EVq92LwWp
rVxzK4Q957yXV4vjnuWKuaFlEuILNzCW/ytX0wMSCJenntI3EoPg0oARTQqCuVqJf9O7LjvX3r0H
gfrK00y9tlcQ06t1e3PvqZwciXiD/MZYD2o41dH5y0K9sUGMDfyVbvb4BYiHRcyaKV2rsD397V2x
XpYIsgOOB4sPH3cx16k4oziqj1edAdbW18YnP+JFLNLC7AFkxrvfafQke7NTw5iHNEKGBnRryWzs
Jz5fejvZ5QJti6FQ/26TKjLRINPeFpan3vmwvBSJ8Bk36yvvHt5t7JgzaYI9LlhVx1Pvu09LuyWp
EhfvmLndUtToFjHgYlGnnZMsBudSAJFwx9ffNeYxbxBjAV1Z5Dt4fSqSltMI1AAGyYaQXJjT6YEe
1MMWFTZfHQrwintQQX6fOTAANqtrqZ+ULvgJykagnz0rJsFZbEw3rEvYwBICZGJErBM7nAnLZKVq
LVtH7XjboRMweSYowC/Z/0AFJn4jbxRVT9r9I9BeeJWB9IrcPNdq7NiltbsIjnp7F/sWS1txYjgc
Ps9QW/JsWmfYrKnyUcq6rBAK3ObdX0+HDspWOeXMCDHkd9+o9gjrsPDjZkzYcRzWRUsmu2Qfdrqp
57da09bM/iv8BLLE4NekcJ0c7u5Hrdm7/GzCx8EJ5CY7iu7ce/RxUQcsQ447pDclwLB8vv5a99bF
b5W+6+asbj0+R+l6UT7K3M3OVRrtQZkDUKTmqgq1qh6ORR1s2ssqAwuUt9jdU2F5WdKO9nV8TW05
likbariSz8CpLstnimoODpWaCNQUijWA3J3h0sk4BML/xs7Er8Wh4RQ5WuBo8JCIp5Aos1hAOtjP
K/7e85ZA0QPrN1jc4sh6mGl4wr4Ooux5zyQAUyNeGIEh1EJ8dvY8/iAYiQp8G4mBKRogSMjFADH2
R7ECuWAX7CduuwanR7NvL/ba7k0N5fKecVWWQuKpH1iKisAdUX9SUCVN0z7EKrx7OXutthUog+hq
FybNE46S4oeS+VbzP4fRPXV0eRudRwhJwYnUH6V1wEZ75LjC2rzPC1IYdkaxxa7O+2GCIyzNFW0a
jOIp84fnfSX3EBlCjHgjZADVVZUJLvRx4L3poh+ZoPz6M/LrAeL7gBLu2RoHU8/z4vId8p8uS6P9
6EDRUM330sAdbiKDhDVG7dlo/+SK0ZAxBuEjbdARU1IbmgccSVhoukbBfxP2INQRzoq6tyIhw0tG
97y7VrV/92Sbn+EemtXH/7ezi4BLiR0I3nmiqIYnRBNqNpHgS6yepnR8Wskyplw17JiTaIiAJgih
Qo+ZgT4MOYZ4iphuhnBoCvjJXg8vTfuBVgqI+CP6vevDrMvEo8tHS6v1s8MjtyR6VcPwXZDGFAuL
ZyA6YL1cGr/VRj8MsRdzbrL3JguodbYo8fAfJZfO5ZYoWYgnMUOukf4VXD4vWHSGpQfE/3gLW4rJ
fWUhWhmu29Kg+1fMPuhrDrOrPzogwHW7ViEDQRYDF2ab0LhQulJzJxWpMa3vpI8SXElPjYbWsOb7
veLYk05bMc0JmjTzejsyBwd/vYYiDOW0A3C4qa5uLqy0IMySjC2weIZCTmU6fa6o8xrLF+seWlpe
KKEkYMFowiMMF47fWvGrJpiR2tFkVnH4sdizkANDBDiRFWn9bH9QFo3YxOSz4FRKLftWQLykFgFe
N74vsa7UgrdxUBbH0vP3nH8CF0C6bWSraH8upqV89V5FYDXfyje8Gm8eOy4mDvwgYn0w7Wt4p9UX
iPT569iknDG54agreKEYqOCq9ahqfX5VtV17R2qL3KDKB/PxaxMvCBx8y7kW71JS5ActHDfUsVDG
FuGREjyDnP4+Rsfz4Lqwpns0N2+rnT0kcP9sLBfbCX1iTmnuXu7CJdaiS16VOKeFUbVq/GKsJlUg
B0CrnA0skbpS0wvNhwsO8xgvHW1VkyJbGWnHpLcezFxBWq2cuJt0dQdLUw//npxiDAXMChnpFY0C
JKYCYgLTKvJ+w5/7aQQp4W3ys3eFfkwEUj2SaaLdYoOwZyWMcOeypDf0aE+drKRfyG2K8GIcn4RP
j+6qn2j44L7cVKQCt7uXISDgFYcjElQYh6uCuKg6xKWUSAs8Xz5xkNdYfMqdyBSQcFFvSZmaJE4j
pi1RQmXnn5sT5vtnIQ65uX5DFhA8hq0I/PVOe/Gx8bw61j93X+T46ImtzBVjuVndg9w7iOOQl2wt
twlpoIorbVJ2guqKMwyBZ7TBU6x+RVu4txJxxHndK2aDsrvDMyMxh0645Ire0f+11H4caIGhgNRT
goz8vANRzaLGNsBjSe8SryFfhSbFM6/C2/+6rmYPs0/QMpuBRB4hZ8wToVCPK4BDFJmNEsgZkyeH
PXWFO/Qd8Z+MU027j0vkEo5M+olhkZm3kD+vgp3VkMKC4MpVVy0RxYNoK61F6mnEvzYgP8StrYZO
fgRS2X5sTReB1xD9Muw+d0uApJRm4yUjx9rGIypzjE9xS52QBbzoPiAUSIh9H1Al6sY1H8uhuNfT
WKag2NLWXeTaJNNtz4eVSTrltCtOXyFMpU5pmShCPt6B56ew3jAfX562UXIlUe9wpw4THzCDNJ65
v4aCQ1+hR4nEC8hjB0KiZj7VE7Xunh/m6WLOf54Dxo+BaeOV0rkZRaNVXLcgQEsFULQ+nEjV3c8o
ntC5irc593V7ZJDBDs/KGOFFfkU66OJV+01K4PgE0kMona11q/wdFXCh9wq88LrmwQzsIANToPXm
uY86a/L+GcRHydfbUcphKjnWgjrGFiV8zCi/nG132QtyiY0XMEFd/KTot36FSh+Vcnd6Lw86uxIS
/8q6mCjC3nThom0fpZc8wrIpTCMMhHGDujcW6z9OH4XXcZuxinhs9Ii6c+eZWsyi9MdocdJ0YHXm
3nSyCGy5785FMuzlG6vjxLzET6fVRa2EyH9tyMeUZnH62Q6Job1hf7ayZtD14aosMoJxwvrBkcDL
AFC3Zxzz2sgZu4T7mJ+KUvfWs5S0Cg/qy9LFcmyT0pA5ikfWYjHY/jJlbdUHcNyKr1A6o93lHkZl
yk13Eju4zw5RCSWZvRuwX8SZIirNw5Kzuaa1occUeIv4wsuL/YQYuWG50cgsfpw6pCs2AR/vFxjh
Gc+GNn+dne6PvFAieYbOMe9pLlSxvL7AuUTq/ISncM0nDZmcsPCidxEWEqHXUuAD8EalJhkMQV1E
lhHsx0IccpT21htdd4cfsMfPkUzyGtbI5QmRajuB/I0X1QxDvThTgIPdS7eMqBpX3/c8fVItdTQq
ttD/epLdq++lHFiVybZFwk4GEjfjbE4YP7hVLzZvvWm3ZZqjgAaiFEeFQAf0F91JiUKw/fnTWDdi
hyksIpBFub3HwOdNuokOc/GUC+EIAItAgrGGomzUeWjsFxrPXA9qlH0A8RdCSBXOOzITe7Ds9u0m
gEAOwq8Ds5xQV9LpPIKcDWHDLczoL/74WklDNTc3uieAE9bsSsDxSuJDxlYeuR1nMUXVTGpZFXUR
SHNToiH3cj9raNfm6lUKe091EzQGt5Oy1ZC1oTZboRk5MBNlfXPvy7Lv9f26iU61CvIV/Ok3J3gn
oSPdq8972tXuIlqGghaJUOXZsS7LKkg1BREasTUAy8tR/FWqdbxVAH44lUInvgpK49XInY45/khQ
jJzufLbsWFKISM9HCwwwPh1Qrn4coio7WbxZ7y6CGxYSaDsv5/t25iBLgfD23J5QtiPcgbPu3foP
jSFPsu+IZMKkdic1soHGUit2Upuq9KofdvPDVAzVFXsbDqsOMoi3IQpi2A50NnLko3EIjScm/Oyo
ewOa2gYnzpV8rnyup6xPABQaqSNkZ/I/pY9Gn/XWTswVWK7OvUxHDNwkIDdCPF3wIGtzR3WVNHF9
6X+quNekug5DOG7oWZ9xyOnKQ8d/5sjbgfKO1Retz0DMyvfxNrzvSwej6uJ0MKrLsAtD8hfo+/uN
C9RUVTn/S12e1XgvEktHcnG1MTc/l68OEUzf9gkuAdU9hLJRoI6M6a0HYLkqwBUVPtodGK/B1Zo6
G0FeDtLVl6cz2DEC7hxH+9SBJbpfh5NSf3xj8YiXWFxlfe8NNp8FW5m1wg9BJkRdqNsNUUrArh+F
6vQW5eDuZoE/EaJWLUCMMnOrjVDJMlll8RWl/jg9Un+pCNvniHRaYClxJR3sHgKooZtiB9cymn7o
LsSyMD58YuYXrND7fXE9EnG8hs/QdIXz6iSXlK1jsvLmzY5FVWsW9VIInuFt3xJ6zsAHOjLiB9Y7
JluHVvNh1Z9BoL1xz1n50Wf9vzWuU0eTxhxO4bRajaZZEG74WbB59fhAau1y9KjJuvla3OBpAcSa
g5LvjAAbbZUCrpe5w0SY+YK05+4KjjrObC9E66AnRxcXGWpz1wsK6QPWTy7iO5dHT2Q2qHkBCFFh
EnUoOy+wmhDobW9qPktQZOswcGArihYtcst35vDdeCzWjirI0T4vxiXN8i2Fr+5wYUa6ZLFKEOzm
3LYl0BVSrOCs412/2lFi5vpurly5ur/FF00MtQ/W86n/VF5zYWtFE2xAC/fuE/u1qobq84vsdqmf
p2v8KwlcvClHQCb3Q6N1PxJBp9tSn8QhqZM+lj6UlzvI72SVWSchkfBHEXkK/OffjqoPdaCamWcW
Jo5Xc0L7EdyGE+qG4x8JnbDNDn4vPieH4vWPPUgI+ddrmr29/X3V40YpDFy6muBhQ/sBTzhJvdgW
y4q1jD1Ilxh3qfLC3XgTBMzGQViCm7ZHq+FGBtoHVTMml1nhQSOfnjylbuxWwwMD4YLiTtcq4dJG
8HKVgGuieVCPOSZohldGDv+4/rnvCVO2ht5JYG59WBM0f18DaWrRKqnylCFf9NCVf/vkD9/L4WN+
9ZWUU2I1ude33pbW3EzM7M/bQMDjtdmUdeTjyH0g7HkgqBH6wXpZ2AqV3EpS2aDH7kVKNZw/snF+
By8TuuRWrsLliYTmei0EOC0DYCyfeo2qDcKkKCL3R9/YnAHI+Mau/3Th2THicw8s2MvvAv6N3dnb
AxOfOyZek20nyz1MqeLAvYxTd22AXIG4N3BzlfxKGPSaEnsrpEmhoRycsuIgOOdJuYHOgpziotvl
nCupAXDbZc8wn71VdJLoMTNavXquDQ5o3MJVoFVdg4e0GQJGUm+5vuXZXlctybqEqM6B02vzgoX5
5UjLIPizcPBqs8EKBjF79xoNCXsjwWFDEkt7OgCQ7/A7hEtH6txDZEFYDWbJhfxUK7iT0oul2jcl
o6+VUzrjk7UD5UQQAmXEN+cyfd2EPmz7slYDLqmJBkrD0oWjppDY6Px1NRl7OYgrryFbB6JXaVuj
K3I9Dg7IJVIxG126htkIgpPoxi6zU//Si+vjO4xUv/cOwGhSa2cza8bj5wtML64o8cOP2sop7kdg
FQ43IUpXuS9ElHcTeFGWN2qaNoSBotFWOJF6uLjCEpMeON0VkV6IZQthqXJGhgnDjBXdBsFgle3t
2gIQwoYNZX1DUhXgoNid/JjamK4cfqlXAjJoU0kfMxa0/3tNX9tQtQIud4pbC6LknZoCyfMZVoNb
hcQJ6zHdXZ6S21ZdnCvu+VqW2g+F8f1VS5edDYh4RaEu04nnkFNzY3zxsSqfvs3g567BHXSHQaIA
Pc+hxjqt1gDYaliJGTr2yvsUQiEndcjaAPUhgdx0SSDc3ilNNDOMcb2Zc5oiSChfRZT5a1l15nSO
PDJgXhkpRiLfFAkYiEI34Su+mcYjEbnX0RY7uTsH3zOEA6Cm+1GvCAihILB3SShpHJpgKNQDVat/
Ko3i/jKOFW/IFEGxJS1wjzH3E011AeyllxXvTe0CTLJt+rFPt+8h1w3XzV6ksfHShUv28L8U4qjg
sc3Rp3PCyGcIRWVWhIE6QfDwrZ7rczGJpgQ9r7KQdoi40QODAQ7eyIxegHAWA8V3ri9dHqhQHb3T
35vx9sxmgO6tcMCIutyzhqLtctGaRDO4TuvGcMZPofcZ3fbjg3YFw+iLRJzE3/Ae/5PLHxWkLjse
VN6fRvQQR9pMYi958jYgxQxVYjBhQCXVkJNBQ4GY92gc0ROSpkq+Y/iUEQ42C5q8/18eu5UYyCkh
os7xTybDlMC/DqRZgk9up/N8vK1jlo+m2dYdO/JvV4eWuZ8WgGf1IYr43sCN7qEnTFDS95hcsF9P
F6UsrRsf9ANJa7u1YKxZwEx1VEHHRsDoRq2BKrlbnEcMhJ3dLhE4Ka3lARrH6KRHuw1DDzMuYFnT
+ipIRLs84myWCTez5obffBgaPtFczFehL70NYO01PlOvkV95sYZmA3jkgV1zAzCF/PpncBVpY+Hh
Oi7/A8JQFXm3FutkgjPE3hoGVZ5t2uwthVsPBDAnCgcQbDh9RjV6c9TyK/Tz8xuK74hrD6P34J4I
B1CZk+cKgzDuIDYUuIKiG8iRYH7EIpgY/HDw60bD7Vk0umPQeNGQvpItChcFqj4ZbOCIwUAQYNGx
KVScEmndQLDTaHz8sCbgk6Emyw8ucNjzAGU9Dqq5opROTfPp4tT1wM3Ytc6vIJA48+CFhPoO8IOz
/MbmcsNgcPRYwjg6kSKheIVN1clTu5h4pBATmDL3uftB31+W5SkPHdFbndREg93kSKIqukNrgmDI
h8/4Z4GVCC4YM8FBTFFc4weyX4M8Q8yiQSbu6nuNt7hBelk37Sqx2ooyoErfBh7QcUTmgKU+F8SY
TCU0NU7YTFoh6n6oIN5eSj6hZjCzC4sAlQ/P5x5e8ogH+XTnBbEEXS7gdaRMoeMdDtmb+Wb7Jopw
hlTJqWX05UpRDg8Nhc7bMLlKD9bljVs1ddu4fHkn+oLFKpbos8n442jkQ0lW+6OIHGC6jXkXn7mW
ZBmwNYsWrJ0zpAP13nqX6bD65PHf4/5QuWOOixMRhEp8n95e1mB56eeNQDEkRzpMvN83uKSiOtXP
25geBwckeIl+2Vbm4Z/cBfWIP5OR3mLFLK2dBYxuy1tv7gP/L6UjslcJ9mlDRO2gcvNVcyNicpo2
rTHyqUb3JheRWpCvGIPNMziaSkrEThQ2ileHPNfzFmleebNTvJztSNBIbet0Vj9b7gWLLXtzeFXj
OtAJ5aq1XnOHKBgxWOZc980sU4xTLUYuUUPNhNHr307efIAQksKAOOBR4s/aDVtHKytZtKXuZX/l
77GhhOzC0T4jQR4SLm6noph4TK+HObu3tZcEOmFNXKdN/LqK5aTQugnpefkVCf+QzdY5/kVxSjXa
eokQH5gQXbFYBuPAN5qgLFA0ANiBfJLPzhCp6OqMDQONFZk0kjBQIvhF+3rUJglsD+C3zGAeDjOg
ny+yowdGrIp/DyRhY/hktI6fEotpBzSIsUg+SmZOHA3stQqU8bQvBRuAB+rUE8MLxGdL+txKcuJ8
1MgnacUWdikm3ZO/xm0OwD5AYQLyP8PKf2xa4niXw2jq+86U/k/NCy92Q9hlibGw65drTUIBYkFw
21QY8dhm4WwhwNsZGvMQxgT8K5ywspC/zLHSSNfz+tBbe0ywBKrvI15K97h98fxAzEsUQIQxWFLn
Hsj12PCdnpyi8DqVfFJg5i1m2Z4ItuKWZmL+hTX9D8JI7Vk/GrXa8MRWAKj0cEodoFOKB9DkeT60
0D83ZFkGRiXfsjZDLO5pGJUhs4F4M61iGyTSEw2QWmljl6rXQ8guGz0UVOxf/nCIC6suxwPLfFG5
PPRYDx+kO3/nDJyiE79+8gL9l7vjkv6D86gKz+STlVTI1Srx1EofTzBlIKbkAlzceD7cv6UsarcZ
wXFIavrAlorBM9fgAkJdi8nai/JPvkqnpqSHn7Q9UyJgGbhlaaOvnCX+PgqQxmy/aKM0AqK5LRmo
bKGyZn+uHKJdZKmjzfYJhEmut5qu7xGcy8gNaKq+8xy1z+rN6OFJPsmnHgndzpyOkpa6Lm4y/fe9
9zLUPAvYVpR5OOw1RqgQYH6N0YQfoJ5WfmVC1sslzH042PJI5pXE7FUastt1Aq7KEDG/jwq5dw4O
OOJTJyt99kmRWDxkdebKS4sI/qRyAieci9wGSus9CUJwoqeha4kwlM04oQDgZ0Y//rSppf308hcU
64k36XzAz1mJGGsC8sVksNTq/eN6c5P18nTy7Hxr5mLZ/88BWrsv95hDH9HReWgwzIqalNuJA09H
66wiGhuS0Pq32eISMDkLrjkHbN/U7ySwYa8diW0RmIYjLK/p18CreCHsZLmgRgFJDvNzbM8FytxN
vJjdhVgQf8h2hxPHkXkEhl8VuWW+OkZNhkWgu5iHcvJsqY/XBwoKj/x1GHHvEIqy4hvRIU/L8v7r
K8RTJ/lXGh9447ykwc69wgRuLU+jfJdW1WS0TDnGHL81mfOgaMF2TLik5s4vPGi+7aLv0BtTn3QO
1EhSUcEtV6TU0n16iWxrnDJslB0bL4bYCwIVKbLTXEc3wEbthqsiipufvFgvsSKnj2ayRGMezukN
4ex2lu7GI3cQz02nuQTYkgTJDJuUutggMU96VAFQ+fUqpX0Q2uThaisSu15IClxmWOM+w5WUaXaE
lXpOt5bhx9eM2+p461TiixyZ6WMmSH5/ggQX6I0NP2rK4oRWkaYgCh+aJlkaRnZshUehzFJZkTY7
dDV4S8qCztj01SJK2RxV2mxM03BWdqVP4xcD/WIXfUNDhLfhO+teO/qRWKdzMyvQXPnc3ZJT7eDr
0cmSY0cdCueoouHtfXaY6xhw3IVpwrhJKaenS8kbEuxKFktMX+PFDqBSu002J4sSjb76+UlQpT2i
5n4ooypsM2ddr4gA4td8uH13U4LSrLkk1sATtEcUuU9MDjRoLIzDHAmbOq87gkTBCwaTkApN4QNy
ktcUIQYZrDHUK5dTFp8XFQpS1lbl7x8MjHXNBAW3R6Q5AMgFlCONkik7Hcg4JUW/sWq14QNvyQUN
BRjPh8x00qZQvR7Ry8HrIxxAsmJj7yM+mC/MReum0EhNkkqrXCeXGjzxwVqiqnXCzOoc+kpQvOw8
JV40UZIXYkRr29atXs1rLrCTeSxxWYg7fEqXsvT+X5ckUzF1FqUlvHOL3I0jVYbMvQtaT1D3yOq1
MYHTtSmg4okp1cjt8UVJc1X/MJ2+kCDfW8JSz3Rde/8RxDMm3YbET6tXQoY9j2+RU8QBPxIH3Zcu
P0pRz0XdHIy+cDD6Z12vjZxDeIc2+8KhTzLjYp5dt4s+sZev/bhW610AUhf58BiTtcmixTIZDHWk
ODvdmR071/rTeNDD5XEA80hMBvRAqaW1kX4ZUGXh+jNQ0CWOch1DzfhMbbGi/STXz1UTz/jCPyIh
/zDZbr+RoNdbTAkzIGkEAryfzPWXpabUrLAJxv9n7tYr9L8wGV7f3WjpsW7rAZ3428Jx2zf+08jj
Nfm4umMK7/OK6RDN1YezK509IAg9OKCRvQWnGX4tI08r1qrONAV7A9eQmrFcTPx8QwOongnm8/IU
kD+TmZKPlaDw10X99pD2DQXLWYpHb7awQBaP+hGj7m674uKic2gegm1KWhTIGuc5Zs4Akq85reTL
uRgd5DdrVQ0FOj4192p5UAY0p37/tJKGshkuf85TNsp6pSAN2nqqibyBubQYCoIOpfC8JWlq8ZfN
KgeuCy78740bn6jdE+f/tGFakqeDYxScWXfSxoJP892V+GFKZDIfly1hjo46zDfh0B5LvbRjyJkS
fBVTJE2WOZ70BUTWYj7O0pjv/sKrCRsYNJPo2E0dr1dHnqmXUsPvyaWXzVmAmxjEK+LDDFXQelY6
P+6fNG8yID2CrH8b+ZSX+oI/9lNW7KipC0GT2D42tQj7A0IbHJNI83uiRc7gfG+tZCngVB8Rr2lb
BNwfj5gNJq7hfoQcA4Igj6FL5p2qJfrkmZzrU5AD8Fa4iU9CF1IzlpYQFkWZEzGZN61VmG7vNXmo
xcRPYtd8isN3EktdCHLwNnQ4siV9fb9trzgZqYxzDT1UQEV57Gk2O+bTKuLSUbOc+XlG2iO6qz9a
A1EjRJIHn4ybSnEaTSk3wnKzr0v7FE+wl5yxlsTkjX+5C0EDq8gd1/5xpnLAxMe0trISRSeEPaC9
QyQHnb8uW+GECuaK92eS+/BPVGpqlJ4f1YIW7uhxFQg5Nljc3jgJNHk6ibP3Ov6LA1tPPRWRxzoA
i0hHDN7sPGRxHo+SNCCmrp738aCz+XgUQPCBvT/oOULBCZKlxM7PXuHks1UV+YxtnK1aMdD1yPLM
TWL6QZDGi1vyXmC/dA9oiqJHcD7Z5RorrN0tiszyqJdMAv3WkEzMYznvxhHxF0kXBKR7caurECmI
AoXSSgl7XoTCy6ETXgcia+hoeE1DiSrE9cbY4DZs8ONrX2rtsJ3Nzg+UXoG3oBkRkejHRoUqBd44
aZb+jYioqRS2iXZxkQaUL9d3T4gkMegEAX2ZfKL1l0cUuB31Qp0yQblpf3MLwh0WzxhOrgqOtenl
gbmW9XMYhYVsFKU64fr+aNHtwHdjToErBFJrS7BetJZyxRhlmnZTb9RJqTWnRXNEQe2RAM+IL+vs
9NOHGrtWRcMA0C6ZEUGmhNWQ8opNgwfQpMdmvz3qr1Zh4ukItnN5LRB2YhFBhpaZOmpnk2yEgSER
ycQBhVPPNOXrsEFKcCm6GQZ6bq7zPE44RyD9sJAHTpHEEo5NdWaC8nLiZHLciGYBJH91VvBFCbNX
1MWWbcpIR6VFcM4r9DE5Z9rl+76lmdChGjs6U1MEg3tNfgIgxYCzw6mHrUis5HNW2Oss6KpqPwaK
FTB4+66Ng11uM9Qq+cYTQQm7ps9TbRwfgP0seSeImPVWns+Mz9CROoDgWcylOiLuDWWnzxm8MCkC
mx+q3gxI6HCd390ealBwXywqs5SlAGQOK7kFl3S98H5D9A1SnUzxtML5uAwxOqt1JThmEZ2Pnikt
8Zp1SKazqk3+SU/Bg/dodbyuChKI+d82YtQ9Ymsc6NPVjRp4PWFIpKDIohqu5Xh5Vxw3K4Sfn+tE
idjQVFJegTw5ELbrtEjZwWu3JIGrW1Lo0Uusyg9N/W21n4rXFlOmMvwaYKVL/MHjebiToyrbG96A
f1/tYXdgc3ckSc3lV7KilJKrf8EuxZVYkLzSt50+CQ+gO08qbdcUMHSvT5HFoa1stY2SCIDFU/OM
2f4/AUgSER+c5r9jSt7aITgdM/+EVwO4G4fU42FppHCT84ck4dpH46dEesAj02Rx8aOnDZWi2gA6
W+ZdoqOFuUGIMiYmnhyHcwG6zvFYXUHx44nsmw45vjM7+qnaoZUCNn3Tqe8ekWDjd8LivJxlsVZp
4Oj46nt0y9z/JwIMyYucmpC94A0krJ5WU3gd1Uszsotcyc0n0pEH+p6IWF25188rAAH9IRYexr/b
P92WxLuVp6fdrMwV5Wh/gG1G1vv9rYgbeVfJUTQCcNB0u1+b5OZAaakqAoQEY48j4jUz+GVyDfaa
zBig29SFsm2KSVLbq7vV5RZXUDeKxZ3/k+GmqiNuveNHnkEDJSpbfellgNwRi5xIAXrGDeLJBhCF
1rho1FYgQapbnp83qZPJPGXWAUYVH9O7a8G+BDDwyeir+lIUFj6eEnxWaIYUWhaKOvsAS+3lCFk7
yxZqgmgwRru6+DViUt0OyFiUWZrg2dH/FvxDXhqbTVONrrNaScdUsYz8EKJ5dCAz0Qdf8fUkDP/f
CEQOaI9QAd52OpT+9eJUajqHOABiLXcS76w8m/JVUIUVkdp0hpndODuSIVBEjc5R4+1SL4hoXw/J
VACvvfOc924svYFz5lYRVt+kRcUrZ6wZI09bIqXJHBu1QQEelhW3rVDyrqmHVt4emUPU1ZJCUvba
pPMutBnlY+YUR9UAAggoGruXDzT7s2aEqi2JE9IFD0YBnDm2ew4MsZSANvYu63Yo7a9z/v0Jh2YX
p0sDPw0lXWhjWOnGuyYtRQGDy5o0lCWVhNRgmkeTFu6lMaUabQRkH7mVjm+tpTJY1pVH3mD5f1Iv
XVT1KlTPP41SaTYP7Xh2d9Od3oO3E0HsYxlsRR6pp3f3O9C6ktwhP6sknCpBHdThHjefmbVoZ4Vv
UGqZBCbnPKN5LpY3m2NhItZdAEuEB/2QjU+ixX3wti90GDHxLtUDY4IoKLEtpfzFRYKISzpGw6Tk
kVs9FRnleQ+z7OrAhG8YqYphfG4i81YYYHD3IRDUMMd0XF86QRGP+SWovWxeyZmBsnZ7kWZ72aaU
IOb6gkTM5hFPbVX0jw/4g+noA1CYRfby+fn65GOMvTKHf+K2lKz9wXFG++DQ+vDtv1I4A83CB3Hy
E3EoRjHMXZmGW26kKNuhLYpTD4eET+uEOUy/TapZH/p9enMnrfdDUrEaSZD2685oTccZBcnfo8wO
oohyp34i3bTeHWQ1QStHfYjrmzJMFt4HBTf4eZ7+/4z7ry7/bSHp0QZIqa5f1yf0xGKZfofvy5rl
SSOx2CyHo9UkKcq9fvX49D9MZbKwqvYrtxOzDqQ5NaqvcnrVuMl6wojseVUBLsvkbomB7++33B1C
QzfM4/vvTmYpwQWRdKohQLk4K4qtd4pVnJwSny86X3Rs4HQOlekpoTJ5di71tQpMs2yWqgEgmRrV
FXGRidMoAmyYh+piRu1AoPI4ESkDowkqe7GwZb2dkJuTO5FLaW2ptkwRL4t0rIFFCHSHEDCqhs3W
I086aFSNh5sDhACyqTFM9kANxrKm9IL0XI5woGPqz5mzouIqtUY6clLqFb3DwkzBTIEqwSMIVY4H
5noU3xq+3sBo4/PFAmp87j2P8EzgcZ6O3zJ+ODcRBpxMuP61dE80gRzaCmR/D7xXur1QVrQsioPi
25Eas0iZG9NSp3Glfb2VatIpDw/bSKM5nvduQsba3s7BUXlTAktOCx4Lktm5PgIpU6cAFjqeqTs7
sYdpgTEDiYABc9Kcj5Xwf/Eum2TJx15KuAatYMSBQAXVn9S9nzWZXONvWKQ8GQmXOJSL78ZibAhV
myC/KpvM3Q2aqaMWHCgUqyG7DM7uuZbKziYdlauLduAPaEa7b9M5Ly9FCUBddE86WIjCoZCfOkAy
cX0uQPj90/gXf2/yoBY40276CezAPolslfoCniv9clQ0b3F2TQHx0QwwCKLo9aoE/zTldNbIZQ18
DIT4YawE5Bmq0hJOAwEizwhpNZB5PTm6w2OnbX9vXyWmHazbV+9S4RCq6aOXujZ4GPPdyRS5ZHne
tvf2Q9UDVXjswW3345krmiOvDeB09PDE9lljqoZ9gxgtY8UVyM6YKka4UPJDJC2ZUbEy2FTpdDIQ
Thh/xNZRAPnNJGKvuFmbIXNIy2zeSvr/nR3ixOSTWYO+YqeawPIF+n5KcbtFeR43Urma1r5vkfA6
rh4om4nma+1XKB0iXl++wfed5NbvyZZsVbTmWRGlb2b6bqfid8cvfZS3kIiZbOR915MV/FwfIj/9
hlrexNCarwtdI8LXRpH+ugKWmRjXBKxQvx9EcTe6zYogWsM6OnAopZ0ZPzclPVTPty4gbOmdse8F
b1sQOPE8WwGOVZ4wjZT36vZ1ob++FwTUyd6MolZelohp0CM2VfcnsInwX8A7mp1mJcGdO1SYXpbh
Wv/fnwI1QYg8W34qreAL959Cm0r4oCdtXIFMWl1Yv0mSNbJ+kxZ8I6MnwjGO/koDGs6b8AoNuavk
dYjOGRx2bQdbfhWuzDlwKSRDcf2IPDCz3/n1u7p6gAHAcjQ1WNoJZqW4xdpmBJNuJ0qBx7OtLm3Z
OtFYb5FAxj6MJs48xWueBc+WnH5hqH1XEOKTm+xHoy/+oij9HmksapfYLDcdE9bTaIctVIG4+FBV
Z3oPSXCjieUj18einjGk+B2UZcJN9SPTPtBT8w5W98x6dBnS4t8KpjDHV6V1tmv3eg0VVKhqMw7b
1OLymhdD79NPhEHLxLn2Hb75w8NrGrWiHIaPbenCR4F3QHBYdWZhSxh3TWGLMpBGaWQ3S+e9FtkT
8/wnRNnaRZdTAIzhA8BhDGuCqKUlpKBWZlt08iACFVzdB/QPEIzrGnOnW7S70T7KsXTeEkKsGJ/s
kaaf5kBE9iIKWyT8LHXZc6gQuQV/d5TCrBeIcQgPR36qg5053szp8S0ecyEaAJat1IK7uX7KrHi8
ZKGzIP0S6eW3iyl58ogq5OqoOsVwagD9UuoICtw5o1rNcIjrnballw7G1+UkC3akJoRxF4gCtTYO
++W5CGgKz0dzBLERx4xTddiIay4zdh39H4Mm8nTmpvWrFeQjYz5uojO02DYmlXE2+RL+Z9oM3XdH
7xorc/ZpeGK6fqF6scevyeuKOvypp/5MeEsXW2ybk2DGq8yOmVHugo81wVGehPAlnIkWXgTbI9Jx
hCKQ+4rGQxtwICJPS1XEBXunq2qgIVJaPfU4Omn01urTEF9h6X+lthf7ZbB+3F8e5UaOC5cuwCfZ
5TfpVOo2dLscf5RTC/lILZHs+b7ONSLas2+kH41AjD3Xcycyn/PwTHwNbonUN04vpJ0+XCpG1KmY
uUM33CJ+J4TrJdsr6wbtJKWsgFw8IL/4YaPMzRwJn33K2brsqDuCdkNkdPwfZj6A1Qy+Vz6eAh8K
fNpdLT7trd4HTxIWVyXgCDsiLMvflDpLdeu4WEWUnJ0Karxzso2x2I0C/mEdpS+mWcNSmq2dNTcO
aPEvsO57JQRpEq7AcETl0A0TlMKHE8vgQ9JlGvIZHO/eXl16MGaK/gtEDho+v9aLYOBVtxJgtt6P
C1mhSkgAj9NxULcbf+LM2v597zNjSiifCehH0ZZbuLjhoEOxZYaoduPzRwZXgJacX1kxUcvhBYNB
+hzP/SYESXCzSiqIQbyQkrVTg+j8HElRF0le7gB6KL5faoB54wCiiC6BQFz4FyQj4ezuuzGW/JlE
SrBvI8WmFsLbTlHtbmJrmxz3+/QzULGwiYWcSzsz1BOrdlji11064VBEVSo+hOjuEV0EGcgsulRT
O0pWxHQLE821tzxHKvyn35ZlDr92iUa+plo9CsE9a35GazalQAPcXKSGbkfHQyhBqtkqRQo3skFw
YtZjpQcyIELR7IUc3QLPiiKeSX0aXXqf8RqDnHNgBupuTTJ4NCDCQa2obgdOU0hWYqsg7o7nfC4v
hiRW2XKB/6/7qTrR5Tc6MeiVA1WGr2w+6F0PJ6wjqW4tIdu3oyZxUFaNQ66ysc0tuFbJz3g4CY6X
qldSQXqttmyUKXt71ZkII6v9tIZx9g96ba3VG9u/GvlmxPHYmQgXBKm+CfVUQz2vhbi1QHMF1WtA
p2UGj53YnBijB8HofWXIAj1iff3Nl1zeSKVyQI0WUbRqpJlbAHuL53t5CrTznJ/sPXAB5zAZWqR+
Rr+OLLA3w5MLdy/zOYl+yc8awNmwPgDePV65Yeu5jhxs11TZgR1WS1h1bDVlRgFodriVxXLPLf6Q
DOXXNUtamHk/FTPoT2YVPW6jK8seq2utfkrRjeGOuf5pcNuvc40VhIUb30HfcKA2Ka2Cwh7P9dyi
4tDncYWn8VOiX5cVbx7YN57yuHUgwRtx7XMxN+BtCrg5O8OQQCFXjlPOn3vsx4qgMJV03z7+fbsd
burbCiZtjVrRuSYc7fCAIh0pTW7Yc+NTZwvOaK+lJ3cFrMuPBsV0QB0o1m+P+GwXCC44I4x8m/68
zwKvzf0G0koaRfnU3yqTghbpEQrvne2tO3yGTFe7qFYw81PcZ/r6BBLyObl5Lgi4ceYuSuJ1dKmC
leNBlERuzsJhWEnr7fGGwCNPdkDzQQrLDpuF7m/XZqfIVAOrGQdnM3eh7i7QghBTQvJHd1XGRi9H
wfqrBGRaqDGffRgfct6Vd+wabAZssUVqlk8kvvWkj6t9yRinlBjfcqlC76Fcz99daPUApmowBCSv
n6Dq0YYNlrh/hNL2AmXlDiLmhIvyJ1dYWaK6VADLc1/MyBT3Xq2uMm2s3jWXOpo3ZeVuVoMAI152
dMcHJDGywSX6T9ebmT1Fw1uKZ2hIC0ig/VY5+mBr2pJtD9IM3xTiRB1hMhaIDC17zgFZw8nQqs9s
VJpu4JKO9HgXhD0rXg4s6m/+RaYJxkuNUtFmQ1BboH23896gi73QkuATHIgxSVbc+iwIwFvHYBXC
8JsDB+dYszWZlqlSeavU3xBaJPhrIn6Ecuwpw7gIfynfAJLVtG0Jp1nUVRRInQk9AV2TbmFENPQZ
Z72smyNeUhzPDNdJ5lJLbSTnAIh2gVCsQkXpQ0vVGOBYkzKo5LVEjxU7PHPmeBqiXSRER4k2V71B
YmhxrMZYo4v/L+nOFXF7pcXL9nqniWpuPDSwDqw+iGZerG2CFaD7A5Lxm9hrU11dtT3LL4rPUfrQ
fB26eCQ2tSAxVIoYcLy7kHuXb/lWYQhttylnwmz17smc9792rbGLhn+Ml9jXWVKPzwIPkZ+rgreb
Bztvsmj0Vzu2iwMGmwodFOVfdyi7OxAIbB+eZsonQZDNzwxFhfSTV9dx+pJcy/1TzwNBcJaWuI7U
7TWLMSWhGkZHlrn5B3Jsn0T2fBXP/jIEHV4l1JP+JwBpPr8+ukGnDluGsiRGY39IdjH6VOTNFgpg
heFNi4NQatHoGD+hYyrwC9+hNIRxVYQdskPKNVFv2AMgXVb06Wnw/nHtXkgF9gUIg6s2jb+fbk/S
kVzsp45Ki6/0L8qvzT37fPgSINz9c1NRmlwPev7bD+Lw9Hn2ups5dhxL/9Zw2SUVuBDFdxOAO7nA
DjTEkf+RuwK1KmJ5cNQGvV7aFI1yamfoC68tkpXCvqHfUIrxmSf/Eq2XT34+IN2nTm7hO9X0Qaep
syiWqp24P5bOnyVFiA312h5pTLfuh47DCdBiOwJeTE6iX25fDjj8gTQ2uQQ9PUudlNhgaHhjkulC
LQycUg89VDPMYcMe/a1MJhRMb4ApRNwk0ByyNvX366QNCrORCvcuge4hY9dOsH916dJ5qOZK743W
RR8bfFRu7FxNaPbFn2eEBaB1Sd1rQvvQxytimSNgv03/lg3lqclzPLbznbD6Gaa5nd+EUsIl0LIe
3U9nkcesN8TjaSIblGCAzpPiXMZB63Kov+6BpdYStJGxH4Qdkcu6B/+sVLTJC8XsYL9PdaVfvzN3
v0peIApyOId/UjIuhriuxXzZtMzpn7vnHe2WbuF0OX0Sp+7fBz2FYuCS2ORRW8ztyJCw0cgB9XHI
y31V/zHPWUZpbqjxb7vcWYCem4KB8lykBkqAP22J1Z8uMUS6fCq8MSS1BIPnfiHYXLs9NbXijGSh
9d6eSHXDjxtJW+fKMmeVhIAOcsDYEwV7wRkY64MqILhlS8BRbd9MTHeO2i+EzXQOHOH1GgagY5eG
/NjVnIOP5TIgkx171NNDMi+5NrJwG6VitnFgs9N+KUnxUvWIiuEdLdlc6B7l8/20U8TVDSoy3U8j
dl8zStTH6Bbuz8Kj278WYujn9YmiwD7RdWlkPH+R6kdQtylK+bNH7CQqOlzT6/8oEz3R7Unx88yD
UlFu3l/GpedUxGzFkHKwa6TTDSG8mQzGD1rw1EFXhtatyGhY/p7TC35PWnooN6jc9Ioop/u+6jhz
1JI1YCbrwiSA3j3qkvfsd3DJC6pFMF73MdmTXZMOnxVRo4jrt28gWbY6RkbIHpXruOAqv+nG5uEG
OR+xEYYKLTLCHYqjGEjC+XDF1DxUqSoGTbPvX8YhJ8x+PyakO47JnYsycb6EEkFUSRjJun4uZDO7
AqmZo79al1jBfzKtQuwZtszwdsnj8u1FUc/c73c3jqlIWxvya0CDVApMprBUwXTuMza4oVvFmNZH
vCKQbJE8FPc6iMuFGuSZkAaBdSuIoJ4DPjxLjB1/o6yiEe0npM5+/XQ8YuSanRt93mxjhwwJClB6
B3+agb2MmudSQ94fRo56yrH+Qbqd+szwHpalzq4OUnB6edlFNxawRKoa+mDi8F3Huo6YvajCmIKa
vveiWad7HqPQpTy9TOUr8F+d4/XDp6yv99Ud2LWkfyq+lXJC5FLCiPZx0sZDw3geNF6K3O1B0TnF
105PWOvT2L3BbcvTeTTHo/gB5t3cmkECDISWh4xdddh0u15bLZnLH+IG/s5g+HqrJoZihShli2X2
7euJ5dOVtRQPdb0/qTrC8wjru2QiTnB4uSi38vGy2tDrtM6rx1URBtn5FnNfj6nW/AYbz1Uzb/HC
DyvuJsnEbIG9mWY63E3GBDxMq1wQKKsT2+KIF4nYtzPfoEf5zwyRzj1MFTpjADqG7Debq/DirrqL
0y8GCt076ldFAlhxOWoYmAMFrFGvMUY6MNuZhgwHVGRVXHtvR7OTPkqctW7HRxmkxnj6nvcO5ZxV
4Afj5UacUIfs6noGEjwMJRAIDIIgkAxXkP3fPOrcePf6w1+p1dr753wfudzLtilTDLDE/RlEx9PE
lhnjgsiYliGWu4mhYvW241XJ2RoSQA4JAgICFqtZDgn3jliqhIYbVuWsrpNj3lw71fHh5CjZNUmw
9ePLLwxVT4dnPRRTo7PET5Cj35PUyD0xZD2CwCg6ttcusoq0Kyjhe7od1iHgD2fo3sOv/dEA5i8u
mmXeAKMj8YZsUBUxmQMNmixh5HOxfx+dfwqlmfsi2ZV8XYvoAx6CfSVCeRRhhk1NNe/EXHvEBnDC
dV6MG7fY8TfajzFIHzfYcpGZgzAyM93+neuJR31cl9l+RI0gIj8BA1+7uLhR/zzWR/FSUSS0whwC
5CXMHXeTyCS7XonXkMhhfSQuj4WzMQaRpDE7o+jg89NgfSxSuvBHZvN15Wus41KdWj6Sqtng8Abt
4ZxglrkMyuutz9zp2FoJU6wsrIOnPv6LVaCPfDv3g9TF7RF6+isqEDADKQQh3RINqyvLwGw+STs/
cAKXjmlmxdHkwjTuC9DFp2M7I+vGX7unJ+fuBDOzdN8XguGsXDRMCyikTEUSJUHbV2FunnNmj/o9
WVey6H+YnUgpmzZwq0LLLVQJWucXdrOoQQ9d9ytnKJ2qgaMjEhTL3CBu2QmvzqomUAs85nmD5uqC
P8NMo9orhrQBEaZh7LHJhBWtgcgZJ1hhUPAIBldu7ZuWBaxcSwcPECCc3KXuK8BEzg92ryqVLWzE
4qvLKUb7597slvIwC9YlQM3jWqA24KXObfRjjiRHnNigchMViVmE2Nb2hEH81Fb10klJIKEvyL9Q
nlMB/4rWVzaNUm6CppRXtsTMCxIewy77lJmowPDvPiGw0uqzcnGvGehf8s3v6ZTBqHc4SP5HfIXo
dhnTTwetO9iG6E07pIRTQl5IJVsCNIuM36+LHNPrkgHJyEVSIklAD4eFfdlLBM+gQgVg1dQeAQYB
ax6aEVGei+sIb28Y4gZYdujq7QBJ2rkpgDxzgId9KMPD2u6/p+OqlSFgWZAT3mnFXAaz6tTpC9Y7
AbmFnd83ZYfbEso5+tndZcjGs+ZH81CRXIVi+i6Hj5uQFYOfvMIjzHXPiJRdyFUGYb55hfvQiyBI
Pz0HnZNaX43S0c1Y8izS+kz+QFjZrziMjCKwnNHQoUPg24afYxW62yVyKSLl/G/NNsHS0I0u1u/+
zk/7THqDmh1UtobkROdcvQNrsh7ZD1BbWannxkYSSBfWke0YgYzNRPWbppmU8XmjPZ7awV3M5lv3
3sTfQNosxU7hL4OI2aXzojxKru0gSoRAVMNkteIXZ3b4/EQujBtelWz+L7wWrkhbx4/tvnEcS9r0
ANnB+91uDcUuKGryGxzezLDQNAUpGGFSnvgAitWrakLYICzFgOmBSF2LWCc7juxoez2nfqCbO60G
6KScNxflTm2DwGYbpzDSCQ0/kFfaAJqY1n+0xAmjr+LeqaEEums0lbSUMA6YcMBJqVpc0GuH3Xde
m/Gu3R26EQLadAcJfFatniTMEESTiHjkvLW06BCWClrpXVRNVCtEo9h8J8YrV+u7vs4BxjM47Tvh
Lf0qf1okZlWYbNuUL7UgPYeT1pfdE6nSdayxXCwJh7EPBNi4MZo1bW/+iCr6BywotRC5MH9NA7ge
5gPXMfq7H/ZFFMqxSOJ+Mg+Y8kQ974azivaBB1dyoYheMQt5k49I8IF559TGrha5BMts6QxnXx8M
6IbtOHjFe10l2st4EXrQRq/0vG37VPKMOqKwns5Rzm7ERPBaEqglFWgxfbryRodFzvPcOyAIx+g3
WrTcYmKHNTL071JmLx5fhzYIMHU1bXaGCQJdc28UU3r/IVVCtPl5YUEC4RVVhL2LhCtCTHTv31Ec
8Cp0WZYR2alixL5A3xct9CUXla47OWTXLUxiBonxEjxyVfkDY6Z0iVCax33HwiohwUjQT3/kcsWn
i78qUKaeW64klF7UPg6OgTQQl4BSZ9CTiMezwPrDRcRNSY+Ab6PPw7o6P1RaP+U9zrY5LXXN4tli
xPUJK/ONroCv05SIA+afZK1vJMQUSjcarojF3JrY17ef+AkypKGyDhfAUXbJojOrOCOgVMp/NEn0
bpDSpaPUBzXICGYmWKpa+kHsEKZGMsIw9Jn0kVcnWs8l71exJJNik9tndzFUXrNIDOPJknhartY6
esKWMQIsYx77XK9zbMAIjrwOLgLHxBn8sp2/31I7I7Q9nZ7IIayNLF+KiePJlFZC9CWent1TeMnx
vssnrB3GkuFVfsQC55gr/712aLAMpCt57Ixjy6d+/ncK3I8NpdHInTkZrpbVdg2TtyzfxYUH3K3W
haqCK3Rd4yzx+TrnfP1Z9ZISWu3wVRIQCSvzULd/0XHbei9arrwhFN4VzXszgTlnGk8CPGip/PqC
LnW6lWzQPPOL+Z/ZHmDa43wDqPahfHXE7WgRpx3jqIHdWgjEEMbOUlkTU4w/ixkl4/JkaKPx02n/
xmzWgUULffGFE8iUPD9G3Kd6/taNx3Koom/2Zm37DH71mVzu/3xvOPx7dpCOhtMmScnjtXK4ow72
YwVAkYFwpwsDkd0xp9mXfydPKVzwyyOMpyAF/dZWIv47565JpqTB/BHL2xcolu+cwHrcsiBtBomX
YEaAYwwN+Arh+aSiSABr6hwmvAG0rnOXZiNOaxobFo+q27zD1Bsphs0BVstgiQ40VACJ7aZpqXhQ
rjPs3Js4fh6jLjX/PsRtCRUztYhqOD7OQtFw8yxW/Lu5cYEgKKURxrGdWrSFBp7+gNBxQsLF+30S
QjI9+b7rMcISDWz6p43wW4HJ1erKkCE/CZ1+w7y3uxityEzpW56OqcpSS+PeGusaEKh6dMCs8+/m
H6JuOtIAYMTTGjIqZ9+u0VVeFzbzk215pn+39mERSH2FdHJLAYbyGjfY5LSnF9RpfmjVC1DxOy4G
hhPVqYVX6TbBnUskJX9qRpCRfgHALSmc5CE0Hd9jK3y/yJ26osHAN9OsNG/KAeq1HIwsOsgx5eXO
Rc/+U+DJXds9vjX1njuZKOt6BuTVCMadVvFipH/TByVUeCrkMhD+hhzQtz0ovlcAc8LGkT7RpmZM
eKre8v/4pI+Yl35UvTD5grhDIM666f0JVbP5/7uPAt0NGCHiUqRMc0O3XBRG1xQFQtBtGaThqKLm
cVRI8Ultfd3aW4nzwUhnLuV8tU1bBqCLaqsCMikV7Rn9SSOluW/zTGWWH8OKdpaMzurQ9CdMYlWk
WKdHYSB77C2lyKlMikwxCMGdsff6fzoJq4x2HVEW7uyjZrjyhbhjm/A/1NZL/70KFxd1N+tIEUFV
CTon7rEGtegldaQv1Kl7dXAJMdABt/FnYDgB/qOeHztqV0mq43mtsKGT1+6RWRLZ3Sa9JW/HPAre
MKtJvtd3yZtUzMdJEoiwkhVOSUdrn7H8s3x60a0q5M65vVBUKiHZpF5/m4FAoUuIt/RtmSYBjPF9
mo6EVc4+5fSkVUkfgI2b5RDcumUO9bOg2+a6yVl6QJKlhP0Pkf28MuSn3vkw2+x+okOSuyAbwLuS
UZtfCzG0Cb/77RpcWGHrap0TNc8t/npusmKWxSMfyisPLfdppAii244SYJ0iVJ4H3c7jYMM0Wu4I
I57Y7YufnkSjtwCRSki9KP2M+8LhvujbAmKaaVnmEpFTEd4B9BCEA+jeLhBclNWHSmOZOCNa80ag
CKMHHE2CYggzUGhhTrtL5PPR50vWUlZxvIBpbeJtyaYwN8lXPy2gIcQ5nNxXTB52oO680ar9YPol
PR7RxABUH0cFXsBJ8oXLTSgcAVVgDCwJAc/3o6rAgvslzFapWTF0To9ffyk2iZZx2hCWIh508bU+
pVWzaGzFjWNOl0S0jw3756J5N8dty+uhF3XIyUriTQHoQDrVTHT+Lwc8cAQiYXXTW6NcuP6YAG+s
kticC1+Kx3MlFC/IJXnKfXucRJ2GemnpaQDCJEEInE1ZJYTByZlzjzpshCCoCL5HLb0QRVg51wdr
m+QpyOvfeYBctpCr+CIq/NyhjHVEv13cmWoKewHvnbdrybg4K4Pv3W4Mcu1YBzRJ8mPp/VYZn7mm
4GQH1p1tdZo+8PliInqZtvh2qCM0tnklasHllAsileYOFD9+t+8KAjJni7NdJmSE5C3clYmM2ds2
AcLS2ctwIXeJ/gMPdj9/b02Dx+qg6zYbhq5LqNBvl//F+cB/noOliP041GHjInvNU6XT6nV9hFcT
PFFKoiC20ZO8/UV4ENC/gGcyQG1k1fsGa6g9hstBLoky9Gskwphp6WXxzeiVA6rx9BanMQZofy5Z
UJUPH4IIAFeRDKtgNQx4jinPQ4xOrsUKfG6Tj00f6WNCLdEdD+hHecxBBtjc9/xFJGlZvHnAdWK8
+vw0OmngK2vVvsbHaEMJNABvtzTR5iyvNGdbLL6XUEwX/VFydlnbZwS4IfmcTI4/w73FVQvFDVBM
bPz2V8RJ9k8At5HO6B7s3VgTmo5XPpacCVYVYOYj0KKQiOOJsqEi2ZfhCd+l05RFD1jcodtk4i4J
DADD4TfC8iFunf7xWGY69EXxUrr3Nw7pKSK3yshMy86O+3gClHf9vPpb3KL9lagrrF9h+xavOAJe
fZfxHn5BluIe1i9anmY3uMCDo9PYJv64J4lGusL/s58YoWjmY62bUDQ5lTGK/Vwh0OluRtByqzEF
EKWd0sCJLRZC60NYGMunViKQN8uDRP2AMPaEmojed/vPa1Vl8RaPC1ISOAekAQUOXtlCR07oDi1Q
VbRyiZLcvEBU6yoIXv7kKiaT1qkyLai9CIYqec9Tkc7xd1ZkOG7bemiTJME7eA9eM7VpbLgKrgAs
En3FuEZ492TMS+eN7rYGcWntC/dlvWG6irc6lp67EnpwyINDLMcLTWbRrOrQqvacAM9M81z1Qqrp
DZ54Z9AzUFg32YMUP8sg8132k3n1TPj7tmELS89OROO0XwS6alJ0Oqf5tML/zws7hZz510cCV1we
TbRpo4oFz2nvzCc4gx6KtKEO2t0X92D+N72Cmx7+7+i/Glc494CLhn93WEr2K9YpX/NErJZ2WtCV
Uxfm0kF44pcE6m9WnVhowzsgvKbnU+IKYkj1CqpaFRpmJcF4p1YSNIG6KfPkjjPKNzcWxgnKHNut
dB1YaxSpqsPvCbNl2erXXmdM4wU8kMsqZ5UQsn4dDeeCcakJiaR4PDsh/Kp4AErCAFG+z6rmmoDY
MYChMwnXJe9Bse0VLuYbfmevYwDL9JMpW28upQhSNTYe/ZRH1hgcgjeX6jZLsHLTUu4VWS6fAg7M
W1uWGEYgiwllLvcqCnmLGwqHcAqOZlmXV7QKNF0hPb5tVKguEXV6HfuXlrt1TFp+kq9zoz4dvIGF
MTZwIYxmEvJZmxLFN3iCX3kSMI9fs0cI9ITcNLm66IOVsxM2vuC4+1QByy4YEEAjOTrGV8+fctoS
bxw+ujzfkHpU+DK/pB3WbSVUVu14XBaEoNtXrsqxojsq8TjGpqk3L4p72kRYUc0nmP2rVptJyFXx
KBWVO7JmVDVD8iM8AEomqhQYBE5N9go7wv6Eiu4B15Ez3y4Vk6AmJuingvSj3ONZ7wpXxee1IcWf
Y0Vl4yZFIFO9znBDghe2iSaloWPaPtykeDmPcg1GLgnMPiSVAgyjjTyQrQefQX3Ol1fpgUCwXNKx
YjBSMc7iV4ljiuHjRYv2Fo0zznjvQVByPLgTj7+6xexCmQns6Z+D45jwgao0JIP59rPIAnO0Y6ok
c/T3U3s/auBClFvnrhmOAvV4Se3ULstMt1laNHkA2og0XO5yH0kfsDGJUQRM7VbY8S2OUluvQGRR
A4rsa/ghtJwSitVrdZpryicXGpUbfidUCAB4VILwAxdZwlIqzZeGIIO4+ByFVswHYANkeF2DNsNq
IctsT8S02oyGPyYQb28+k083TKD+IC6NA8Z7+WOPJu95/z9PMCx4I37xCysTC4UL/3x9dnmumDkQ
rV6rtrJ0rN3aOUFkNqwaj21RFB5VkNrlskE9SwduedMi+J5NscUjW6dvZ0qYayOIOSlH1lrGqizI
1p1c4Y+e+qj1zWwZI76c5OAaaJVgfnZkROnpIvjmojDml6gcgupCEXVU6oR0rl4L+NKlzLYOhX9I
G/X6w1/ZWjRXb4SqcwFd76teMDvRWBGk8UTY5zjbhf9FGiLsgXzNQQbnVrYMeciYgXUSgR/yfko1
YKlLPUyjOYSn08EMbUQYOhTIkb7rn/ugRrydwxCjNZfPWnzRxdFMv+iSvCIRoLAETzcN4sQeEJ02
BKA+t9PXjpy0RSKOzwfLBYHb0scWK09O8b0m4qwxF0DK24oAbLM1mL5RvPdVwiyaSLw7iyXwTlwQ
ruu0VhO1aTOTpeGpGrpRlYl6e46me85xBwkzy2w68XxKKyppWnoBdb03Cwjr0E26NnJM/7YWnoSj
BxgxR4gAl31qkehTt/0ZksQ1Vq/uURyY6yH8Wn2i9oVYNBYrpFP92iXxYCMruMNXPhpPPD3Bv1ZA
DxOBNzUE98gXt2WyUR2ns6gVIsFr5oXWay7LRa67IXrOeqm/d5c0GoRHQQ31qPeXv/tdIEmGpM2f
gYECSw1UT12aZNFw/W4cDy1GXBly6JUUclSNqfBxde9l4p0k0gDtvRrCELLxRfYEPyFnrbipj2YW
guVJgbbnCiKTFAu1LoEVpWRIO/ac8oW7DzR964gCY78cWoSlOo2Jm6xIHhxX7vtqIeDuy9JJqE/O
zArximauIsfx5pUZ+rs6xyt9DyI/399mkZ7p9QpPFfiWTQFV/RLNvpom8F3wDXoK6atXnsiZnCbK
OsBfBMHFNIpJxa2akqMMpNcf4JxxEBZt4YFCEw301CPItUpeF04rT84hayePEXCP74Ex0EBLGb/3
3nCIbE7qPFVxewZkHSbCRL3dhjYWoui2wU/QDI1N/xLPXQqEfRbAoseF5T/yJScCLgTb04aTI79F
qIH5ToiZYUt/qy72UVolmDeC4SZ9U8L4zSFC9UgnJl/0Gr0iaefWJoM0Bu4J3Z+GqaEG+UXdp4Di
Uy4TQNwyKNkvxk3VBotHeOxxJssBUZRKM5VwDhG1+EJz2P2BA6LrB76u3CTg4i7jSWKghGMfoiOM
R9oKHE7gN0+AY+vdSw+JL2eiGW/bl+Dl96Bg2Pm/tanmlOVtFLrs87E4C4OkfWYd32SLZPAAa1j8
0jK0R5Rdb2c/SfuwWg47qmB2sdLFaTOqLOVsdw6ftfnFG0IUDR2ZBd8VxVJPZ5k30N3rtXhBzswr
rbTpkvqir7oE44BoyuSNyfIwFIbUz9MjcME/0dIcVjLZtoNWVMlD/5LinZ6q/o4TIDLlmrmmQyJo
KM7G0phGT1plPdLRxAHUNGUBhdin5hZJmBm1PDl0yy5b3xzw2nBaE/a/9BDy0D/5zMbKskaYlfwA
ORsqkuT9VFRC1SJ2Ln7uwx0z2h1iu1b03ZNhu/QrOUAk0Up+sZQwhjIkdGrdd2P4848CDV9wVWDi
hIuNDQ5cdemcveDTZKmeoQ4Lfe52ZXJxLefEF6BaGWgDWm6cTI4h2/1gAJOqM/hj19k4AkHGVRLl
dRgfMYO6zEdUF8n+VW0LlfuIEiz2qWynXE3y4XOHIHLbARlQrEbAAu1NhJelztc/be0dWDY5GZMM
Y8LxbPk4LVzqAQmk1EIsXX0gekL13imdxf15dwU1ReSmQci46B8LlLwEzZ1xqHSP2nrsH/bbExjC
r0MV4dyirTmeU6wiYH5kUUwnjnoO6uN/Cdc8Nv+NSlNXN6U61YQYjD0FEJMKltEFg5IjondeLkqO
w03CtSJPIBioxnt9IDR8iKOgnZ9EXjNbLzY4Nsd4tut6aGUO6oc/lj2MIiGN+e6oQKnpO1LkdAGY
CYkh2sDYSbmgRZiLovoxJNldh06nBS6iXjzjK/qdbFA31ed/zoyKKmdbVjMRbIkrgEeN1l94W+68
w65fNY2j9SS5lGm1TVGiroHDmnAwVSfgHx1ocBYVarMbi8QefPx6jF6xMmzHd+3xRpvzRu0pYZ5Z
X71FHSoVabpLW5tp40Ny/HVOeDzJnrNGxHBjvF/4CqYaxXDchiR7ADDVbEOHzG7ybHVAHOrl61Xf
pRjmOAAPd/NOEF/iqARTDCw3EkAYJy+bQFFfY+CG0HzRbcEwjFkgBt+TBa8X3uBDb7ZKRgOg5UmH
ifjSHDw/mFi9ommgD+yRO1Ie0VH0T9YfPKAOi6aeomG+EVjxn4xk1ETmm+87xetrkE4FYSesWGU5
dqAW2BYZi8TjdwhQwVq+jTWNBZ+GbajxkUtLzFhd9YBrbdg+/aa+A1X7NHN2gFW34G1AaIp/ANVz
pr3QdAxEPUjBPDlfev+DyvpIs7hmDVfeSTnoERUQAg66Y5CBltAZJYxA6NlrwzJSb0ZFH6oSRMWc
FqKMicbup9U1QTpf0Oe3frOXW6qIZs/FucAHQRFWVNObiHFC9Fm6zO6x+2uBzxY21Y8ouu/GC5Qg
uCPTAfJeEjRwGHGOWxS+FeosKs+pjyGnKf1eyDySZimvUTXIrlx0GXNau4ZaiWL+QwIEXiMU3F3a
o+EHAtmSGaCLpLgJ4WnPUdfIja+W2uFwNTw3KNHzausrQ12LLbXVBKyESxM5DwNI+HC+8+JBVF+E
ReIKghpsxvVY1wNX045BMieLbD0xNFB5zmKJmaRepzUjW6dwhHXSJnny5IFWoZ8mSuZ4cjJeE4Hj
oYLJqSDuJam1legFSI0NPDkvaMQZ/5mV8MFr3y/NVDEz7hY5DidjQ57i0erTeT1/gyU7n+xPIde1
Bn+qwe6S1RUFRs8XFb0cC6EIiIzVE3H8YUc3we3PYPoIc7ZmDkq7UgnTWDv2l+IcwrdV2hiuQrbh
YierVJabM7qbEOIbhK+Tfjx1sfwc348V5agLc2ViRkvE95ct3KFN76nE9hhEvpbSrJqrGMGFL55D
PWILosP9rgTi0GcvywNG8fNs2oug2hWLome1hicG/vB+E7whbfcPlPIhxaDG9JGjxfO14opXjf0q
5naZTAL5InXenMlzzfrsxstiOSuVJXIAuIxV0W3GSlxoWcLDxnPlIbBjZGY3YnEvtgHNz776KZYW
WxmReK77SR0j0Un+Amg9DhVHl9txs4zTy6LzysVTa1vg0PBB1fDWIgWRWdd1qdE4wMzl8HQVRWXp
mLgEVWL0JkShAFlu4u1RoOzk6dFGzm0txQSh/TnywALUZxs6xgvziF5BruNRQRJDzS7LgLZmq8i4
Q3PUczJCPmyfuRn8oiR7ZKyrWYIDVQP2+svkgS5UFORvToPyDyT6xpbpUXrrfL5YAnWLpq8ZgVRa
g49aj7G9YqQRPDE+D5zp5ByUzxnMmEl/JoGZuYB7hZFtzoO+rM8xczrCBVahQipye4XXEif4TVcC
VGFiAXm3wI5kneqyMMiIrxYuwamFEl2CqHTpuE3iSMRrYzFtCC0md4XNg+CMhV3qA1D81/YDttDp
sL8MigPh3PYqqGFdjgdAz0mK5SIuWgYpDwBBl6RO5T6bR2NYo6zrDAk4lYM4fVd8nBvFoV18DB/p
WLQ0gk6Dp71YJp6vGFEJua/r3DY3eCyU1nvP/d+fFPUbOKePFoSuw8V2A+gByAKoYVzMD5Xb07+k
YNVc+CtC9/rSuW3qlefpnHdfTHLVcB+RnYmLSAQhAenB0bF1gFPqKRyK4D1MMgGIewRVSOkz4wHL
3JwZsd8NmW9sOYRY510X/VISmAB5AOlnmhr1e7uv585alCGMPdR4J83IOULpXWd5vhk231sASiLG
iR+YCxiJoE/Kdgcvwf/RQKFzKAa/bStQlyjyGEUWjGH1cjGKW/cKVJqR+33+vGnh0Icr/W02v7tl
zCxnY8At6Gb3/gHfH4j8c2WDvTtvCTn8PH/Zzek7viqg0kj+/s326gz/a03v3PWOBQMIhHVfxU/1
XAXVO64eIf8GjiVzk5RzkDJJWmVSUW22UMmvPb+lf8/BpfIJ2EkVVLvxXooS+q4p1YuNy5dlqIhz
jp5mIgD5Cz+XpN8XEWOVfXPZXA6Temi+2UIBWoh9/rJ3ugdu7CNt0Xp0y85ea9SHs7Gjg2dHqXOh
vVBB+qXGetqG9s2DmdASrxAJ3Ua4DM26sQqSm5VquvyVGYgqEQzwpwrASQ/BhtoM27wtENh+umfp
1CWZLw9eCl1+OYZtDs84LD1iEYrFHofycDrVOakebzzCInchl0pOMdeQwcjSkKGsCb80LbBWvtYz
05rPxVaupv6XvT5S6uHgWmqHwSTkf+2WI2SCkEdmgXTIt6tHO5NkpdJz7ync5jxOlUQ/GNd+4ju8
t8tDfGkaGwNAhcMOETjVpQd5j6q3eUIvsTb7TkubnCZ9mGM09LqZQcS2BT4ia2WunX9RAdMH4Etj
clRBj+yNCbqP+htLPTfKD5RuXHKzHKHCplMKqH0K4AVs03RYUtA1+edS9uOhUmqS0ztCKJenrGnQ
elmB7vgT7jFCu89oV4GmDU9KSt2KhgatjEpFmEgPavM4nvSAqseyFXmZ+fFkVO60PL2YlUfQ4qjh
FXSXGJeSl6tgtSLqXBe5LF/RydP3dA6RNhpzNgcYvU5QS99cEF4Hburvd03x1oncpNCHJX2iRmHp
Es2qzb9seuY0gf5R7RLI6p8kdjyfONfkuHlQgWG/XBs423pExjcfKeh2wZiXswUagQ4GgAWbKeRb
Lq31m5AiUxZIJ1JaPE93IPLoPQPK5XlsixQpt8U/tdtjkPK4uUHWQ6VSwSd5Pdne2/b7jTkO9OuE
8pqoB9SOfFGNFE23tRd8DcM4wJ2/LnbCx4RWbJFkzeDPYt9VRXCwkfw7YRAyacL/MKH9noBaR0ly
I09gJ2aQA8P0U4Xq4TeBwXWK4hQ4OL83k6fv1vwWOagDfsLrnW5y+A0gzbBz4QtnidaQHIuGw943
lhMlVyqUNAHAgfqPaYE2w/UHp7TaI+HhnwTHax6CyhFUEUvrPRr41Ezkpy47nlidmF/rP3qN23z4
t2t5A71ppvRXVtWC/JswIz+z6GZdWP0EbIaFKGLx+89qVQdjEaUTap/pVcbVt10ETTOJVwpP+f+D
1kv+XX+VQ1muGsbZ1osN2lVBaRyNWD74VsY8KQaEaHUvUzxCbOE94MsGmcV6u4PApoxL2tgY17F2
sQJBTfQrn3FsWWm1Bwih8HFQyPY7HhYCqELZiriNFCbggpKCVdUj9HTAUd5j434ZpbD5GNha/Bhf
n26drymiNvqV0H/LgNAkJv547U7HOqdL34jAq0ZZ5Bh5ssrlufpniVfQ7EZCDe9vxOCWCC7bpI3E
Tdyv2bYM2oEeGTQf//znwoYwIC0B9opiZU869YutGh7aLGb1zbb2A9jM8jbVeFfbjbzKYFL0A7dP
nsEFmr7wHq/NymG/ZPNp3NFKEYGvmKBRMLInTIXjj131EnACiXDDw0QHZP817Aiqu/+DQ/l/h9DB
5B47F35JkSxPPi6L7hlsc0yZbSenPQ+TqloLstHvKR93QfxH8PgBaBQfc7XhNFUM64oZsUusZk7D
zwUokmbbdoMjLU3zza4zjiTZlepUkxdQ6jrhh8xsD/LEIhlV3FH4hlBSHAjGFRt5QcA2szMXrEkd
4Y1pSWAV+TUKU2xggwjsTj7rvRkt7Bc5PGRMF7dHPIZl7im3SbnLPa/DbLQQi0jRnWwiDtYzewTX
y+lrp2Vxj+yG88pxr1K+8JDu0MB6uSXZJFMdobpQHHqcfptnNLdZkLExdLHKuPK8oL94Cp1WSY9t
cBtout+nNEWgt6dBLYk/jIvCbr8JZwtDZDv/pzebOkdjPpxobFn7VYa0dXTMfXeAfF9Eqt44LNXd
44hNYZvWCzG45nD1++R8LROrzonvlz/NyargoJfwkVb5NDzFsBNBQQLHYzs3qKdYPd5XMi/D1dxe
Vr4bc1xBYqqme25VIRV31nIZg+dsZHaUgz+903WiH9aMljRdUbD+DTKIJlNxreDGVP5Zs0ffdZqA
jARK8tDnyFuERthpkd5Ma0lvx59HCFSkTfYj3jBb/q3DGGLCd1dk2mAc0cFTflI0vrkGy4fYYXeZ
gh79CHAw7/2WGDcCBE00FJhhBTgDPctwKGEyumneTGh2zhKL2zGkZNBIfns3mDTIYrhsIAF7VDWz
YMmEwL4fIWU6a0Fq83yhOR1K0kJYr2HEHk7+223XQunHdjoYJleElGO53oraDWLqNBoBJCIKSnhA
9RuyGUrzQ37dStn7VORuS8uhMNVFEzsLHd523QBMu467TsqHghSPdTO/QNuXqka0fWQ6yJkQgORz
i/aDNJcumCPhcU11kFFijY3qxvDv09uI7AMGxdxNLt6Kun4xV7NOH7CaNICY8qbSSgZ0lprNd6pq
b/R+BHfmSIrqW91Y9wK8sgorwPM1K9L5ZYYqgBIlPdzv7XAj1s2v78sdtlpwXP8KuW+UdCv5zARJ
ihGEMW+mFBzIlGBhHs1pNEeoiFzDsURB1C36q/9d6MwdbwFgL0LLi1sdAP3k7wL2d2lNUaBd084m
6E1WoLzDI7clVvo/NgfoASdZmfKBHHqriBlfE6U9wxcH1YBGFzLGmaBHUHni7t6LAh6/O9WnkRqw
swCNT5ZRS23TEvbE8eWj36NxB8qvwMP6+5nUAaytj2YZ8qrLbAcIMC+x9oy1TX5OUTRhWbrJt9/3
0HbFVAOp0pvbErg88AN/DGtcL43h1p2i+xpAqbkccdJ45+7oqWZd+1DV49GxhG4wDF64cUJMK79B
dyFAOPbgUMlh4MXMVRULvW3P0+xgR66LEgdeHmxDiMyt4i2zGmmZ5pZU3DoefMO4QjU7dkJwqDv6
QVsjnAxqaS24iqogERTZuZjKq4Bk1haKXBYVSW5JK5cT5cwENsUJaAbPBjUr/JbJqfcLM8iDhEf7
lRX0oqqFsBdYaITdZTtEetkBRR1xUqucFjCF5lKuDjxCy2wD3eqaAjTgoKzo2oIhDbkmSkooK5ZN
aUYl803HzHEdl7WbJuF6xEaIrqhEDu5hIjnBBXxg4DYT/AaJ/ULj1ZvspSt4EP3RIm+f+iXKd0xS
SwbO4mgZCglfs1arWHDHnMVikLwSCTWY/wmDKtbCRY9VR4tXS837EVGrgtebNFi5pYaBR6nuBNTF
IFTg/8XoMMhsQJfUBNdalEbk+Jk8QapgfTOwHUPJ9LhHnVdzG/owW/ajh1a2MpB5RPfRMwi4r2P0
z+iO2i8PG7RewEewcpeKtBeeV9Zr7AwtiK//bPBZvu1k3gwFakoq4Eozz27e2sPhwizv7OO+38l0
+1dOssZWwbX/YqLJrPNPZqlXs6lMQ3dUaFEVgw8Z3QyxpcdC8C84q6oK0am1h56oNyNa5vZUiCCU
e7XA9J3VVDP3IJfiGu1PXnKFCRCEGyOFlEaD3EwSlH+WI6byH4dQoA6qsDV9ADg5YajKmhuJjP3I
3DqyBAcj8kGkxbGJlCZ4vBEE0OtNEcEpI31Yccvw+/GC7EK/dmVi9wP0EcyEpN8yHDP9a9nJx3rM
/9E+i/hTe+ctTxW0Ob0np2IZi83y8Llbq7+jrvWiy5xRRO8A53XvWbpObt/QI4npaYFuW16vMjE/
AyTFguUlHyGx33hOzgxyXKCdsX9kMFQLYxIUpc0Wf7R2y5T37WszvN6eqN+c/KY1MLZoPfAIfXo3
2VBSr8Mo5qRbnnBfZzitgL/zYKcIyluoVOdtyHzNAERpxLULd7SchINhig4PvhckPlSlavI/rjfM
mekxKhZiXeu45WMEbU/t8KenP0KsPh5EZEFnfaUa6yv8aJK8EO4tU8bhAqp1mS+yj/A7hRioc54c
A76ItceAwxDnMrRG8akgZhl2DxurBgKX3mIxupfPzRqdbTdnu3MsX8VgULzTdw3xr2ttubXpcsqn
bQQuRrVCtEGE6u3Zh4AzOoSThB61g7YlTw+bRGjVkFhBrg8qcQCZxjZBdcYNk2bBmcq7JmY6sCTe
qVTmmPzTU6jkN/0Dh9its+Qa1mGPnSZa3bGhZvkPTDpQ1Svm/vJOxlHavWc40DnPryf8Ok8irg7D
CLOgOF+bhKoHc/KZ1hHR/XwC/2rSEPOyInSmRK+ONrk1pdPpMekAB6dWQwBqWIeile8Zv9GII3BS
3VocDdVUy83pwtaliRXtK6/ayWEhXEDCJvk2Ydqzy+6mEorSEbzVgZrAbK2++tC5hwwvyTmqQ16k
hNvc2oHgUwgLbSJ3Hsjy6k7MzQfLVQ5G+A1ly55hUpEDmB+pVNCesuI+VXJWhX7lbnHpxmQd3V2j
zRHsF0FIeRUxVyHCMebr9DiWNzDv64ktPF5QR604jckz4m1RhIX6kOtWw80x9ORyaHlGtFkvOS8P
uiQwo3N/HqoKGLs9PUmOozuWhICdCiaPAHqJCvNEB7cq/UVfc11dKNaX0wAWxzo13mdfXyOqD+TT
IscERQDXFleMaSPGhpiVo9ZyMlc6FP2BuPXgmgj5lxlp4zB0EH/bVup6lrJwO9gEOBfjvupubRlv
3FbtzF5OfsgpcBmMzmKIiMxxP7nBlyn5OBHEXY3BmsyQJuYIvZfX+q1FjDZP9FIwqMXSzjF29UAd
BgpwiU46kEl/Ps1rc14YI0n3IVzObROm7Cw/4OE5OiwqtvFNPVJCO6d+rVb5CTmTrTq+zIXH2SQ1
Cu31lgRoHgiWbIl8S854mzOoxo3XrmkbNpDXjWw2+Bxm2PmWkDMo5DnILLhLl4bT/PSQjgsJ39SO
+/diZfLuiK5PY9xCtHWBPmSJ9zvzClbbTPKc5eaBEH1twPO+5nEtHdE5aaVZ2Obs9YjBmajTlpxI
dPosdM5RU0CpirdlxV1SMtxhiUEjMqV3mzt/SIvqFAHppKTURHMrz8vHjCvPqvbVREDk2Bj+xaYa
MA7TusBKJfcKLVEjYDIKYFAaKBg32VTXWR9peuzudgl0zCgJt/j7wyMg0vMReBsp6VWo7oMHvjiq
LtHQO2vu7awgNZ2URM8JjieCGgCnZRzP/gdIso3iufvYwn5QHx1DSdx0lS4nUhtMvDAtdXV/Wl7V
9Z9tCOJhMH7HF7UJq+1GhOnfeMUBpn9jWkZ3qhJRqooXBoT6F6pZ4wDIPuzMvIw6IvhI6TW0+/zv
W9XzTIDPgVn308XBGQZAw+qreyZxnNUiXM7G+fGiCnExBQQwbPNf7624Tnl90gKiDNlAvBl/NmgB
ahamBM9bQ5L5oRN4zY/qREZmv2SgdMOub/9m0OhUMCAUWm/z+yWTNeJRDQqZ+Aahu1O5n0O/Zr9/
ZatslLtUeGdY5RkaFuzAwiyvdFavyoDbE4ElW33/fZ+OfdjSMZmIgF22IuD8+PY8ZYQdzwE+G0Yx
akBOTpLR6XGr1CYZuMvr408sq/BECHSUZ2DZ004kUZ0lBDqFJdHBwOked4YZ/DL6iGCQqZfKlnLl
V66+I4fXdVRp62XsGcg+4yODiyH3BjgNhMFX4VoEOmq8lksSeTvdINYkUWEdt5Goqb2aWQ7dJXjp
nS03DXXz3uptqxW/PdQyu0NUV7g9z1UYUWp962YqwQNdYdRsCahWVi83LI7cM39To21IVP3aCG6M
CSkFzy7X8xC8rBiyffpdIH/HhTwOgNRwvc7tJNHenxjKf42UOI9g6wpJ/bj3AKkI4vBu28Jdo2fu
D3zXHE1vr9ug23nnGpkNJzinPnVbBvpAKbeCIcME7DL7dhNtGLPDlRb8tlZnTWSANSZCZTNsaMnt
LJ1YMUGUYhrAWE3ATlRA18Qj2WBAdid9Qxhj/FUciwqJF/iH6XwFmvgwEpkbSuWFRHF1VWYKmIXe
0MdM16x2XDyJOlK14SjmSOWm2hQPJ+lXf9XIPq9C7CHiB++NMZ4Pcz9prkqJUtkn84KHvb8cF37O
wRebojh6La/A+hImjz6rCaWRhNY4pJM0c9L+HP6k8XrCsANbh2LAf+j/X5FBBzBY6rDZQWrW9c9v
nWj78yzz94aBw7j87yq3JGQr0x4v5qWlHBBiJDBvDDsotixkh1UCrCi5MfkWWswNsmGYEuVw2UjG
6xInWhcrMwbf7LRbF+aUejhTA7By3QD2AOy+c0tX7WSqBc8RTLeurPN5XpJyxiT2QcCG84FFI+eP
zksnOoOOL1iOxt0kRSqxdkaKeFy8tsWo1V6CxPuxvILlFXLI8LDMQ1aHI5m09AbvOmXgU3Sr94Il
qP1+HtXtiUGkbsfBVS4YF3XWAASrjRSnQZaS8NCbCBAwtvdYelkGyg+kAOcBTmfexL0SAaiNaYWP
pk4njDD0j2CU/mBKtFt6j/bxDKhnTPWi5k8yzAbKe/MaPKj7pXD1yOZwIBTBXK+EA5Q2YX+x5dL7
fTn3Kg0oUl+Iz1g5NjAxWt5Ck5zN+4koINm4id/Gntebrm+Y2Z9VZMFNHFSifV3H+C8Dn3E3CicX
axd4/W4mKT60o7xTObNOTHvz+UX9m1DS10Pa8h+n9VkDqJgqK5dwRoqypQNcDOuDPLKEAvB1AvM7
cK7AYHD3Bb5cb1qOC0JrBEgRYJUOSLzkP/eg329CYksvcUKpdSG1y/vTN7gBg8yrs2YJp7fbWfVp
wTZjcBLzylp6f5zktO25584bbp6+XhGQSbJZVC244SYNuZR8mRSV7z7pPQZwriaUxOj0JZWG/dZT
NndsklRIOC49YmWuczRR6PbKXMh8vdl3Sjf8emvqtcpPE1b3Y+eg6V7CbdJ0Crnmc+ZR9PoEhbNZ
2OxHMGb3lYT0oShXUAZaUOKj9rVPKHjJEnxciyELM//JXOik12fhP0QDjTrDWi8mwillW4LZ0J0S
pyJtigpfpBIMpubCy/Er6lGBJN/wMhqs00d2COrhM2mLUxxPJxhkL+UZDPfKvSm3zfnjTC/6Oarg
yiPBaSA141rdq1Dq4vrNtXXbFft3yEACDE94LL7SCAQchqjyJomPmvaDb06Da0DXgAGAVIK5nyDQ
1HuF8tMYuAag5kk5ybZOkNYIs22rB19/LTBXo/Th1+2aXZK4WkLJN531FDvExZJ4obrFf3lvUHB+
gCh4UrESMfMP1jBMm4Agt0jznp14xEzEukUMLGruf+pXfTsrxtIB3Daz2sCkQAaJciAw8xp2LNZ8
sMK6BRTitV0jZ6ZmlYbN3sholBMSIgwSlRtjhklTq4oO0KRwwH0kRagKrRc2tTgzjN9y+nTZakot
+MBBX8BsGHhnTVlHiEh9bW6QUVwbEqIBdLGKMpldaQpfxPhjNyhW+mLymxBqwhq9C2QCo9mSEsTD
tW9ebwbxmD5ftWWzAQmK/rtDNWwKBrBkk2kQlBwBg9pkrOSL9MYgaHEhsm/AmQWFfHOT3/8IsYuY
kZBKSKG98ZaH7XHYjTze4BOlHkx1tsDm/ennu10j83/NWtQ8f3QhRbXL4VxCbN6Q/NGVFAbv3wbA
DQInchHOpatIAl+kmulnj3vw5gynCXV+oDCoPKmq9fO2sqJKwzhC8qeLUE5oHfzhz0LNfoMPaQeS
lMGSe67pDfvvn18S18fzOs+WEjxDpWo6FPOlPh1GCXiT64481M8oCsCh9Xo5kyB/stkqfmIuCTuY
VIT4Hq0HZLvO8UcZm2pibWyRj34G28KWlPMvGeyCJzHx3KGozT4s5luvRpODVTDRArrJZHNOfU3w
tnz3MJaPYq/wPBnGZpKzXkLnZ3DzYwggsL74aJHtUQzErvyRV7HCePW/Zrfs4LVW1YfjndJj4814
bjOzctknL9+w23OZ61hw5pQBbSuDHxJrhYT6Hxsul5SKhBkfSp6xrEcbOpw6j3fZCLD6nDLYjFO/
0emky6OH66uoYWc8dSN2SSNM2/32NVVR5qyx/TY3i4foWVWYtKrHCPVkS5oih5mEc8bpdj2bafoD
/mmvgpQDTKrGZFV2+igBX1qPUjQgX343mc4orpLellaE+fU1wziIG1td6klz9OvKAF2kJACH2S7B
gJ0K6HkFnWjhM1H9wzPgmhzgxVdV5ZMNqaQtQB8sL69xdqdnOM09rhf3vJ8vJ7QumUryr+fijVro
NhsIJWrQgDnr5pevTYefnm9YxzWahZsPy2Hz16KTpX74UMs9HUjk9e3zuV+wevBvNJNfyZwwYCTF
knsyVndEQQz6Meg+DZyrmZHAwF7nNFe98kaFzEpgMxATLVEnJdmuOHu3dO2t/ODiD1pgBmJc17p6
wm9KeugQIYuWd/M9RtjUfoqFtLWloRFIAtbeftWW1tuOhhIax3xdxNIO2h6rDklARaOBi6upfwzx
7YWpIyTx6n6/V0UsSlcgwzKq+glN/pUrPfRdjItysDB06cyoeeO4+X1rPnEECbmkLS/vKFtc5hJ1
YWzBRGOBCtLo3ZLLRk5w2oxVxH0aFe4Cmx7VVf15bsK4Py6Q/kpCzMxlkuaKVpZzCmrWWpdFxqZk
f304x+ALZNKJsMs0ji9Wl+VH9hwg0tKtdnccM4psxwQnYTqE9cD6APGgKchIBFxKvApLitXcyudg
DbFGq1LHTNc4xzzlQOmdNBgrgMPitS0Nqd+8LuQoy2JQofHOVIF/2w1zLJeJ72yv7u/YEY8Gb84R
lUi984RG3mHh6DIQrZOqlSMdbgCfwb259DAiz1/Zw70mYhKXTX8OnDMDWVpHOAvrMcKkKoUQpaOo
zOd8fZkcYYWp2LtrySUAW6ORXy14JxhGbnQ+F1bwdW2HiAq7vPNZc0fO9roI1oDej3t462vJalOs
Ve5KGlLd5E4YVSwzf6s+zsUl7IcK5vv5dlmv7dFOQgBer9X/KOXxmz7g2qtjB2cEugI50vc/lLl5
h1+ENCcLmdOUXs5YrUc4zz5gVcoi0Dp9V+pzdWZmaKkzaPpNv4481mpObCKBk0l6FSOR89PK0bZf
h300/egHTXzabpRKBEFzx7Z9UW20uWEuw3FHyxqyD9ZGnZFZNMssc6SS0Yfu5Hm6SjbIgu0BT7q9
CXhxNLCfIw8to4wPu2uDownTLLcWOGv/YkRNKcnrzE6y4TmpAhCKYF5BMSRMbHqoXpRNzCLU6z2X
FHa2sNWeYSXc/xnbej88fGT9LUvY3bbH4zbHf/DJbI6k9ZyO1cfdqf2RjncqON2lE4MzC+fyyStr
cYRy+rF3aJv2GJ8rWLeDgoL5E5uxdRf60ljDyNyWoY5U2Rzq64smMjAKoh4A10JUe5c+SyX+qBrI
jnDqPsIjq5YeAdOktlDyfWqSG0j6Su1YnJM+dbLq88glUVvgWrlnP9GWEE1l2yHXKYJAheg08YoT
jDwfneNesCLs3b85euDmSf/wyYc9rPBfChVQvz+n+u6iRwSNDyfMprqLyP6lkmhNlUgNf44Fbcrd
/KH6ICU3vHtkOSAzBLzsesp5R5X98iscvoF+ifIuN0l8w3+R+bxY3eYiSga/EVwXxAbxW6EmtFUA
2XmG4EoQoQwwEDeACIWtoY4Kqf+NBNC+EgLgag1c4CgoaOHM/eKr6V3J60D1SALkuSs0pUniUN4f
Tt5kv0MofN8XOeSMT57pJM4sv7fAYU9Gbd8CJ5oySsFWLm13p0ljTLPIMF53HF5K24iM0cZbwZ1r
BWMn9wNK5u16E11YCUE4ShQiV4pFxRPIvc0PEXkT34aSDBFMGe5ixJllaA1tquLWlR90rfGyYI0r
rr+iu6rs1AHPySzKN6gAJgh/hWjy1Pl12NN0h/JWk0fgVkQonqSJ2tcIBPYWiaKVMQWvpMw1q2Nr
jaWoVVkvCTcgn1dd7pXz2T27pXedkGGprtOnBOMhNTNCmB8SFEb70MdSg9qMawUPNgUmeD06fHCU
gRvXpWwwsB6LWJD66dQeZ9IEpxIPZtre/287u5BJx2YPBlADv98AjDNO0TRr//N/FqLyTunG8pfp
ePjdRqeF/w90mZ1HZSE42hJ7iTpX/pC4gYWqZgpkAzgA4Feez2rZ21beI6XeoVcw7u1lAOBFKA6w
ZKPYoHvYHXp9S0LkXM3KZNYxgVhkS0Ag6V3EDmboKNeD07RQvKVI6BQMFE9TpoDwpd8A75IS3uy5
BKN4TDPAqBr8aNREU7vZQZWjCoiWxPJlAT2/6r/Lxi+NroARFyFIsPVTagrKmSDWcRBxEdSNZ4oR
nKjmJRpDO+82wYWCrdEZnkCzFeJr+Xs1oXiJ3eiyLEFAc8dGqA6NdpQEFQLEhovfa3w0os+oQEB2
L4RqKMYKMlefhE+SirInpsXqZgazairCqKLmP7OoSLDgedK9Cr9S2vNCKkKHVT7Kvv24QH7FFPA5
AZFyXxiJFuvw7Xb0GvYnJ4Gqd7V4McDgkUXfCVL+zaaL6wPh+wC/Z9bB2s3XDK7ajVQE2k2RSbqy
Xd7Lf1LLjC6M3LSqNs6xXyS5UkFYJtdkWakjL72LpbnOaS40e/ty/djcypD5XygJc5oqVp5Y8Qtu
W9/z35pyrErjdBoG4GYQGUtj/clUHk1D9H2xMM5BA3rFRC4Ipki1INrcevdn7cr6dwjY3pL8X8VJ
YgtEBKzXE03Zk0oqEOBey+uQk17gACYgamWxEX8kEkPOevJyY5QNHKCk4hnVsenu9J7eTPzWobE4
IAgkuzklpHyv37212n+sc9My+qB6pji/t6b6Ar2QAGnKiaC8U481cqMV/Cqz1QZ9TjsmQSsueCy2
t3xjEB9W0S4AExfRgw6whK2AKwvC/8Kwvwwlj/f9DAkIoVJ+ef/87aO7r6wDIXtwNM4GFnRO8ULH
dG9q6FiOgurL75w8ZG21nAepIrFnGQ7IrkIVg2Sn8XBq2er1xucS7HaS0eFMYG/LZySYBJXQPgjJ
B+Zy4LQ8yuCPFeYsQxSwxvdBwQUTglG0dq1uLx4PftTg1+i4iXJncuo8lmFXtUnMI5MMWRKkJ6fk
3xtiGXFYQucWrgJMbD/LcHqc3MbRuBHMgFMiHRlKCHtCKWGw/hsNCM1A+qcn/hggwFFvXtdHugxw
r2U7dWXGDO5p5zrtD6RiA4z68O4uDQZ9NbiiJ9L4iWwCjjL57awja+OlHf3lQUWc8Vcs85dW460K
1XWP2/RpeGAaxEbHT0qlezcU1MeG8C9yD237S6yhmqbUXD/kXuAHMlcrJpqaxE6PKcD8kHFzX+KV
rYieZzz3NNEl3qh5vjk8PwlVAhOdDb+Bq3LrSNgtYOB5WTc43p2YBGSZg2og2/3FZv89kJDicAt0
BjDE0XbozLXOgpizJi2hHB275mDkh4+Bl00jrIZl85gEZ8wHd8q5Xrq+saGOwXPMesANg4fFMlO4
ukk9hxmoGwg7dJL4gBPkxGsVJuzq6T8dDRQwBE9QClP/LtDKPtpuWNwhoBx11tF2cRnVzTfuo5bq
M7T6ZBLcDJ45yBE/X2SFa9g53XL5EYy4oqA6pef0HVj9pCBne9tanNXkmw1g+w3Y9a/quBII56M4
0rpUA30oHokWDXh4P/HWL8UWOjzR8S6a3A53w77vp9ibq9L9YOqEq+welTLSYwG3yZRg0xosr9Ed
/xmkzIhAthWBxRiwMNV2tLX1P/DXrax0X1bMQ5z7jUubM3GVEMeVt+c96ZiHGIBdM6m+6mpqN01i
ZOvc8TML1PJED9VZi5/7V8SN5cRCblanQiRA8fu9SlX4O7o822o4bb5+MofDpnxhrLeHxRV9Rj/F
gTye0zjXDXSnIGCONWCazXLsYLERpSwN8EimwHC8zOD8zTXzLTLqEDJ6QcP1ZOvQM8pKuSLGfVy2
jYxZRPjAFDRnf3TQ5Ubgznmu2h1doIhYgvjvFpAqBImRBbDeLLL0XGH+2y41zmER5vBs7ApXKECd
i9vSjce0u9aFy/kGOGRCGo/W66iJfflurm9MmpXH8qfadfl8gejBW1/MzCPzZAVoyzhQ0ExAPc4t
heVh03mmwHMlg7s+I5C+hwc15S3je2MBAdpWCETi972JPbwvlF1jJjDeY1hUBJfzfcIIIwPuNskC
bqkvnSP6ctJCh5Nam+d5kiTaRf7jtvFj5JNcch700Noe+0Xg66GCgfAm2/UN/JxBun+5RENXku8T
W3MKNEZoP8mOrrFaiSnJ40KnctirNlnS0j8cV55E0gAJxy1/8PbZef6ZD0zKR9VJPTvtgS2ZysNF
7UgQ15nZ1c7QXvhdzueDiM5qF9ax/FFwdXihIm8t3G57B9r5wUO5Gf0KGPVVvR8zlXqnBfSOvIPu
aPOljrXKwzArmuO2amljYbNWhoDVvWX76/6AChBv/vkiFDybr0+6Y4ymLWUQsLnBcwW4odUQKqoU
L0A0++DSdXabmlPYn7HipuYDhG13QAH1wljCjLY0fGk3GYaC/lsOiacK1asuw00fvghKZaly2PGH
YwA8iVWL+UCwQi2jvdKUgm0+pKAlGt2kpa/r5xcVcB0jmZ280QAQitZkMA0kEGFTU523WJRfnEFX
DEgnaZX28JJFPyd3gQ2Y87VCFE/lMLd+neq1dLpkIbQ0AudISmHsOz1XPYb1A9mfmZda2qi1Krnm
5zWPYMw0iy+kuptFHmABXxUDjWtRcqFxrwvEYrkqn1CsLa2iyBKgHzKIv8kpYkyjYd7UoLQoEc7A
l4AnHoNzDLi2Z6hsZf9qgX8x9G9YLyVzI+Fxdyoh9vDfC3VyNyfwH91eBrwSvpqhE9sUEj8VHc1e
9k5ThoLni91yXFP2vhYAwcxhZUFPZ9+q5acTaxyFJySHgX4x2wMIoHpBoGGsnkjjfUPOnpiOdRgY
gA2sgr6gfOFCXpTg96WGdgJKhBhqRlG5GvuqCxpdjoUrh4twrH8/gMx7lvz3drwU5beSHLaJdh3O
pblkzKCUL7bQ3d1zvo5cnus41R+M+NjNeXOm/xdXC7kBTsHBkjLA4ElMqzsr5gqDx4166fcLWAel
DdpgBFAdf/U3YAm7B+sKL6Z9wQvD1f7CS9TR1/mEIBa8h/cw2jttyaBsUKcqoWxoOW5wU7u2+GTX
WcYU9ASxnljczunQHF5KDvatWhMWQg7SAgVQrywshShiDmggLlOC+O7f8bAlX0BEoj6iZMQ5SO9b
fSO1S2si13kuhs+xEd0dMERZ1Zu/lGNN2zOZlNCF3WYLsIFPYi+8zMzX9fhPJrbMPuRs1pWHCLCt
dHbCzIIaKKCKzoXb6AQwFJGlKjwgktl0Vh4fZyqNfJRxxmy+vFJy1MOyLPbkBQTReies75MpUk/q
78uJikr/skGdlmUF2f77lYh+YAmvOwpKS8aAqzrnaww4G85A9P83kVZTW4H/H9wvnZdi4Wxiw7Si
NbptPShAcwNHSsujuMRdZnZCI7Mi4mrbMSyOF1My5QQfved4kRan5euGvgfA2IVZRjeLGk27YxO4
VevA8A7Q5eYHxCacVzjEEQoDKmZbkdXTa+CYeWitOcFjQrQfHswOI1p++r7I+jjcOf9Sg2vQbyEi
oONtO/n6FMkOmKxeJp1AJo1M6hDN2gc/21kqz8GloTrjacyrl26nwCWkS6iUHJXwbbp+3TiwQrFw
ybPeF7Xmr3o4hFHYNBRS2L7EhvdF/VydW6H5jACE5o3UKKl9NNONyFd1sUp4ew8Z8ciP7PIVIkSg
qiZkyD5gI4qx0Hx86Uji6fFdTVCHrS2wWL34nMM5cv0jSy0OBgPK/ztOPQZ8nH2C9TQ72ADoRWjB
oRbAOM6ziY7+7tDQj5ODHii1bC7hWmWlTNYJCNDzC1JumpMvx2d91LR34NE6nE3YZKajJlE+JlDM
NXbElviFiX1cLw7GChmtMmwK5edHQVsTRMGgFNHTAO6ikp4eeFwO9EEdKkQ9+elHYVbCwPO9YDs2
emiuTMbWyJfJLJ3pws1akkxuntYfAk2fY/eHGJzZ9QACll5qi1XK5i29QtZy/UkX9+zZowimuG4f
9LxNep5Rh4fLmauAgTdm0SKVgsCJ6wxHVNnZcDbVwET+LtR640igyNSudfRO02Cwc7rjM6ZB6/FH
JzMVaWDIYyEInTsWUWVvR0mNoOoiG0IX6lCqwpXA7ngdM3rCosJ8NUocQ+RzqQrtNiO0lyTHtUfn
eQQbP4FgV3kyC94Eeoa9pWTrNmhBgOEw3ZsnZuV8QjG/BR/lBlBTcNMliHqN9dW7EfrivDkK2PAg
6RXBzd16nf1Q44Mw06go2QRDfOK5slAwiJMKCJdSgBZScqX9cHecfNvBpdscCEtTRFZbHy6uBW6I
E5nJqtKYIyCzMU+D2JTroNZcr5jsK+InpW6kEb1fE9XYAm6jx73xXobYm4QRc/AJ0xKkHLXLiVov
g7uy4+9QPHX+eljc1yxlUvMm8yCEOTA/Q7lBS0gQHNG9g/FJ2+25UbOFaxloxIZNtAlRSpxwOqVv
DIbjLkl9/B8iN9JPKi7zpzx8RFEwnfqq4tfMmc1bsP0wz/3fV3iC8Mb9tS2rtAKpFdcJogrgeFRl
svPB4pg7in253/8Z6wEev0+BX2ii2EcIJhC3NAhTevejoWDmud0NjFxOBZbg6b42/vbugo6FX11Z
oVVeV1bpB6N69PsOj8TNLUtohHDBEkqLyP1Yw8OcP8Pr09wDuR8AG5NqXNW+EQsnFov7lPbl9g7b
63ZHHRBRCuN9qipPNgfYmq7UZHbvedgUskPH414IQZbf01HHp1zyK10QURG3GH7B5Iney69puNm0
EaxHZCtftje3IVdcmDP2K503XXMJOU/atp7UyeZqXK+7OboGe0Rl0/IGd4kEXNkhZZogZEAizoTZ
Kvri85FYQ15ozFAq3nqz+dY3jxZUokn+7wQV9aRgIoJOjT2Ua8MsDgeJdfBilFdpHElJJQUdslpn
Agx6AHKxVvZfxLYhYvAfSgi+LFqnR5e/j1kPyrUXuCDf7EwTsH3f6/ZbLNxVcBvNRznNwYrbZZYI
wv/8rmjuvpnHvRsuQ8VehOKoxtt6aA8SUZWZ8PVx6s5yGryFejzyldyy+LOPUz45FiwW9nkyy4FO
dPRw/qMj13/e6/gAJNl+iKx3rOI7xhi0SrooRLom2Tjbp7W+L18BUH8yXzw9rr3fY7DLcXWjsKxW
hhcRajQYSoEXrrLf7YT5A6irRFpXv8EA3yiO/aErpCTlNTQNdNs0QIIMR2xo3aYF9DhsQoYJndIs
2b6yHtLz7RgU5OXe5IVDl0cIJhyF9BWtpgsjAHr7ILLVQmZBYsth3IrbtzFxSGj8Erh/786g1rHm
64UEDPvRI7hW7AKlLRzvtro4xZq5uQI6Y+mcClUQHnWVRTruyFCQxo2Cz171XfqG/XjuaCS5kWyV
2IMxBOtrPZe7eD7KEmKDQbtbYvujOjU7XrZaKRm9ST5bwe+WWByV/1YZueKcqAE6Dv3nrFgrfEIU
94xUR7Dgy+BQYw1ruur4Ua1uXUjnUuKdZQlT8JL9JCqAmm+NszHXVBPYJYjq2qoqGDGsh+GrAmjn
C0m59gkL68z9Jb7zh3/X1WH+MfRHMzbwzyNB5FOo95Z/ZPXBdT5nyPHUNiOgC2uarHcS/XtURbZp
5hT4RH67AXLh/l4/0qwqUmetoHOLzPDohSofja8g/eWns4coF6ITIKuFKEgynq3VDgQBLw/DDTJK
8kKcxcoivj8JqJOiDC/6q9k8K4X5uW2IbBl8bm2E3leShKzbvRfykwaz9VQmpUvOfDSCnJX2MSS8
dDuhfWD2D/HhEsEcy4biqin6LBAkQfaOWc873feyHl6Ml5cXskRTUOfTO1XHsZXTiz6/TG5xpEmX
/vEdpuVeDmMBdGBkGXuVFcdzS7qkGaqdujP7oip9dTpEV7OiJLOBNLaAbqUgbp3owDry0yW74qm6
QD9Q6fOeJLKN/ZzXr43N8znXS0oLi1KcyaId7fzm6f/8/EY+WjkfhECFUXRNs2Z7VLoY0CSm67qS
4n9UKbMF404vYn2hLM43Oh5l+Pa5zjEueN7qBSujHA9L9d0llQbiH7aDaKV9hQ9pI3h63qrXfodU
Gvl0wlrJBhgEyjIkaO1uZJ7bj6GF2YpC+rTXRuyEq6CjzCxT7Dnom3HdMgL0j08cgQGZS7tJnoPg
HG90ntUO9byuTly4uzdJ0JVJ2LfLTTe8d8WSZfz8qHp0AMbRTzjMcUDPzjoLSHBOu3ji/SzsinUs
7THkJe6DvxP2gAZSksAel4IGO/lZ2mo3qYpTXNUQQBJbElEfyGfU4kMrcm99bC5g4tPPL/dyx6go
Wd7r8A4DWmBNxLgHjdWWB9y3NBIbGPlDv+OQKwLZBs1ES+LsvpPMEZkA+8FIkV5DMPRAywa7AkHM
S0XKbDsS4BIy0krYkz4Fal+6CTlMZcjbnUR3+GfMTmiGaw1zDMMyePuGkARRa2SGYbudDLX2YL2G
Wg+xD+heuMECRGzirIsj+HEy8G3LV7ohsSqOlF92eUT3SyFeN4MaPTTvhbIrP/06v44uX/ioW/kU
KMs6syWo5m/F27nwX7d4rgqcVGz26HvK6VuksgnzMpoF/Owx0XrlLUh+H3jsKIHmnsPRp5Lm76Tp
5yOPP5fiZJtI03syNXetkVFXAmLTO42Tzo2LzHhao7j+rA1C6Rhn9rqNRoXbmrGmD+o5zKggU/e5
U7UVHNaAOpZfirIV4E0Jwenf6JQHOoo3q7mYlc6+bqP4riUIId3Fx4tm2HXunQ7dhWzeSiDohsNh
B9CABWnGCdu3rwDbn3KiCAc0XW50Zdz3g4YBFqxaHAk2s8mspYw5l4l1Bv+HgzQXN+eT4HEmOrsC
VhDJduXEd03ugoct5h8Si6h5nTYOeyGTWHqblQSW3/YCYlkKknlkt1gw2lxI8O9KNUAYK18lZ8Tu
TkK+s3Fk1EVq44aeJoAyJjkv2CG1Wh+2DzRF/OpMXeJnhG6QogghexICea72P/tOlMp5LwmIohUj
Hi+WAZfLfeSln0HMlBZhegO2l41bGNsAgAEUmlBrvZz0SC38is/4UILb6n8EfXOKaI9Pc80OQL1U
LyI4nLPv53FdJd1W2IJegqaicVJc1pLn0i7mABk7b4j/bJB46clrtHjjg7TqN9xq4FIM//MwuqBW
nGbD/nVlTHDmRGq60rBYk8sppcIA6he9tgTDdgqYnWKnGFhGNWI/tcPIb6Nq0ZrPdYFTTHKMEHdU
6CkRHkRFzVszpgD6rXybJIfJQtIAgB6ogyDtLKeLQt+7fz5wovG3ytpUKg+d+WMyF9m90RLUBt+6
p9iaczAcGfx3K42ICHiEHYA/zhQTenH8E8EeL9jCs3qrLWL1M8JANTovq3v8XS1S1Lc6swB1MwHB
koqq3qvUJQHIaLIQEZ7GVKotpruVl5gRyPfbpfX9RC7mcjJ7EjiYt7JC5KqSCVoqJNRHtvRaeAVT
G64T2+73bT1pUGi6XdoeRPhh4S9c9+/VHhfpiFi9D0nciEZ2F4r1YxyP3cadLbAp7AUiYQOQ9Q+s
8XJconzaOV+l9NE9o95vJeFtKatNgfwG/YvNdsRnalM18fBYzz5YvimkZ8VdXdMnM2gJgqCmL8au
vhE7BWYJ3Sv3sAffob4HjXKpln7kzDhxmH+0dD0DLHkvQJi1Rkd1jL+yptlqtX6HxENQoMue+XQy
qgYTnndvC0i1KJMcAtJ3vnTXOvLyrR+caHcFqn1PVbnUJBpPB2oe63DoBsHq85RKyUQLXcrGuzAV
1vmJxDPjIA+ckVidUAJLZMj7OcDuQrPsYieLOBs4CRMYfZtydbJTA8DT9z0w3MtCbUw5X3Ar9J6L
oZUDdOxaQsCQoko0QAVUL8tS/8TplwzNyoh6+l/xQJaIDXiQPF+pAE7bZ5lN9HHkVZdeg4J6pQ3S
I8tyhL3zjnLLu3H2C43iAhXv5X2ZDFY8nxEoh2BxjG+G9+fPN3gx1C1SnWiczLwSwKfEmCoV77KQ
f00SocsHvF/mMzhUYCRuTH4Q95unqO/0shiijivqGOz9cLStogYLi9GzSsAVqYvGTyzhXSzm1bhr
6osYyBhxu+YVpO+ny9nSwq2BuMmC0WVBr/QEqE8XDa+X1GdbMB7gBPeWffKzOkOrSLeZioLs9Ezd
YnET/gwfkU7jDGcyTeaIdGX1pRXMADFy/gTWS6520l5QMWCCo/AnXIEpvsUWlbMtb3nrlTOLqPv9
ZXjd/Lrco8VEL1NMHyI9M/izQO9r8bLZjNzF7JkUaP3OccBb1eMMDPaogoklbHDzDG99Ao5pNCwL
wDLBf2JtuibUNb9mJgr+ejAwAcKUXzw03vbVroQ0ChDuhE2fbyz9FtjbDsk/gC1sCQrtVnLnA53g
frc2pyjpyALiDosXagMOZtP21mKDgu1POM2Scgq3eZjqBeX2zYMkzycGazsFTb75fZ2cfmXy/3Wo
c/9Olh7mDXrBl44ZL+61XOjHiqLXz6W0+M0uJ+ZLJCwcXlNv0pOb46ymjrGsLQvBGDM58JsYEp63
1VDFc1fLNIEC/1hSi4HZXllwH66B3gdl0PKWE6WcYDqg3IN7J4C60dhobLg7WfTKazXOAFZLPZOa
kC7DT7nllLNnK8r7wsZBmkoNpC/nuQvExRHmLDtkqluLOjgJ0XmXdOy95YqZZ0fMfUZNP2DNK8Bt
GKtfaZspvIyMSqCvXe2WrpP3poWbwNHfKTLvmT4NPC4QW5xeV1LvkDNNkiTEeaYYTawVhH8D/zU9
fNI/FA9pXd/OkdUEYeO91Ni8531FJLpgaRlVu0Rc4iBg4bjlIved8GToqAi24xsgim2+btZXGTvy
dzfq4NW0aCehZvn3VvW/tPTl2o3mhCC42t7hvh+XPTYUNILrLncF6ixICOwJnAJsBtN2dNe1tejz
oklLwpdyucCLqSInfRF+KjG82UvPqeMooX0rvkRM6VBQP48UArdMzA71yU/vgb3pwHPrzcHU73i0
poLZycjn74yFu95eciZDkOhmAgtyY/iZ/rNC2ryXbXwVzuRT0NC1i2rxZ9SL94nXlO3/By2FYOfw
OD1IKwgehWcZQkNY/XHNN9dHrgshaAjVS2CCW+MasVrqyJskbmDx8hvJMLmzUINo4eX5Fwvt1Zj7
FuynIPIZ7AsAzYq6ZqlYGlnZ/t8TmZaXPQwA84obOqilVzqYSkWdcpS4Q0BMi7g/CrSc3QIa9Zts
RHL8niBK/L37+hZ4WBJatxeNBTDJ/da1Eb4ReJs9YqbdO5mb+3iynM1gBB9UPa9216L1JWi0nUM1
FS92RPrvtdZZ4copzV4NDu7ux4rrIPrasvplmZ174ESkZw7luSqLp4oG0Nie2sym3fljLaIrudgj
K1flhdLPTRTk8VETXO1M9nsUfOlsvhrPHN0ELKCXrE6J5MO14Uf3eTCQPpFYEuM17rtBDKKxqIs8
VBnteYHK+1kHGRmtOhbCC2MHSIYU9cvmBpJzePAt4AS0KyfOvFFOU9q5uJWKkJTFUuiEICWs7xVe
QeekBxgxKMEP/4k1YOkkzu4Y0Rbb+5wnBR3TEnGCgBCvYf8QULNPIvAJW+X8tkaQBVV/7uuduBi6
SipBuL6N2Z/C9nmrO5RW24vDOz55f1/trk6Pfm04K9Gchq1BJMf94FGSQcOVdPC0Ro52TNaKhqUp
r+nCPhTfdqdrIw/gy0ncSC0mJ7SQfs6AXXJbgoBHvfFgwg7L7FuFc2iFLgiF6dTkA5781XpVDwZN
PteMHwDOugh5XREXTHUd7xAz7HW+/UuW16c3Sbt4/+IABoy88JW8Vg+XUUDFibWksbI3EJJhMbym
i/wrhFJvuthV5pkaR7dDcAddJMSt+PnnMnkURU9P4H7CcnqBkxGwmBmZRyISuG+RTfiuauRNqH/m
rZv2/WK+7/JcKJDcV5NmUlLO+33xkyLkCcj5dHxRoryCALuVMsR3Edjgyt/cOIgB20c8FTRQsQO5
hPdlnNlQI46kR7zSHjQzg0GUAzEPj05rJTYpkL8WWkZSTJRh+xErEjqYxfvF9pwvp0MyL/U7wvry
BNxDYy1fN3g4j2s/S13OJpzynMrDTiwcQgLYPb0PlzqS+z9YVpRjlb5IOHWhURVsNwuRF56LRZpD
AWVxEWM8ZmwyANH1hlMHOSTFZb1G2bnLnXc+3GPbqOrpot/QQZtp2kbhlHF9y4T3MYPE5W+rTii4
ZVvUadK0goa6tF4ZNkhu8Z6ei9P2C6eGefm2WBfRjVTgpHNcaHHV0qt0GO1XzSVoNJwdSuPRBRHy
6HfPWKcaaOfosMXx4wCO1iG01SaGwwTN726IsCnVSSnUDgr+ZqslSLq9dBKVvp4hYDcG7DmChExv
FnLvluJYgdEnXZI/0QgkXaihS9AnZ77t4cXnAg2Q/G6+emY/kTfeNPx9jfck2uvlCCDoEFPkbITK
o6OtK27A851kJ8WFG8rlTHBSvUugunQUPpirYWCsP7tFI5UWWWs8skdKAUxKRNGEdIEQA8ZuuhQz
MgTf6XMuXCHJ2S+xZPu+0Gcv4P489nD54odXyywJImJg6RKW6KlQF0dlE9uUIzZ20OFj8tfoPs79
Ux4QjAgBzcVvPZi0K1bxRpLm74NrNMb7a69fCgmlRt/z4S9EzzS8JjQZ9RM56cp3D4YaYfv1grHU
uH1lemvLQqTTdZ2X263ynzx5kl2yGcEOv2oZ7pzXfTLXREFWPBYTQ2hFT9oDM+WyYo8P2cTAsdFq
mwk7HpOqJ9kOJAkjvCGADuxzWjaHoeg3VLYm/5jGFDy/PEHpMO+lsZALZG3BIMVUVVZYJrg3ujoB
SI3Xhu8WWMyjAaJBsnytI3uEwbgIk8ZAL7cvcsKxgvW+TQM9nmV5PQquuCZ2L1k3F9mV3bm6wRzC
zBWtDQRGODV7qlL6z6mh6OKRz3xtDrX4x95m+vR84dyL9hVKQWFm0hfPmBd/WLGwbA5+olhfwUJ5
rce5TTNr60qzQYUraCzgy55sGwFTX/c0nNSSx0AYzC0fSLmIWIPVp6itx7UCb2UgOPNQ5vRvXYj2
bSZSXJD2sIpqusgM0OppgVYojc6KhL/a/PXO5bhDnGuj+uRKqnomy8+WXNt8YQqmucvN+pa4Rdm+
tRomttzHPP9ejHJIqOQB3zPtkhdL4d9qRydrc7zJH7KagSc50oMw9Q8HAftbqABIfcvRy2N5KhPR
feKfHZc+d26CFuOzrOwou1LNY5dtDAqxUo3qcMIONZEMFSKkxg3N+IVNYbtUFILf1aKMerv20Vnb
Pio1ycT6C+mZne+1+Zik59/2X1gQ9v4efty8Bm8qVUZpzIHA60wCQZaQe7jy3lhd2AdDmAIR62Cz
cZb0tCXEbcwdWCxGsKDl7gD8qInHLQoLBjn7RIs8/FApSACzVj3NvGhecWyCWzA5uIwIk+2WcqIM
nKcxa0Zm1q21MQvXF3KTECtNDZb8rm0qXKMnRBegblPmXSfm6HoRIqWHk1+YZtEfqBmhDHuFM4wT
W0IZ2M2ftwd8KJzC7NUS7y3TnPb07ZflZ4ZE2PXYndRr8udZS691U2cUHr1Zgnfm0ltgFMyJFcDz
8Tg/TWJEVlw3ssG/LQ+sNZ27pl+thGUuo2sKbWKCYNtL1FFJq/RIvjmxue/ZqeYxwW81Syhe1OEn
ol+n26UooJGyA486rohV3SM/o+Y9R08xtPB9ajMl5vDae92vO7/Tr1tYgIPVz8lGE/GLyb2FcrDQ
mkCM1ibYsEdqNHpf49jLD+xgTSLp6z6nFvFrEBsU8lC2YDQ4k/9vIXuP3yUvBBNv391QzoA7Buz9
bNiLrmjRF3o9tj+pGgPGNSSy5fvQ/C2Fpj7V0E0qWayMHSW6LfhIaR39EcPMxVW8p0iIRxi6EYzC
Prkf/HK5DKLEAUg7ce4O25HC41+YanV+VX5LL47sZcBaGt8V8b73oqCjeBf8Kwoem2/g5M84s5TK
k1owb9YdilDsLSCUdyNnZlYBpuYESJWT1EsgfwlZgr8mzhtC5RpMSrFvoDFsUqNnm4zBmWBc+O/+
xgojoJz3+eWOZoMHeqzLHGKbLqpQnU7dOEZKHPHI3w6E2XvNGIV+tbKGhTvhHAISZ4k94dYdxDGV
GekQCf/zQWAz1ucMLQwmcDswJ9X0zHwz0jNvyTi4M99iSL0BOlUfuLQhMQDdPJBvE0HhIjEMc0oL
Kl6WHVPVP+GJ7DgLq8CJigXha1wAjZoBz4uzFlPTBVF7fnT/Y/qEzAte7//B5OPofsxh7yzbuVZk
i2jPJr5gmPKv191VqfAwoVqBAnh1g+ZSt39+EukUcQt68bNAZJh+ixim0Jjzyf8BIaoo++MXdV6L
GLWkL+Y1W8M25n9pYfkv58AEtfP4/Un7GD1ZxibS4K04bV2cGTmwEW5lbKIcAop0X1bWNeiilAq+
CVRDUbxFi2AN8a+qJ9Ern3CEP7RxX0Y8yTQlOdgrSSMpA8pKSBn+ZOv3nZt59hBtnfl3oBcARwre
4AIzgvNWpWsFd7Q4iOSVql4st8NNXDP1a10JsMl4KyE826So9TzWKOt8rto9Um+L5flHyIQNpf+Q
4P0Z/sJz5LK9sKtgBDVcCdPQDhhIoxnpYtisr0wfyz8Rw7v606glifYTUOCDAn52xjF7vx11Y0U4
k5mIgMJPo+9IoPsHKcaiNxy6bQqs1PqXhHbPEVKDVXngD9fSpvZPRpVmqznXprWuTXS1mv/6/lNF
+xAzpEg/JMzAK7HkHx7LFi6aEQ2IOmCLU0BTKyJPoJixJYQO5Xhruvx7q1AXT6dEX0CsF26xN6rr
krvc1U2mKNqbeSWG9TBN8jiw8yuxdPkQLdIYX2mJWvEoW0mrTC/cCmEtnVBUZ1gcCzNvCa3rY8uy
EGU0lSpu/9A+W4BmUxeZJpd/OgpkF3adJz+EY/rW45ZPh9kEj/9fkVK0YwvbaqPpN9OVTGf5N1yz
AfmJ0Q/rJVGdwUkumGxPwaF/k8o8LshrcY0CefVj9KrrHO+QdsEwxkROIk5euw9gqjIrcAVNcIeA
ujiD+3EXRDc5utsCR8jEyDG4TqvM0VpQDHA8fNWI1VuE17qStPQpTssXPjlPidTdJ43y+yIhE6l7
v97QBnK36dKQgI8XefpsiBPft+R1MBEB35zNrSx5bNc+BSvcNJ+eCoReUCjekWM05thb7h+V+9sM
cd3DCwhgGZcFquzva2yH7FKlK725jZ49/yJvpr8GF9oRPWKKUFKb1XgpLXLadE/R9o/OU8QLnpPQ
7xJpKi2XefzdpIMME0LVFR0Qo+uVrCIdGl1+8Pgrphbtq8HcPrJVtIJkA8kKL5I7nc8uctD1LRh/
7HMOTahUD6g5ttGY97D0fuFp2N2I4BRUmZRw6GtW8U0c1m206uRvs1DxE2uKummh3tllLf7v+IgQ
4zUn3qHniGHZ9Nx73KYTr1YENl3rGiCom/bIFZWdiLHVhlKeKVwR42e89iPf6fSBtE3YjC3JxbF3
vHcob8vWmlw2C2yGcRaoLGhRac1mv40LFhMB60G6hglf7DqLKCi6AOLpD7HwaOLvs3je15f6NvFc
T41weyDHKB3NFeYGyHuykrG/WB00Wxd5W+71WUNVUVkgkZva7p1UpLY/iQem17YFR1Cpg9BeHCP2
c1mjO7pUW6vdVV9NGwfPSNiAZs64+K7Tdycok3sVCbm2RNkpMT462xjO475DkkWeTJWTOz+oe1cy
YIMVSj0bkGQmclp113Xw9AKZ2Ex8JePQ8GC0UFn2VivMu1emCY9IM2PGhxcJ1ECUHPyOlbe9ZmrZ
9ZSXQsF2Be4BL5oqTphA1NP+pcPskg9Z4D0YmjVf1MIrVZLV0uyuT05wZgs3D+aq0spUqdodTIBD
2kwkA01B14toZBYqtLA/x0WvukU/y/WU2pB+9JuFaGx580nLP6ruTOAkOthHvpFYn50cLR6O8mZC
IrHKfB/2qJeSO7OjsUxKg4CoPUUwQjZgJDR00Y1jrD5NP1L880el6OG/5ZEy05shswPDR0bMA8TI
TLULV2fwxuOH9p4guxG/sVYeHg4H7aUznQ+rpcbrWhldYwMbMBGd0cJLXgO6uDfFOchLnIzJnBQ/
zro2uKTREwneBLtzryOHFo9fgTcbC1RJ/cU32e3tuwNFE4ihx0PyyC91Xuh0b/FTXZ2uwRTEpkPd
UDWSydzTa9Q6M3N8AI6fT2/mN8CPHkspRUDAaIZfTB9fzbOYxm7wyLmEtdMSMRLRCjJlKWROIeYb
XxUU6cNqnSUp5WBINqh77hYgsXTOudSRGMenNHgjANnH/UIaf0yBVtMseA4dmqjGbkBascNgF6k3
RDEJ6j5xMysvD86jluDPc9Xw5596MQ1WRnciZtebZWFZoNVev/CaKJzAbWnkeex86w+usqGtcert
MNVsGLF9H/77Bzd4OYoe/9MuYq2xhmy3xwpyaJxKUEgTt6W3qmtHgy9PAF//Sh9d6HPp18eKpbYX
yDtimDHN1dPAJVIVSjX9kfIlSFq65VWn8CP2lywMFl3G1e62B3iUvsUGt9g1W7AzrK54JJ4hKwJm
h87OBumJXMk6E1Zj3txo/ZXseJWsFasORH5t47/yxROTBDA+OpPU50bKJsRKxSVHNztGOzXDHY0+
/9zpdxYzhkB+B5jrm4ouf9Btjm/H87q2I1V42M0rltKQCgaxJnYZl4Ml4/QOf4vXjmIo9FGxaTtn
xgspZKnTxDEg3tRzNXpYSFOqV+qGg3+++7YyKpSb+Jh9NLHeRUS1YZpi/GzwEOttp7bzskgyUpud
eZ/2MP+jtBCZ3Vcg/i0ALYbRHu1lnJ8U+kosFginTeNzaFZmjCvQl0i9IjsrVDGFLODRt0akHMss
/bqFDtOwwW6tqLPCWVAisxZaUzxSfkEn42u2MYhOs4DC1GRYoT1CW5NG3mQEFk7Hcb8lart1Pqgd
hVDHvGLmjGFy1+Ehtmf6S6fZP7gRebMVg+ePdLlhgNm9WAy6Djv0LUX35lzwMvWAqbSepGi2f9Sh
KKHG4VjzHJFTS/sbeF8iZrKA7fwfzhu5tsbVdHTZzvgwkj6L6o3HRNMhOL64afqF4Uwu75rsHHWV
8vA/t2JEYaqqxTE/IYfpszc5+WdVLDhVkz9aQfLStJ32ABrWgDM2ZIP9cKplbasBlsj9bTbBf/sJ
CuzfZzB/bwCjzAmUdR0mHbCzTUo4sALAM9DQte9C6wKwyLvX0NKmEvfzYtcifEU9ySE02i2cDchw
voOQM68Piv93p4sstAerjYXBRwiHV6Hzb/DZQxtlkiWe91JQqGUecaf3cdc3q+Yyv7FMLs85baWD
DVNi9ZptVWDOCepS9SDoxX1wDYEv7SnWN5B5EJ29YN6wYPYZd7AaTrJST790E8DUQDM/uRmrk03I
texuSP/MPI7pz1+8qABtg9exvy2DKp5+GjyiW06t8zzmC61Z0pDAUKVcmt/dRSiU4xqUmOdIh49b
sdtdfa2jQ34pFtW2uAYPcjjB9EgAmPcvcgbVjzsdySj8g2oUw9raJO1pzNMYG7uEKlBXrebPtZvM
HKImhr9nOx+TIf9sS0eKnyHjSPCO2McxtSQtpX7SO7tSf/LyfOWCOgWE+DZ0/OuX7P04DlBxUWTH
EdDYOVZt0Xogx8yWD9RCptbvskH86jHY6UGt5RjmPrIGZ0LaAyeDL+Imct2k6G33QxUThiVbkDVU
mjkz/TI633JAqD7EsALMP7eviLbJwnay+yoCU1UZj6Xi7oK4++sQtRlANKu/soh7s3Xnl4MIeVGH
YOPIq6e7kyvq5XMccqmBSg43EUHw+tRFpc3LTMIVczW6Qy1bvdO6ZQrLPxPo0bXH8EswIChB1Ges
DK12ytnyHMmIf1XjQmDowycAJ1HbzqeRgIQD/4QMyH+ilSzzqXLcX8erYhqFPSUMiiYoayEW5x7t
xrBZsQ0WZAcrxbTY4PPoeCarKVPboSF1veA6hwdL4igkZ5XCFJCW2H5m13+8oOT2f5RlgWessEzH
FLNygNxFnnPfCTuYqgMEeOSevbKV4zLf4qaews25jQmkmMVZZ0bJ+ewklmMmOPaqapunfCkXIlB4
VwdAj9y+cX02vm5JBOX2DlQf1LgiFdRDmRsZEls97zkUHVd0tsKqBtKLL93IkJM7oMQMa7NxTYdD
ss8/bj+6sd5Szx17IaTrJOpBPciYUD/XiI45pil6Jz8wzGkkq7oxK7wiBvwMvdC0lXc/PwrhAz7k
vCdg8YyVwSY6+U7VhMPw8i7964mPuVvR/89AJNBDlEovDoBa751Ndeenmqew+s4yXwEJIXkhqQnm
tr+rlz4HMWNY1ayuPmKeidPJshVV/PBKG95jPHpi+mXZIB3ZWZefKXvGJaUblmOZp4+QmaVkNTOC
xitb2vrn63VAjf4WNq0B6C/9kx8AuMJCO65slQHWh7YxOzQusQxyWXJT1S8Qo6ySoHB2LgPjcdUo
MeaSRZewlpQ0HvZYn8onHBUjhmH/zeT/lUjoYmyTiO15OSxYeBSZ9bThQXakHEfW/oOrt2HjxORa
J4+IJLScVpQhvXrm+5LI33b5M1G42qlOb3UJtJ7xuW4s7Obby15v7vpuIPmXcL7aQyhmznCj4f6R
9WV3WSz0A2mcZkS8meMNP5TturrBGR+rlgCO8R0kAousUZsxxtSrOzrYvKCG3rnZdsLvTSs76crw
4dSk8c6R2VAsH3RFNsOWz/xllMV4TQfyhRFjfH0HS8rDYJinL0Z1tKyXiFCGvIyvXGrZJy9oMpiX
uMdu7PH3uOxSCLqogk+XwP8ZXzPfwXnwcywFZ1+k9PAyPbLtvTuRB3a9pAmNEGCiLD6wct62AAS6
fRAXIe+nX9QL1Uj9qgygojWV54lLVx5U5Kh+/19y3Ub8ihinUhnmsE+/4ObQFRab/kHNwv2koz1b
AsOU88VD6LJb3wfTkHaNK26EdpLaolKc05GAlarN6MmZuRqSkdCe8T1jvwxNv3/2BHzi+iZz9cuB
+PO/Fwjx6JX/mWBKHPo8Fc5Dnj6Yz01rsGfyAXYO4QXysm5dmnBxfxPpWOAJ2VEUqvK6UP/QSE/K
P8wkMHGNuYwD4qgvL2woczNK+7D8dtE7pF3ob3402G6+GydNOCj07kmgmqM++sC6wILs8i3XhVXx
NUGQQOldG+zQnh1PbMgSeqCsYTBoELSg1ia2QS/xHW480AsOJU2TYHhMzzSe+tGnqEMOuCbBtaQz
UekSFnYaNGrAj0wp8LUr/BdCnt8zVAw+Ktqzo1EvzUaOfwFPAnzWiVx4VDRJaKrdDl4tnxmc2c95
k5ef/S21cQgeqrfkHJB1jYeFwWVL9cj0GogC8cHVWdTF8wxscpQz/IDIJhGE5XfhAvsastcYJY2t
nIEYUAsMPoRgz8jT4q6vXyBpKWPodn0HCOEmFYLBnczo9lDo7vOHhPCQe1Gn7En4qbqkyzUKTZVq
7XN1gp2yFVlnM/ZP4S3PvknSBSP037U1VKdfi5XBjYanRzBov3MEvnWAiPxbjR16kYEIrlOsOXa2
bHX/MjOb/IStY+5AVEZIS4djh0fHLF2iypQL+Q+P6+pbmVPrI7lWRvdInhzs38plOJBOllWfkeUI
UHQfp7aaIbewU2nveJlzEkBoBiW8XWo9ltHU3+X7Sdjh13F9YLDUOfp0t4a1eToYPqNe8yIu5mC3
cspCqnhNyYFMTWi7Gsk7MpXZ5oAgYjt3E5Ijek3bMb9Ig2d6NFUwHhcc6xz13yse8OqadjIEZx86
In6G/Uwa+YZPhinlknpAn3r9AADAMvqKrYN2XhioRXZmd8fsBeNtfU6Yb51ti+hMdcqCxvaKqMEw
ulN3AYQkXcVCnE58NlTWJmsfJ3gLUY5ZphsgZGptENCZQi+v8bkJYh/SJOfcEBFJMCU4q/P7tyVS
yBZ5CHtDHEEvDLsoExIdJF1sefN8mzwsx+FeKqxpyTPDsd85TBNHB5f/Oh3t6gB8rxIyF63uTzBv
SCYmyZbCXGI8SWwfENnlW43RDo56+ko6i2IFSUvSpw+4xx5+wFUbUfTG30obvy5amzXcglplcmg+
3k3KL6bZmNhHrciod/KxUkT5JCKQzX+JUc6CsmISyfuwTPwzNkxExj5lvGkime+ntUh67zGzVVBj
ddxmnPaHI9f29YUmGwMKYe1K0I0O4SeCnqnubKX4umR0Poi1YR1PDaBAwZ5AzbE+gRU0Q3JDt1Y0
EhCTohABkna32d2yROhTRzz7WAmLaz++ATrHKjFc+Jb8OT9AcJFea7iPBeDslrHqgLgNfD/BegBi
PjuOtsV518H3khBiRS9x+IaffEHA8axMJrsTaIydodZp/xiAEJWhHHfsjcTkm760w90z1CSuPY5W
/p9deSnP+7n7hD7DQ0IjtWqrizzWguwDOssqIPE5Pl6aQUQIwOYflcU4umnyRtQF1QrLhACwsEbQ
F1EtNd0C+C1iu2i3jEeITAQOBk9LTk84IlD2ievZ2kRjaPVt/A/qSgDqWfiCx12EmCyld32P2DZl
GvJAV9v6dcd4go39cw9OeirQX6/2gohNcoTOQ5dJXebaykkXZzAe2uVpswzGZrtAICC1hwCGGsJM
ZsQaanZVWCZchGvjk5BhzDMTFdOZzbwdHA7EKuNpv589PsfDhrFkZWnZ4ERoLb77oyXPvvwuKtPO
vfho/oa0EiXAFv44G6n3ALxPNTv+gRYxRgl1Y8YTZQXJseUyQsU1SVujUsfYZP/mbXifA0koYMO0
SGowHgiTulndEf3XzSxifS62/ey3r93RDB8VG+6zGSCQoZ8YKq1rj8j7bnkwtR+YDAiNZE733uhF
YcNq3FqHRTxa09krnraueYCFA81U0eqLrofjwTt4dzqPTArBFSgGk4BNnQ9qLSmnICggO6YeBqux
uKNvB0jq34v44Ist5WWeAUOJzM3VeLyhTMJkI91iUKfxiaGxDxbuIus/iI5ag/i1LwVoVM4earA7
FDgF4VuUYL/Tnhx1a5KITMdN6d1sfcOkkp3+NuS2FklSZjoeijjnm8Hv8ZbkGdFRPHkx7Q1PYdOx
ejflWc3omaLLD5XL3i2jv6BnCiQFZx0SOuArmjP38aT/7B7zMwPr1l7I7RV3Iy2fjnF/stlVHnAW
bREfIFM+T9UaD5HM3yd7OVU1HiGVRNeQsuCaGLntYDZJhv2lU6VWA9GC/rTH8ew3WDFokW6oJOSK
Xzr8k7t6gP2zmwRBy/Mh5zFJ6Mbyi7BhRbHUgVPJPQve+hZDTMuA3cBnASxKuETP9XnyBtP8SCzB
kj1uVzA/qmuxYsrSgELVuydmj5GA5T29SLa1QHoDVeQPEJu7uzNVEexEUR/KOgky14CNLSmwedSD
mw4Qo7e+7fb/XNFN6F8psLlQIHccNCQ2m+eD7Ol5NG9pdqBBi7eq/gIejO3MJLXQraw+D2VcyRJV
cZSrZcmWLYTi4TxIwouSIjsn9UoFyZhsov8GjUFf85C1wbtTOWX3SFTFr4Y4hd7ER8pWlaI6LiQh
MxfieWzoWQt5k+RoW3R59XFaTgkl0YMeD2BvmkEOO6Z8bc0r9HYZX3xqAc8IQC/fabYLpCNoQh71
DYfWfIiXZiJuoezANZ0BV0zmgWyGnk/OfqYVbGsOVLvUw++7pwD/soMOntmwgRHkzZ152NDRcche
YI0IIDrEIcsouncYzxxDu6Lv0o7GMGTZIh6J5TaJU1n/lIkQqxLYVautJw2y7uOZEybS8jG1eHUO
KNasZvFO8vCj1ZubA/IRfLwn9kDMmvL8JWPirGkpZJ2b6W7QbqIgk+fL2H4y0P4YTshYvC4bWObY
L8di3DAwbqrL4iUOQIVZFMJqOxapNpbCLTTd5ZSa+ssWz5fT/S0VkdlKAY5bWNGpvGcPv5Tj9usj
GZRbsNEp2fy/mlmNDwBQ5DhWjWnnz4QDoApC9JKy4Y9FmuatYfBZNn560NoS+9OK8unO/VUT7sfQ
8l8UTwtJ03cR1KtqbrttwrBQfLMPR7HalfbJNl0ciT6nf6wFECHmF4qXVDTstXD/GM7laS0NHiZs
xYdCCFEupyAMF1L0VbvrDYPKad7i59F1pp821USaecesw6qX7AZpz3BjTaAvDtSOyVPpWKKV+Z2P
MET2G7fmNSlww9o7+GMJeWSlh0SVX7JikQYvdpqajO84EyOwaAhHBqBZ9a2Po3X/IBVJspfkWfye
kPrUsj3d44JO8eDk+suReiWe59ZfOdtOv4JGWGTELiMD61DhytBXRS+orVLKxe3cegUvcAgLz/Y4
IF6O8raW7EktC+HZsp1UhRNSXYjYOfmatBrBSUi+kGlloF/lrJneiKdRjAKxvsRnUFA18TDHE2jY
8iv0h8DehnV1hYGjiVmUVgDC1z3aGit6FxQJ/KcMg6AhJ8nmPd0035+nWYkJDhcM2LlG+wReKIBe
xyV3S9sTBwOrFd1uZmHUwvCmUwFWwUfqCc/OzZ8yZbkjoSW4tHfeHbWG9OXICGBgcuSXrkuXih9y
xIhwxpiDP5vJY3ldt5dLnldqMgou86y9xa5KW4oHqsx4fUV8H37anv0jrEOWReJVD4QdKAlucPHd
NjXo0aSSPLP3JP7ubNjfypMxmDmxkKSVqVjCUx605XhYsgK6hwHuy/h0/1RHpzKJu7947TmBd+TJ
Bl/wenKpi1+tyLwn5WO0t9MeVwIpfmOPIlSWS+3wFN4QnjtfLpJOFevWzR0spCfIk2QLjETnf6eY
lDlhOllfLm48oTZGDcdBKYidbnq4TaKuWopyhEuY5k0UmuTBLfbAqynxh7PYudbdjaHPOYiUdFH7
ActUA57Y5RqZx4VZddcIXh59YAjfvUQdCSj/tRvmewOovUrFXszQ2uI4oTW0ziehNTRNHvUIlsr0
r/rcoEJFVmXLN/+27+0OuAQYU+7MbhSJGHz6t0SXn+/oRmuFM3gMqSBQa8uzgaNB2y14+YBPBR1x
pUqwVje2V+TdGmhN0D0r4tFNGrnIZ8AMLeVSg2rNc1fm+exIvTbRTuAetl4Wtq70McAg/6xswKhe
IuOV6L2LkyitdN7kt3lWwJy5IUSVYRMh3mw0dgnjL0qiJKlENcaQXBG6A69bTpybAne44GqgeZ+b
ph/821MgPxo8Rhje3QLkw+MBRryUYYZcE19hM4IQX6tlo05RuI/36EuSd21bEm+qWJJIvoUvaff0
Ebn47XxSG9IeA0qVgv9hvKqJf2w4Cam3Mp/35SCE6KoDfeLfWES+PlUDRU1xwDB0FqJ/0+Oy6E0T
O/qq90/e4XdhQNlvHOSuhVKJDEyZKFC0Zfyu65nkXgx2G7psKHlzCANMysTR4I15YXcjt+yLQ7zq
JvSVNyXxfSnqYXlz0/2Gw2c1BzyuiKlCos2RRgdS3ypDYvsb2Dasf34+3MKO31UeB7fMKyrkuzeQ
YCbY9sF8ccpE2iAOP4vChoyPQcGPfsNQLzPGWxoOdX236HqrKlCSOga5uoGWQxn5plkwOKPOACfx
nJJo/MmByhNWmrzZg6hQ8YPcRjPsuSw+dhrv3LKaMArrx/432cclS0OySr5CFfwPV3FE7zFtsEF/
g475ixJ7avKBPAxDAXwJuDb7AeoF0bFthpzFA6iF2FvNykAm7NWCZ9rfCmgmrl86KIbEVC/UZ6cy
T3eG9Jg7YXgjwF28ZMC9Sw+rG+XtTj7EoZWWsQ7dnpr9NX+PTyxvxzlIph6DXGjSJUcHSA/6+wO2
3iajqKV5aGYI5rPPuITRIf6iIH1DoE72T/8L7pRov1r1tuq/aJRxSp1ZlneBYqk+Gclyl5ktEK8Q
0f6InBN8JKrJ9hsTXDwzNmYv5hLBnUFBuhgw5D+yKo25nOrBH2tjwIY3X9iZqefxnb/4nfeeFZ8W
JnACv6LocrZeghxaoat6WB4iv5lfbu40pPIm9zlRiemADmL3K2GzGFsvwUXcT+RaPXGm0QRaKX9D
T6BXWxLscwASND33CvE3OokPhrt2vX0fbC1lffpnqEcQU/IqVBPoDQQEPBZceeolFlGKv38RI2YX
siqFUjB/5d1CVq3BuuiC+XanR4/K2nFpJjtTWoifvMeKKxUfuCVBDGi7kNj4CAbFb00H2YIgRVDD
nyatb6XeUDpbck+2kQar/PW5evan38Y4mzmpGshuH9na67nhEktMg7Htg1CN3Cl0sHIpikc48283
jC8/NL4VDBs+nBY2Fw6YIYcYx5P8QccSA2eQTxm2bW1yU3QTqCcHZW1cxc0TmzGlx+REM8oAa7+o
It3nhGQM+/sP2nc7J/7TBzR7ZcKyExPerdwboDEZTRQ7BPqnztkzHhkT3MhUBdwkpw0d0lV4QfyL
9GGatpUE2X91x5sHD2aNEt9Agw1ygjJXBm268k+9RbpnijBFO06Z+tpfvCidmIRd3d8d7HupKjIR
FtZXVzeGkNRZZ2M/v4+xzrLdQNYvj19p8qO/AWtS2wcFUO2L1ZURGkkHFFJ+Aqs9XCRLt33w/nPF
viYCjdiDV7VipXo4bEvkw9FvhboSAJSNplkc2Y4Oz7lVVgTlCoDLUoIyPqQRHp3IS6pig99milO5
RPw/VxhADKEDlrjlA+q6QLBZ7zLHG3bYEDxqE38mQX1L8UwOUNXT3/gFDfwfnh5FbfGHsvwivHJk
R/Z4w2ReC0u/I6wuvFs0daSAOwUnnQ5d49QURGLZpjf0hQNGBVEPObujPQH0m+DQTXj3icKxTJlE
XOyQ2CfguYFV5vZlXTQiGWQ/lHw4m3hyrU6J+g6MIylZ3NsoE47txuuFbywpWjRYMbUkIMNhBAwM
ChMdgPfI+N7Pz01AsYJD4Q5qlivDhF58gsUeUcwPPRG2BE+SzvwnKUDlFVv3RtVHpbbmkNPkUz/v
Py/xAM+WLM31Vg/43mZQEoHb2/tX+Pvd2h9a12805S1FOxzh4Gqon61ewbuwTlUwUybmEMRq6Fcy
FA1LBGI6U0WqXjy86+lWlmJPZP4Xy+R84Ae/vjtEivpi53UjHN2EjQFz8+n8EaqfJR3FMVf9CjBv
NT5A1ltvMTdPbpQTKnrjWA9icyNVVoXqHjwBoNQYM/dL+WHVc5nGVfhZvR1XEUCStIwIANyj8NmF
bS9+CUzImVH6DgRfiQmqaNzeBgCVFbp2lW7m8NH4IoTpyPh6o4aR2edAeduTx49ot8DhsNOARNmm
tymLeL/yLZsYYCzGV5TQ5cczeCI1q2S9bf8yJh6x/2F9IE456zkR52Jwe9l2sQWOpgQtdPv1Pv3j
blTzM6vIjkzdrU0zqRil6XIGySNdz5rKfGl1anPIaXzJNWZO2Un/KAjxjLEn5IktpG1ASYO62raU
AVFU+NNX/1GPANRpjMlG2ggCxRu8cifIhhAUXpqO+JTuE8DDvT/BDIiXnjkCd6UpHjx3kQ86soHt
juR2t1tju2YtyCsgdn6Y06M3fSSBjUpgEI68SG1DVgx++huGU1rPRytKd6INzE0izjoQjVKFSAuz
tkv4HS/kHU5rw7U84iz5is4m5AQgRKfrA8PdviLsWx37cw2KXj7SyIzid3D2XFmyAloZklaCheWF
DH/4t3Wl/jjiCHWWP32ZkowIVn40lJiebVmvU9sQKf6sI0WUhO4iqxrfquTzmAjgQrmqQ0z23ydg
ofNtQwdFcuImZGyV2yRps6jL/1dFWcrCPJKwlxi0yoYOaMAmcNnjK2WZRenVTDJ0w07Aa1nWKers
Ns6+a41blsAN7MXGPxOjUPJ5m1vDFsQX6ofixzq5OA42umR5CfnlG/7XTiToe2CuXkhceVH7WJSf
SSpu403D1nkSXTzi8DfvMPielVcvGBVISyXf3gt6mB8Um4xuMKBibq0AeHxmpRuR/V5PhiqAXAu4
aDkJf83cLiHKlT7jIcdQ0tuPxvDGDzXA69Hcylu2g2mvqqDB2Ck0n7GQlHOOE0xRw/HI78N6uSML
5hyb3eTc+a4tYf+kcwKS1d0Cv3OTGW4Yl7RwqEPqitGkAbA2hdemR89PDBO3sFGy7zi7JCZHHh0c
tZVvPuhCzHv77t1B/GliHGRf9a1facR/2S4Ljj8vYrKwSt4a1yXy8dp6o5gOuF4RY7E8LbUL9iJx
S8VYL0hsPeoqdHbA0L15B/SdFoi5nFjwKTK4HOYwGC+QQnvGsSPLx8RnLtn2Pp+kZ38xQEoGQqjD
uiBMuXvZiDpThGZn5Yd1zBNm9EmSDIkuOPUhuDH9rjxLmUrK319FxYF625Sh5d/OL02//Fy4SPqW
GWnLpIfjm5ZdAq1YaF/N/djkLgljWn9rKt7Z+lz7iZ8x3TYIHbTqCmpjpx2d2Iy9sYR7pXOSedU8
2TFYJ2x0IIDVR2DhJA8obBJj3yBJEEn+KaYMEDOXSQmSz2KAmIQMxW0uXjLJKlCjwf9H7oWLBBsO
cC6r0ooiiKeCkpxSx/2zbb875Sg7qoxFuv/TaxGtBNucjM5v31Rous838Ia7QEByIN3U5QFbgzGO
SYwJrWWj8k+OaA26NFReGeFA6UYLaxRmlDRmJwyxrQw4LpzGiihl3Al8VyXL0yidqMTgp3x7ccvL
8k466Wr8QkxrPvIkPaXw5dUq6AFfSqMGjB41vBNqGKRJqK4odUA+RugH2OBVxGaMl9bXa0l8lNYr
pq4h+vfGSQsA7PeE/9pDcKVTvndc58hmBJknoPry7U1D4JDCZC25oCIHQlOc/zn4MPuWIQv+xXgm
cGkYI69Femded/LwpQ5lLP5kP6V9gNCecsFhWCgH2A++iY9e0Q8nbTgQzuCyRcQ3xIwdK3pAl6PN
gIB4e8qPGq6LwAxE4OZa2aCTkru/AUhTnufT/NhL+yfyjIfs84pGjnU3o0Z4NH61hQlBsmCiQE+U
jxtm3kX9BPbO3V6T1RCgkZCSZJ+AISfyYI7r9/cDMYXwlXVzECvtXg5RkVvvFcis935chPZHgcF+
zhI6327zcvCR+ePStgOmjyyDCbcStofp9Qa5l1okp7d97RbIHenSxPdM58uop+UuzMZBNuR/yHdd
V3eiao0o+A0weEiEuxxJ2TOUt8yqeuWXu0NNEjldzZYfQRTvUyntrpPRlOKqq5JYBXvrAz6QL4Bh
tOua/qDyt0ndts+gHGLzwB8EZIqTelRW8MHfeDo2St4D8KoCIPXX+iLTOAohhozGgtW5yGkdJ62y
zHKMS+BkTgZw++bJPtQkELkIdVxFD3tRx8nWwMSJgN2JaIGfYbcT4DcwouXXwrIkMZG/ztp5S4qB
1cN92laG91iM1ONh4kGdwQ+PUihHV29PZcgkg3v4P/qpQQyLzjkhTIJriljpEZWMqeCTPZCwiz3Y
HxLm+KDd2BiBi1apBzLNcN0mRC4aU7rs8ioEdnFIs8PSsu4G7bBlZbU9zM/z92kttlzKIoitrVZu
Dcb1XYNovW9e/DX9WeQvt/tQQGaHyShC3x3yhoh+IrqS758oPA7I73aovpNTDaoEU89IpGngFoaa
vCrofcoY17pi4KLyalsLohorB/VacgG3VLODK9wtzG0EiZ+IukY49ImHXXTeBobc52FV1GkZAl+7
k0aXSPrjHfdJBm5Yq4mz4bNkTctuG4hQekn4pEtkS7FwGYIo61gcit2DCzlaEhpxfXX+uC/vf8uk
sw/NEjSk9qw5jCp+TMWaNrmcroTqWwRk3NTaKu2CFl1iYaUNcW1FLniCQxnR56Fv+1di1lKQN7/8
uEMCgzNUlGOIcNjAbeB/1MKlzpSDiS4w47wlaulP1ystfgRSDvE7ILvM+MHuzqW2aZLyUql/lae0
xCW146I+DOS5S587lbnu0Sbl3O6cw9aWE8m/uF7HW56xZRtTZI/oBGYTxv2TT2P6TfXOCEjwBRZ8
1q/pSShM6NPRMUr2IKLJ0R8LRnlbd2ZXnenQ+I1ZHZXD7xK+dEcrTmHBPhI3hpnYdjlYE39j/2TV
OdZABV22/pucjQKx85L7X3IltIXSVM731JVudKZortIihzHPF02lfbMaKpTzsI4NQKUk1pt4LAUR
ahPyvAWp2+16Je8Fmkwhr6y79+4T4YqHr2DXOp73HKcw4+F4RSk4eS7hy60QyhM/tB55JFa8e9BB
rb85hGtJZRHROwo7Vlrie9RdjmNgpNpIIKwajKThDwQymZNyZf4zLCki8JBnIn0WhtRMI97Nf4Co
Ii6/e6H0CLmWDU0OKboBllRmCKNP580Kt5kduzp5pGC35fAJWdYEgAiajM0Kgt022NBBGCKbppd5
i2yTyK3oj0JpGk3EycvsVRKAkakrWNwgdj4D5EyQd0j61/k+2qiQ5N/s7oF+vEXhC7XLWSHkmloc
9hEf3b+yT7qF4jqkbYn05AtKCx8XbANOsShfi3qgFLI3MjBXBHA6pFQhuU5nMMkg+VNZpRUqucGD
WwacyyKgUuzgtexWv4BKQwxGvw+M1ve5aH5V99qw6I8PJylFuurpH+7kknCY+Pt8wvjLuruwgyrj
70RPbm1Hq1tQkPtBF4XstHK9AtWvh0FygIQjNaaC8dWguH+D59ucsJGmq4YxhDW/7RjJOal0nGdo
NBFUZZuEgSu5sS78cO3ct0huMMVDNmJ+psFutmeHCJ9jBu3wLmLKCfHuTOkCGXfGTJbxH1H8R4/T
BCExzso3xXh6CHCJUxeC2/Ys2p64Pik2XSbZ1SN6RED8eviGTq/kFkUXL98EMVtiXqv5F++2pgJz
2tadJN7LAv52pr08FgE/Du57TnMYJYoXsl/iOMpmxNvfSlYCzgdUhzjtZAKtpPss/g110BMdaJgE
5FfdgFJx7p+RG+yTQ6/Z+LspwgpNg9u/nS1mJN0sKJq2098/B3QYqKHB/Mvb5gAEiLlay3hm+KMC
BWth3jac//shiDelyfylbjjy/QuU27aBizZoxOU7LKsBTT+pm/DoPzd1vDEeBR6q5l2ZluWh55G7
OlEvpO2j6N9fLdU7+Gzgcb3pxbvbVOf2m1ksE5mp3+s2EgcCyDyYNyjK9mZA5Q13NZb0/vzBz1pu
XKMs7+8jpN7hB3WRbybX7QbhAsTeC4Z40/zXr+f770tFT41UKKyLC8hMtxT2lLg21EhSONOhmX2n
Hq/1jjVGYlWnXhDwH/+adho1cPP99ldIu1FTQf67/yMWyk0ButGMKMWKdaYPGYSKkVuXQ6EPcMo5
hvoGzKjzkIzvZhnbQ5auj8Urzq+9OKXGe58NzO/aORyHL1plMTlbXM1NNyud0esYq22s7nVr0877
7Mn83LlFI+OkDn7Nf7o+BHdXCHtpQRan4L99F+X/sZ7gydZb5il3AXvvIlfCU9+mwfoAXHrK72Yb
0PLeFCoDJmc3dIv0fuQCLtHLgYtCsyPRbHgiTl+3bdHiqIAODMmBdCWJTkYWBFlqrMwyMlYSrSaC
YZUhgirvpmrJwuCYP1ajkC3jaIIQ12SCSEAFmkRr/uraR+AQRURkS7w1lnMrk8kaLuFi9CinlzV3
ZsEkmtsTTktqr2qDovXxT/vcmx8zOYOvf42Pc6BKfMmLB0CvyrLONqdCiYyjqkIXKbHk8Waa1Ac+
TDNlG0JO1crYo7Rss/IEG2tzETQ/MgtDqulfDgi/Ch74GFYjjRrnRKs5VweNObQBG5zBJSpNXcmO
FMmq6NfO6FdkXv81Fmcybx1vgBMeQaZrjtKzTFseuZmEvtZ8xZ2MQ8962Td9BoKc50EguWgM8y7V
q+YVN8g6q3vYZqnHOVFi36XksrYun3e7QTc3WrcSzTIuEw3IE2s/nSlV6PHC+NtWSawaW3wscyUP
mgds6xnHqFUcRD/m1M15K5nFOorTdZGLm9qZdbqMutWQcO8Xvqbq8Tb1eoVhvxcrLpRNk0504h6W
/YLv9wUmhRfk1r3MY71KEDSOd0n800Z6WCz1xv7YsyE7Iz++ThmfqhRawAYAlpIMUnoEwkq+2Zfs
Q8geWvt4QB0vXaIrZoa8dkmtPhup3QpupBPRkPOvuekLzYrTgedM0oKYFVi9BLoUeULUCqC+2YJW
5T4/odxV7pmcl36P46TBrgSML3cH1eamkDO4tWT/E7Gs/OfWqQ+9ZdpZqDrnv33Pea6lPQH8Zzxd
5mvzoggqTDhP6jYHA7FWuyvGH9lWrJYx2vEEOZuzgdOkjkIyv6r8Ag7/u9jzCCiwDsSkM6uBpEjm
R3QwxSiGJpC86vpVsWRgcsdsAbXHUT3482JjULtVjHBtwWRBfRWKTVjG727m+6FEKULBE2nhU9rW
zPqZWoWsIHNov1Ec0isv3/EW4NlRRp06mgCz8Jk7viNVZYbmK+zo0C0tP+hOvQondVOCMeAIR0u8
AWiTK+XFaPihESTbFH+5sul14HUcaLgO5b+Zu3bMt+Pg2vKcE4eA2WkxzzxPT/3+fviHK+nHxZkf
sc5f3GNHQ82XkKTmCg74q8WFypBWk0713+OtcJ80KMD0T85IJCwGcfJZkWD6J/dvyqRY4OYyLL7u
x70xzqDvplY1KNOa22CrRy601dbByi49rE48VQaEizzkW3z2MGmGtDIVLiLHLgU83MOkIxOcUb6z
auxAJZeoWoxro7RyKmtvxec4qd6/7Oz2uNYo9GkjPeZBVcGPT8W5xcaDqaMYMzQfI5pjo1EBCYby
RQFiid1wMyFv1Yi3UmxRrGoEljvuFQKoT49aRV6Vv7NnWEBkf5lxUQ2MQfbJ6iS0sBhglyNFVoRs
Gydj280SJk7lTy+obtSPgvkdHFiLcb0ntxqcMIOWG2IPViV3oVsitwLEukbvN5FbZkRB3gcU0zh7
wF9/yCFux7cW8agiRdAhBSG/i0Yms0Tm5uY5WqEART+4Sgtdqa6XSIMnU3rIYVRdgCFH3oDbnn1c
0KdgI7G0s8Z/xuEnMGbqaUajAyMFGYbutnHlZyxZoexgbCaHOk+cdxc4I3MfgGh3i5tqkEpiIexh
ypfFZIKS79G4wr+Z0182sF+Y+W8AkXi/YwnDo3aQPL8QC89h/dWEUqEtx67SomwkULGQht08pVko
p3Sv/vsq/0p5m6L9BhxjhzEOMpVJ0BfXu/ukAY4L+hzCwBB3g+BvCWfhyNOuQjj1vK0evoGu+ahR
GD3Ew9dy1g7mVvsjgjLUOTl22uwLunpTWuSN67vCEaKQkcuC0pYFt5A2jPS8MWpQ+WTeqP0YTBV7
RLi/kYo9SZp6DEJW4nXCST/dZyvPyz1/X54/W9Zn29XUI4npGm8ZODZSjP2Fh3cVHdjdsWYGbJz9
+ONOmWGtubz89W8vomo2U73k8SPdae+XKn154VsLUjHA+i5Z8w9z+zDNQBtGfzwFFvxLUvRoslDM
TW93O0d2nhCTnCGADKrMXoIwQ+EtMScn/XFKurLSVSDBawO/8vDs8Y7QoVnnJ2OAUzNsF7C1BfPN
boPwNwimWQ7jx8dIx3ODojCePZrQpUV8Mtlzzjxc1c2od/8X3jsL2Mvv9uGI1cm91TFKc9xTlHV/
KBAY2dwilKzsPFsCGkELQIvm7bV2PsHJ4t3o7xvUrxAF1ZTcHZFt3CjDbXzxFaqZvPqz3X7zI1Ze
UVRrn54R9mVNY/jiUXBY4PsVLZ6JQvdSRk4yeuCgtKxJhWVcOjcf5iM5OFFdeb+ey5CAGL07y5oW
G4seDSmRiHV2hbyzywVM128f09ZUVx8SY+xnjucCLS96XP7vqkFQDhaaiYdyIOEwoWKzGgbjjnZ0
68rrOCeYBSQJx/Vqdiz0sVL53GZ/D6CLh1skmwmxitnjb57Fhad8vWFV/aLK6Pn4zDW1aANGnOJc
WO8EdMzJtEQh9x7kUgkG1XnS5VzFFyWpBdvfO7CXIB8gnR5k2R2dxis6qqvvtiEwrJ6UzM5L7OED
7umrrG6GKpOHyw/3dpwzP4ERTQn6pVY92AiztMtT56smxpT0bEuZDcS3DRB9TNXjZPVVmYw9JTDo
29/XxLy6i6NiOYAF6gByYxVEL5HKItGngbnqjJIIa0yUpDzyZBEx/PnBJ3WNnjiQiTOX/8uwmGXy
OZP58eQ7/N6Xo1AaPU8rJSsu1865zUyC+gzU/CF9j4Cwr3hmU+goYG8NS7q2xRlIv9RPAv2hPmAV
A7boJBeArakERlOFl3KajrVBMIsHcGn1DKct0L/JcrrAKcETSmXta9afyoBC+91RXn+9V5nZacL5
ucoR/IFGTezQanxjY1EqSR6dyNXb7Kx2dr04RfryLO0gp6e/1b8R13cz/m+VTaSZMFFIT0lsQCl5
KXrQREkFMrfDhuMkU2KZ/hYdOXT5MlEw6QSRtzgNlymnQ4eQaTwfm/ZBENaITYwXQxnf3WY09agj
JloDkfR+2X5UxIIqezRamUfd/Nd6c3KxYivF9xH6eLak5Dkpz+vqedAiDBryD1X7usWP90Sassn/
EXpEKp3Qw418r2Sv/KiRPrmUvAgnyjcAHCno6z+tSvmJE6s9J3R8NObN307dl61J3SVJe5rpmxpf
wSSB/XnQvJIVcJplmXVHJ6tHwrRIKoi4cGo6112GCCJClB8QZUY4sJmAiBO9gR4D5Y+tVdFnjDBq
VKbEMhqBMvJ3aumcy774lJAtIXUuiwyfyh2uTIxFMADn0O6bGeRGULBr4XARtKYb+iY3phg/pVG8
vAs5Xp54y2vHhsl4V+v6nwqxsDn+Z4QqCY7cQcReH3tYi9BxhvUyok9hlDC5MwtqQhhgv3nf4lcv
zlCljavjMSslWVgYnkLVPC6TehhnAexic7qvJ9rral1XieLKA6eVnJPYxd/tR0pzgietNkK8H85t
e+RXcjtIwQoA259T0am5txwaNMJQN+419bTjCaLQwtZpc+S0s8bxpTFhv36rYxO2b9fpHEBU76SK
QPvm24JaiM7X/L3D6J8UEWNdXSvbqtg8Aa9Q7eNCTKOaOJLM2I6cQLOqAYWcgAZ4Ir3Sf2p9Hcnw
lhpSPVcLXTf937PKGn363c0lt/hKAVTxdmLta8w32wQvXP3Bbugw1M67aG3pScSWZ6b9I01nPi+E
/thFGKK7nREbeD7MJ3j5DDxqvhxKusimxiNlQk2ZHzILqdA+WihKuztCGKENHKkD/ymhlRmQEXZC
P7Dudj7gkxxFbQi6WDeIQ0tQSTAkHWGE+a0a9BNYj849OVUFLXToz7sUNKzRhdZy/t+QEsrLzV0w
kjVsAH91/YAUBXULg1WMYTdrQ1Mp5DeGwxhC7ziaNb5GNeTuNAUKTbahWMj48PT77b4lRFjg6w2v
QLrQOrm7K4QSaNu2DOu8/6xwBBAsQBHWepFRybnmAj5G3lm8VwChtfQAKj1MdLPX67Il6x09UP8N
0705FpJ0T5X7G2TCmQgT7KRbIqYvcIA7X8vi5iOVB9POGIotRrj8uSRr3gxQ5TyLaEiOxv4Ienyo
UVv9F7RinUbbmnSyATCRRX/44gUGFO1EwlqZ9nVCa+2/WtsGKLgIMy6GbyL78XlcrZOqSBWAvxZ5
VIlvbS3+CJ8LCGmGc+biFF8/q8FClYOBNp+1aWIsL4eT2t6/TBjK7FaPPkyGGZcG+lFj9m9fjiwy
0LpudJaXZHZaYyvQUTgvKvOlmpzvCAwqsZynpTibyeqDny0/o+5XAnpHX65iE44Hj8yPDyZKO9lI
ZxhL+iQPPx6ZJARmZqdfx+ekzadJOmQOwe3jsm53Iy/Cv3OxVHCAFGe52OuvUp8gzNzyIEec6Dob
qux2Lbs3HOMZXT5Bi2Pr2OsYXK1cseyeY9B32SrmVVyUVA2YfeQFJkuSos00ft8TeQwbfI6So7/a
tg+3ef+khOQt2Oz3V4kiHruD8++ayePF8f6AtxHq2IjzAPvSkf9OC6L2hO8xYH3MIkY97ww4OM3e
lyDsSogzE2Uo1ze6OQHob0O2pf0t1ZgOOED6R/dFx0kbC9I5PceagzMdrF/arsbgCVpyhinCSL/s
H5moKAvgmmkrC5/TWqqOJvYIkhZ055z3SLh9tKTvIn/E01edtAMWOxhcdNQE2/WWFLNPsYeQbzZK
vl/RvvrL0JGjhDR5hxf+FYC9vBhAEVDFmY552W6jn3tT8+vYUPSoa1gRZZ1+vBP7YAxEbGAvWF/a
70Xm6Al1yNms+w4Sxl8iRNXAFJ563m5cyWVmMcpf+OrgPkt+2cjrg1Ftt5aiv3Dioo3xmyLQdtyZ
JV1j+KXOtWNl1jRN8kNQKxFWi5kUg18SkTAgKV+wFwOg7ZPiqewcFPe0dO+jpHepwgZXjjIlPK1v
U5MQoHEQh1R+kMl2mY+5SDXasRxuWaurRm0F9MGCVl72pD2CIhtfG/8p2pCfBZoYvjV3YCn0jc+e
ujS4P2iiTa9QtKNq4bjBFJh92gy45nmLRWYeO/JS9fmOkny+sF2qIOesGphkVwZdLgfPQRQ4claq
tjQZhLkzk5cRGUOKjvPiXcEy+vqCKzFUrkWZ0oIRaDIM/XsFnHEKSsfI8IiFHiqgrKvgP0BTMmL0
TJOoqQbac31Uly5yl1yONTrBvVIXo2OfV1KjbCiOYyNeIpruu+Jc0P3hW1Gq5xotMlohSedvV8L0
ceC5Q+mk/Vht+7/3VpgnA5IYrQPxirlJkyGxim8A14kxOaP126G2WeitWQRU3PSK2omjzvNlyhZm
n57u9v2cVusUm33Ol/xFEQl9zAB5qzOSZkerQKHg+eDi8PFMIkSjbQg3qAqNvxdV/hn3uFfIiJWf
EcoYn5O29Gg6LkZ5laIKik58gsqOmaWpr1cSuQHe+Hb+fBQRtMUlgPOyPS3v24YeLzcuqzAh0Ina
Ag0kL0Q/pg1orJYryJc23VxwLqlLaRMs5x6h4G340m9ScrtAmHqj/PPW7EpBUIPjq8x5ui3Y4LE8
vbdOV5dMXe7ZFF9ln978AdN/XskxWapn1nvmEqOHLr90sH2kRcAE3HzGkfAnixuDd55B7c6LxO6V
2u7KCTFXS0qWZ/ju5cvcwYdk0GHofVoXAda9RimzCjRfY4gy/cIQnHALalhQixKqitb70kgn2qmq
OUQx/tZIwn7t6+7pLIfvKvP+RIAD4CSrbsnH0M/Ib+X5jjFz1/OqblBtHmEbWMNHJ0qNpR9pHXAd
6nbHOl1lqozbgWTdu9apAAlS0mRY4eNHrdMOBGDTtmDxXJ7WEVSS8eLGMv3iawDFvITLy07DX4Vo
Hzj2vIyA05jJN6+6xkKoK5Nu51a0XEAMwYRYnXTGmGMj8dDf+InvOe9dcbHbcx+9KCiDn9VT6yF+
y5atK2imBFGHUqRdbvu/5TW0Pdm1DFIp18lmVhmUtci6vyNc0gcfXt4fBDkKbSw96r4lvwLW5gxd
7H9VGMKwvtsRi8zOIUHo9oHTYsGZ69I/jpED24yeuoiY9/EE77uiG2D0gBni2+L03847u3ipVID0
vn67exDoB2YjtveB/NQFrWAefMPVERc+x4OLgNJYgcyR5p8KBpurs8b7amcHaqhP6/qrrNHVEB+X
BtOAgTKGGbu94W6t+ORLbXHqN78avhV0kc10SJwxnC5pO1gK2Zbzb/+BrLdPHbui/yjbQ1OZMzQ7
MBVLMpFdWD6FD/lD7NgWA9yHawgNUHM95kSk/auoiQU023GMUUP5cRvZbmPXq3NP8dWJ+KVQskte
AISPhdGhgQKa5DtS3iB5lRLic08GZcjC361DlUxStC2SoZQnvrsXLIT5Cvqle8+4f9Jx9MeW3xQM
erN/qJWt35Rj0CWeRDK1lzRYEj+Mr2e4HXnuyc9D4g+2tFy0DjZ7MiUz5iIHmGnYVStwtKzPQ3Vr
2IaN2vfh6oaFJYT1t8ddoOmrCOKls9fau/pNYLTD8PBlvHrafDwrEo2yooCxfFzRTooNmxzLv+1B
+K7T/9PTxmRhLn+q3rRSTuRzdjCtoSFksV/TCHjLUPMeb1OzgW11j2dF9sHqnWovkHNKYty8e7YN
hpkvj9qDK24tUYwRe9Vbdchuh0FWYmIthhD5WAZcR2f9Ybb6VjVwUkm6uzzAsVf8WpeDOvZeA9A+
Fi5koCGEVJJi/zM5Rb9ryRNzYBCNMKjvQ+2T3Im79DGk+B81KXFCH/1G+bjMJNLtiaRozGm3zy4r
bqjir53c1rMh0OXt/7xp9kdn1rYN5xWR0PA6woilus6xQ8M+QZEYrslydf5cpPNh9RXJZ1XuwJG8
Af6QFP3ytW9xcdqRLyM5B2IH9sMEuZWxUEXizz4l5OAwt3a8SNw1iCoD08WUiRGxxKCsDjE/JB56
Botdcgs6DT82aL14R/mnJ1hfwgOJXmUcj+VvWubjB1V6zhiO9HE2w1rDuR2w4V0IZxZGoSthmITM
TP05Y6eMqB8aoxcfjBXT9/dt+rcHtnN0IJSCWyN526Ziw5YC17KhOrnTIeOwLBX4j6JHI+2o3JhV
Vtl7M9Cgt0zmmIsSVQ4A0TKQdf4BmW3FKtCrvKgfH+a3Dn9JIbuscCtuAB7q7rFwl56oan/Ca0Hs
Rs3rn2YbB8YW48qqcPqxV7I1KJCsj3O/W8SZJQMSsAkvouZ2cl+YF3wkqQDiFPNO+Tayk/zfWZZB
cF1FvOiu8Y2siNsUOCh5roHC/cBEt5lCz4kpezOaoGSrcHAlu0CsvzLarAKREZpSCYMXcLVSE8EZ
TnHrcWVFJ3a+Ptu6Un8EQfH4OUnNZwYIvZCw7Po1DXs/rahHYtrYymN44sEO6LEb18wah/jcd1af
L+k+aR65/dfh0rtKYbkK+iVFyTqqEOvKpTdwshyNdq7fDT39ytNJXfZ+yqAXV40uJ8Vi9yWjgL/Q
n+jC16nSUm7ernkngfzvD1rDbcNRNjlevRASzExx6PGga4XdMXBm+iTqk12MxMW2MSpMLAXB+Uif
pqNayKPw/ycB4e3K88CN9xdeE8xVw49rzRNfHufl2P78wqhhhcQ7F9LDt/6vIpjaJzMJxWRswjk2
4GZevGZMuVCz/5wGyV9CGmsqzG/dLppKteTm1KUVoSid3FumBdH8oH5Ip0aGgFA1EFISNqv1vyOf
1saKdDbXJfAZO2weQ4nsqEK88J28YT9pXFIyWr0rEm3S1WXif6FdSsfO5LlhiTZYKulJ7coo3LMF
1DXLY6R73KtLfY3yniGmpDdR9NKFM+DaSq/7EEjARxtAlcnEUn2TLplT7rchTaEh/X/yFH7auyWl
6WpiXq+46scvWx4uIba9v3CneyAxyqXXH5IAEwKMiRdzkvB1K4WT2ZeySmSY/4h7jGj+tJRReH9A
3aX5wrK+7muz4b8rDDI6r8vL6LqnQDUZNOfdzvCwY9jB1XRWMJHiBkiqeh4Cre/KeIc12VPp3jRk
4CCmyR6X570q5As9N0iNBVjC4WKTyT5zzqJhB4rl1N6VLKV/ZZ5boJy/ruspOQ2kmlvs7/SZxzmE
0G8nZ8uTap8sRaehM3DO0MnJhw+w+A/txAEEx6dtnhuSVOtjuT3hYdno4DDlta5ayuT1+EFSDs2+
3qnvQ8jOURoyj4cgpPaa4TrxFM8dMF0J0t+pi6BM0/RvJJopL3fPHTUQvoNA7NiQ95uhWAeH8P3n
go12SOB6GTkOuLwyiQAGe28p8cEtuhP1z8oOCvUhiOUg9Sb8eFesF2no/Kmh5YNTvNHJcFXTwRjw
tmGDD4u05AalakDaoRlExEKv5/13snRLAVwuWrvGQUbOS7qg035d/OjJQ1gHwTyWLUqLE2TrGnk1
aCIZzNzKYyWtl4cGtQF1VwF3b2kvjLLXD3YO5UyEsjA4nGNn2ebTDZPcZF08sQcwDZyjr3uwFpft
aFZrn/xG6WCPMScxnVldZBrgV3AQXgcC6n2QRMeQ8s1POB1PDQ0OSGj+yTsEcoKQhuDB0t+Y/mGV
+8aJAwwM3cGzeKytcJugw5v3AoKzJx88SKFDlZcZarBlEMCgs/1iycsg8xp5d5JUT3fI+t8FlRN0
DyTty7fSRbGvL4fvojBhjnE63RVlOZHZNII2VOldAe79VqOaIiYHEOPGyswd3k6ervoDERv99P6H
kUjlGXS/nZet5I+XAWhyxfeAzx7Uy8oUunmLnOnmDS3rib1td6ZoxWvOKFaj1xhg+gsZ5Jg5yabE
mTSGix2NtJcdO2oNqYlfXw71Bq0CR/Av/e+qhRIbgOUUmSfRLKcxLJ2bJMucT13+Ec23pSldfFao
08KOfkBdmAqWul29ORmN24U/lJvh+0rv5G74aGCfY/hx5SZJ+qKeMCCejFPGVJn51qkdH3WIwgZ9
2IUWWl6gJjYTkG9hGHs+bP9DhlhEtoHrUE7dzlYdDvzsfkZm84z1NCqe3J30O6W8Yzr/GUThLK79
v4OAI6NWnK1fN2daKWyiLpXc0oN+aK/O/6N5xOoYM/KGubjUyalaR1XGbM7DFBc9/HC8FlVA/PXZ
Uu3ff5EGqX9BXOaJP2y2G7spT3/MJG777ZdMh0PJY+D4BgmpJAznEj6ha7rP1YgXAO20uiKXIB3n
y6KMWer4XwZbB14+oXP/qPDt0s3EOg5elCncPerQaEthxzdiV84y1T2/r7xVW1EzwsHi0wdMIzxE
/kNhlI2caYNDq9/JmoTpLajen3h4XgeY2H4kIhL/umZW1FnhAhKnT7SNkYkZHM0s9s5P9p6anks9
ZnQVsscsVAmRNLguQMdeeGkdzhoAiHJ8G9rX5J5xSRPR3AnplRW/edq2C7stpCu5V9w+qXlTTtuR
+pi34PbgMRRWRIM7dH1WEiCIeC7K5kkt4M690VWGfx7Yh7fYCtVojoyA2DlHwjF9b/It9ggX5HPv
zgGr0VOh0ERcdUA7lH/NDhXBmqmpaTs8NQXGyN83dVhy+5RTYr8aI3jpwPSoyxEKelL2Cj0QqNbw
424Ru99WeW/zbukRvLiVyq6vjXc1f2Y/JhvDyb6VKE9zUjMEF5/i/05EpUtjFvnnAJhAK7hqIO0i
dXvdoMnOxGbw4ML9seaVvKwRQJrhoh28UeIRjkCceQCFbPmO5gFeT7D3CqMaEaLuixbg8bTwEIxh
JdzOmQRh7TnsEFZ4lirsBx5ly76o5ABZm8kXCEfkX1kosFRVDvsApjzGMv691QZBqTMNrKCX4bPV
XI6Dc9IRpz2lTJPY6YK+u3h51hxYHaXU2g1f/RGVOFtCeKYDHvoTceRH4OmUyKi4inF36KjjZyJk
6H5fqDI83YgAwWBmDz4iiaJ8vowiY3wsd+7NCN6l770zmtxLk1KWpYDlpMN4nxA0idel6I8jlpfU
9wWbeIFCNX+887quB7IaHtJ63suwMdjMMSHrg0iGHUXoAbih7D21dJhTt887xs0KmO3A+rWn85Md
Mf8bzK/Np6wQQliOnBm4+ZB4ckuI2hfouj3GZl3xrZCiJGLRpAgOxgizT5A4E6sCa8Cwen8/cBd+
rNPDg5ZR3VHP88meG396JI55Jrtf4XynfTKQ9UpQoI8/Mp0QMrkHRxpZc0kYg6G2dISQOlazKORC
7pJBqs2XtzfzPvyEiFWoJSjajBvJ2MTDg5BJaHCvKrxeOZtu3RYHerC3mgwtjjRm05F9TwNjBk1X
oy+9iaPbM8kZvlZEkN9+f3qbIGiZdNR3X34Y5SdaKugBNrMhOV3KbD+UCxc6/XzQn/QShw+Z5LXs
9J4GML8iy0qbNQ0gMca6nFUr7V0gpC2D8fg1BQU3whK0RxgPCZaeV6y60z62M4ZhyMAP5UafA17u
lIc+9v/s1H7twYcxn6kywQ/TxdJ0/OspeFwOqglCRyja0EODs9R8Abgu5iI8ZKRguF3Ri6pSoDL2
DRdfH5tLEPhnIPUBVvJMsGNAs8yHvzSUicNQTM08+RQtCTnqbvF8+1N2YAlYlpp35FOcA3o5ZQ6D
AksZtPaOPE5m3Ga8KIESv434YgpmEE2uHHCRvmOT7Oe27GJTQkoBmQIeDtOsoHaqCI8P+dKVOepv
gwJaOTk54loFDE3/87sfzZzsuHVh7dmZJKtGo9TkBTxrfMh2olnjiVf8j+Jb36TFm2PHlqOAhgsH
WZ9bPotJNDPMbNodoto+i3HA3wXop43EQM0Y/Bp4zbXCE4H42/mHCbKnI/4OEZkd9G1+HmSRE3jR
DcU9bcL5jbuUzZDP134yevR1SObBx4BqK+CQ4lFMC5wgqmfM+JvnS8EMFgb1ojovs65SuPwX9GLA
Q/vmn31P5KsFPNwWSVVHb7UEk4hxd37zOLdb/Mq6gw30FFC0YmgSGRHWmJIXlETli3n5xiNz/wUD
2g0i8QPAbOHCBWSr4/ClQgZq8TqcGtbf/Hc4J0LhiuJOs5E5qmDKDOViVS8R8K8TpWDKGjqZvbje
n5LF4u7ISZQMWbPmLpoulxhkrE4KUZyv1En5SW8p7/xW9cEQ/Q81MOT2QK7Rt8LZC1NAr724RLZk
/qRooPVopMWjFD++geAsGpz8tu6omcHVIe70FhE+VJJIEZNirbzFXK7N16ZFiV5+I4qLYdrDnBfJ
PxcTstF5DJwTx1MwZglUGeCZQmTAvEnn1Sk8r9j7oKA1GnBtBriQGXIn11fwDD/eE9TDlLQ/qNO8
00MfOt6kauqCoeyKMFhPmt6m2IbEy8Vxf044elAXqN14muhxTFgWYhNqEoEIiidLY1Ow6vl3L5S3
LOLeJ3e0BLRm1JQWgHubOSN5cOThKc0csH89jKKTQ7frcVlZ6/wovKwx31vnqmpbnlJfn8E3TW/j
M4D03RoojRvSDpWSUaSEfOrbdrUXg3d+A68WAplW0CX2aPk+tNmzMIKE4Onun2Vyu88sT2QdRBUZ
ZAM2gG21NTGoku2tNDOBrkEHkB0gOrMPIatjGWgJPuPxV+rQ7ZnrcjDITbe+voWPsU8sy+cEdJ9p
gaszmFbFVuSAd47p7GwCC/unfmfK1zo6i1NI9vjugyGYo9C4PK0SUfti1hilL1osOaGgZWudxpc3
CeZFKA8Vf86N3UI1PEv2ldl79bm3WLBr/aQIgzcqqpBS2tsvrXCwUrEeSXfpGsPLkeMZMmtgkYax
AZqWaeMKgfx8rxfFAHmEsGJuVpaFsq8hv+vP3Pfehi8Iavti6V7KPt6H13FUtDGkF7AzoK1z0z/1
lEhW0UOeGwvQyMtXdHUu/Og3NCA8YXFRlx2LqKQCdZhxJ/1nlMY6ZUNuS5hhP2wJ0uQR0QqOqJEE
yoNEGw15Itlxfmw2ErOkqc5jDIezZG/xyA/QkLBnFdSHWqJQS9Bgl/kykAZqOvMk/aUFdpFgvNWl
1dOcB26A49uxsFo0ofCUm5V9xN2SDy99Fi+fV9SOGvKbfaoMJEoqpvg/aJbSj93hxAgFL8xdo1Wb
a8jjDrh1wuCbWXbc2dYayjKNhs8ccn1C8mCoBwGXMJgLnlNrqiTe9gAO0AUIcrT0hAtLgcXe4u/F
+/xIDVM/bPcAMl4oKu4mIjHEKbIblSnXFXkHS+NN9+4EqRuODZdibmsgv54oISLyrB4D9Z024kuE
Y+uMTJVS/IbFuWfU6N0cM0KdJgndb7oYegO95+speslbWo6SQFXmphgxHs+ZMJsJNrMmqozCNGBg
bqZegYtd+rOLss50zK01AIz0T8/Gx+8pVti+CwPlvmVX+KKsz3Ld6P8ebtLOAfEhGXEs0S5XqRt7
wB8pyQXXmBM3dUMno7WmTgWfHpNuzeI3Z6RqhE966G7iawNMTEbLzm5evcArK6V9lO8LfaFdTFc6
al67RbmxzO7MBLpYEunuFQt6E+HpxfNQFp4wCI0YRyE3GF9HeIM9ROr/6pUZYDwdvFARE/cpFpB5
fmiZnhjjbXwNskWX2/XU0l3Apw7V5ujgJoAjft8C0cdP0iSN4QAqb/AMOUJQHlYQbzlYudHyOgjr
t6genXa6zvuuPfveJHXtaAI0qT0qAEbuin7ifjXeMUSLIzFPeYbovBf/f7KExCDQvIwjmKpVquZr
rIAGJxCxNHq18s+tx2N96HxSvTOfjR/k1FA6dbRkn1qzO40xYpUnYb6C7ez77BQdbxBDyS0s9GPO
oDCl3WGTJbrnVNWepRWuxRK3J/yHFA8yNCr0e0no5VZq9uLObczw/JrgdQ9YK5RbytAwbRApLGZQ
TWv4EPVi6yqnugdD0wiefjUUZxo+RyTNkRDaYJLEyaVF8tXvSipxrFqjJtnWCcsmlggB/Lq9njYL
rHLqigairgVlPCDylAXaPr8xDAbKLXrgIA5c/oiprW5Wnr8SU5UWx7BBWuVh84/m3PtV/n7o/Teg
PJ3tU/zcJSUqOsqLA0Uo62ZMPOq3jPX73eY7UdBknoQhLM12r3A3+m02sLtccF755mTefwfBA24w
439Bif1iwJknoArjrZfDOghbGET+0XgjVfpic3A902DIsMTbNCBuSYXa208QelVKFAw/VhgPCtw1
E+IB+twHLHkNN0/UOxmP4IoHAmbdjhotZvwBJf3ejI7ZhNRzjFXEQ78VJGkuxWung4lKN+a7cY21
NttkqKqh1aNTY5vcDcMvU4dGdB2CHwH3fYF1/nKqYub70IWmD9VbeAxsfTDBpUOt3s0nGSum+5r/
cF6Oy9fgelPQBZYINjMHhvXEdWpglTTTb4NzOvGAqAy/k/hKRqC82UXHTSIDXUXo86xruzenCTqf
qD2S6NQO8uC1NgQQo2a4+1Z7S7g41mq89DcbeD55xJGZT2vrvEbUdcLCsUtEg0IbAhCzvPKMddpT
ZBkUgcqJVrF46inmzau0+STr/XHxz519/xWZdKMHHoncNNqmOC+oZViRM8p4YqyztDDM4dgzihVK
BWKLkNdmGrEqZbsdM1a+cR40iXZadPK7Ps+L2Xq9SsEQaVl8Ijpr59iHf7JQQRbXGIIXJiB6eEgT
DIM9Z0vwJJBg0OG5NOA4EdGNsR2MDkRGkVx+rMZs5tkgejVbyw99IhvQLO2JHh0Nn5fKlMHMT7zz
26AFdZTMf8NS7SoTkmFlce/4DvtyO8rT2e8JaanfNdsYQbGM9qndvIpw+porOzE6ZbK9GNo71/8w
lRBhcaFBoKgoGbHPOoYOZ7R5lozZZRCnXpj8aSH6lboFK1s1dvrThAgGToGWimquN1e9pTAo0Y3O
jpnibFIFw31bBrZ4vn2BUKBva6Zmn9k4Yi55/209VnpF/NmR8Jssj00j+yD8BJbi6woAlt8YkdY1
MZswL472x7ZXLkv/tHZGL2kWymutRAalpT73OUz3BnaHGxeuS+kC8DhikghxfWaPHQFMLOP0+5c3
/wxRlnTmRZpzRiGdgcLSow8vy0yl9wutHjOSZDotJhalKlapNePBStIH9ovm2fSIJl30eRDZs5I7
5EtsTK1IAZqMAJeYD9gd7Of+mJMuxGXUOWuguGG5rxSOBwkrPljpYwLe7tmburt7oiuI1adL4cjP
5+pJr2ts8VqH37+lQwUw739j+Zm9Aa3eHDX4hKS2LgEjZtqNigQ+T+KhD94MPWqFffx3gbHvs38z
Y+OZm1qju8Sqh2KBlhHD6Q9gso4EXmqtvPXwmNMisIN1EJMSkMh4l4TVCrQP5Rp41FnnQtgAbIUT
k368jltTHEQY0IhzMgw1Bm/NpgRPn3AfXGZW3HONaQ96N1DXj+db0U82Ty3xADPWi+gCU9gQ01fF
xhfPUHJ8k4Kwl0ehr7/RWbeh0pYM/fOU3GXraiYRp+HTzpx1yNYu2N2wEQv0i5tz+jlzX/zAVErB
IFHAP+73r0l5GQ5Z00QG9CBwzl02FRBlPvzKvgTVRL6ucBKJr8JbuUYmABvAkoSz5XFBLi0k0xvZ
q4S67VozQKlqBLAFECvNzvxVGiFEEIQE2s9okCdE6+o2rJy0mrO9LUQAioGLIEHG2VyU5NFT994w
J+m1/Pq5kBRBySb6+QOJe72qRBM5IruD1PETPYambfiOTBM24uGY0iQowmrZpkw/SFykVncoFxZZ
C7nK40rY0rSUuhthLsOqONdIv3lywqiafK/8zYWmyc/Zjrd9bG6CVGyyv4PZaQ+dRFFex93UdWln
vByOmlFFZyHeMjgp2tJcv8gKHTd3zTq1sai8PzKfpEwCFomrVOuEfRkTjH6lusp+nbSp2kBSr75D
kMbmG3K6Vz/gZCVKEVMzFDATHaHpMvNiCfBgEWOcywP/HENG+eWYOwSugmE18ROZMuQ/fUM8RonQ
GnWBH/DmPtutroQ3Lc27GjGAyzlC2shmh42H33qo+zbcuSOeIJGF9or4NZ26W1R8V7HBCICP6a0f
7rmxU/rGSeKvyVfDtUoIX7RQ81sL93GZX4PEgQlk+hMD34k6yuxjKKe2Un7O68Lv91rtsWPSvdF7
MyNS1ayZNF9yjFr3nCQtLR68awoRG79lB7fzxJUjqMIhiviV+6aA3RyOfCa6sfAIFxt+ONvuBXxP
KgwEJjBcVrhN715nuWDR24RtvBH5CiZ3h8Be/HJqOGLQaRQqxxJZOxRmzNElZ9eI79vG8g8qKKL6
t3IwsgCk281P1cDBX+KEUrRVy1+fHDv1VhXurNiEOBCmHnVMTQH6NiJgiFlY4D1V4yqHncpPQDrg
pV6ZuIcZ+TYDGbvl8xwejPcWn/qLON7oqijK9gGGesUy2M7durzTvtKD/EUQNpjpkVyC87pmaTkp
HIJzq6lZJLeNmkInWMY6QYjRtR91dghck1601OPMF4gDJP3UE7Rla6ubwlq4HvSE0qIS7FdaLAiA
VwQZxa3g7SYJHx8iAjUDDzaCfohtluyFXMYEHK4+chNqLKpcgWPtKsryM/2Rii7ZUyTyEBca2o1a
4iOZqxRDP/A4cmTtjhbViedWqPJMk/c5eK8clEL6bLNVwkoq2dwY0Kc7drRCwDx8dOiHeFAmZQMw
6cyF1E+r1x5y2XjeatFNo4bXr/j89DeRvYuGuVFRu//GDHf2t8h1eS6+osHdcvriFE8WfToXRKjQ
poeeh5rXQab3hUXH0M/spvM109nMLBawx7eSE9RlXZDOLKXBwyW3TjcOp82giLZFDG/gnE+98pGT
uXav7d2dA9ltd6zZH5pPX7ftgmECb48pWP+iGyOmbvL1dP3FkFYaQD0XtnDA5sleL+UqNMvLJFdQ
WPaG5dQQ4Pq1Cz12sYs6H59X9cCRb2EhZfijbK80tPsxjm1B1MPRUaQ6KD1hgWUufSIAM6A+fzMl
ilVUDUFqzAnIRX4Ik9tx8F3JLVqWrprMPg3Uoqby1B/aytolusQCmJloRNtHZyzXotc/VSYu87iq
Vcfk/9FY2dbatNJgMm0DJKwFzeawvcanNDy1Qy4VwSChJ5MpEQZGhcCRPbgJg31rV1Kos4FOTbsR
1ChjMc5Yn7vMFweh/H9TbIXSYng/0tsf2TN3N68n5Ljdp7tv29oSuHqgrbbxChjh9p4hGz/rKg+v
5c74vZPqI+bkJHtrhFwI+f0CE1qUOhARbgJdfRHn/wZtwUSAu8vFjy/z1kaXoGZhTpVvWcum+Wh3
teYmSv1jst/H/W3W72Z5OyOHv9MFpevw0XNuXT/4n1wo/l6GdfTuWyciOhfwjPIlReXwQj18cDjO
bAamUYmMGauEbyYXnC0iqnL4R6s7Yb/xDSIQ+GIu0OE06kY06I2XvrWrgSuceSK0NsoYuqAdgOIZ
3Z0Br3hNzIYaaT72RQCGwOuQ7zVEk3CyZR1jWzBYVZ6jJL8FCwIyUCCK7/rx+apBPzGX4vQfQzT7
VaKh1A9qPVoUPMO2HK7dBAYmsdjyNT3YhRd52vDlY7XZmvU6O1Gj5SUfm/DuaQiOSrO8m6q+5VJi
s5YiCZ3LhtlyH5cpiaF5lBMIKZhx3AqbNWjGlw5qJIgK0EKMzrYNvnpb0BxGpQ9oAd+5DR1oPZlR
Z9QKaBeHDwLWxQygoaAq+lLS3KqOlMVaulMYdE+SIsfm06sjKg+qSijwwIhuI3DnBwKKylamJmX6
A2lUzfdNnnoUvI1fuk8Gn0IPMjh1iSztzd2Q17LjG5gZcY9Gw6CTMwTieVd7S0vs8QY2qnVeBMfg
iHB3gIjQnaJhnVc0WJ+2eXfdnvIOohzWBtpHBLS7YaXza28lw6Vidpm0YU1YnTikO5P64u8sdabG
KvWUiwGAuqie/D1rXxp5mn/48YF5yRcjyCwRia9h6p8VPoAh2q7t4dWwk6zWVFDCx0WwFg0OMsk6
4ctjAlfCXnz59b1Bu4NAVp5pyOsz5wQTdvr1W4u1XKI6SrZVCXllMGs8tNcA59N+gbf+xgCAJiVU
Zbq+riY5rLBaxIz7OCDWiIHKCdZ2hNxjxzg2bun8IWYvK8QsCFzAdoaKkTxznPYSNT/dO0qUNpfv
rQbDc4YrfKN8an0IJNUHqqNNgBBy/nZTBjvEgUBWKoRIa8WlwWenCvmE3xlENyrhnQOwf0zLwu62
6/uJAgh414CzxGjBN2iKl2ixi+jJQqVrTf2LAo/yrD19Rs91WTEW7MBZ4q6uIAOT8zf6mzQi2MCZ
g3M3S9MkHHo3PBFwk+ejq8x7a1RIslOjEuBANDX+DxXaO0875lq1oGT1gWJ87rHp9xg9+PkoyvZY
l7Ofyr8miaAiEwsLLVvNAOHOAu+WK9JQ8TzpK5rjXfcTn1fS36ROyGEI4Nju6FP+/ZzaRHe8JSt5
TJxpoPPqLWdOI9qFA3clr/3rLwZZa2gBUMLrWTFx+wrPcmupIqoAHMGrem6AUxumdp99BENZt4zc
jjmjWEDnD+cfvSA0edH2r7xlw2nelU4IZz/DjPnPDlh649H5Q59WiQXcB2f8VCS+L301+2iyDL+f
v/4zyOAXuT+I3f0oXNNrJ4G8YsGVmvT1lBOgHsn2heIIIduQ5/NmnPFQBJh6m6uChB07EvajE0rw
bAg0hRo/GzAM2t+jWBv1Isg7eUDEI0taOxHtSzZeTAPszIbO/YCBEMHU9+RrmS7O6zYYDBz+/laf
XuBZtVZ/Z9Md86vT+a3WzitH1zWMTPGf7hA701w/bL3CkeI7oRygSE9uT6j6Wq6NOT99H5l6rBCs
GJFazLPKU+3ZNm5wUOk+L7NCXY3rj+oe+/+ZzSSex5LnibzjqM9PI7sGTtGpFMGC0eMO7FepWgY8
Po6q1hJFE67rPk4vMNxO3rskABvz/66hImhr+2gAkyilZ5w/BUwaHKOPAzZDl+UNj1KoRUQ8oI1t
ppKEpWyFhyIbcnkDekgtFWkB2+4s3oJ7bOvjc/bszmY/66Q/g+va8DPJ+2nd6LdVAXLwwMwy7axF
khs8ui53Po57frDbACuYffxeL3/uaJbYg0Lf6BCOOVWXfJi3PT87kMjoAQpIWHqD+vX0gGRSh27t
BHf72s2NEXZ7MNryAXO1+iBsDfG3QgBbzRLoMOiVPpa1wFq3Zgocls0cZeZXvCdWAAdaBwqm+6Tl
eImdwhQF8lmqXrV6lXdy0wE7sgNDtIefn2CRi3K/hAvE/uLZiAT9oA26xVjxVXvSltPbK/eNgkYI
jirn42QHBVpAl+HadOONHIfd3YMUhIcgaWP7tFQrzqcQLr2WSwq3QDVNdz2EDaoT8NcbY21ruz0g
o+B78XJ1Y540oFbV6ljIuE1fxfKQOu2erOe7jWhdGHOsfVzr90B4WaAnHlNGZheLQiD4vKEb1gBL
Tj5c/qbiTEahxC6rRye3o4dzLyECazUDuGX8qnItPGBFGgUslYrfEObf6sOVirUN0wski6h1kJOD
Z8UbXQyfutoEVAA35i5GopNsNS7pKFgyB5iIQIr47V1dbgMOcTAE+2RjEzdnwUo9YxQfUdyzc6R9
/g0SCugcjFJizyTA0DAQnFaBBzK1AiJZItxETjWQhknD3KZEfekuoAghObezs5eDPQ+Lf/BElq4Q
xMxfEbpiU5zsCIWxKor0Ga1uwTv5UFapRVW3Ejj3qH+k/Mx9HYQVUvAzoadyiHcLI4jNbXoRnJ0u
gARP05ZjVxGBrxztOU5ORW4IBXm7//VE5f7qMD78YgsxmWMdfzsyMjSelkCmaemS34baKlVdPQct
432YWE2KqbfW4OIaix/OORmAj1HLAO2MkNBsjGp6b+G9KBONHfWQjks+e++ycYldqY9xeUDkCfmS
QtmbhtO5kfN6eJzwymUkfYdz0qsesDMYOuiTEf9/3R/1kenWJK9bGl7aPiFbcaND9AV0mbcSEfKb
fVb82uLlD4L9H/zeE4crftU14H7r/PsANIsu8I4TARv26FzK4O4jaaU+SgCfxqF3+sGtMci70h/0
uAuSNDgI8DJQlQMYpfxp5Wu/8yxCxyn32pnGyLLewdEiEaFFSMd4UVWPcNoM7f8w+Ai3/ko8V0H0
svO3G5IKoZwt4T05RJRsW2IsDa1/yCVTdIZrRaNTBTk/LHnU4OdWivmtcG1yg1DDy5EVTp4RdYmg
68wmBohucZ4rfu0D7l/fRb1plLPt07+HJJj77803Ma0vm76pKItwnOebnYMvN9eMuqJKXf3369AH
LZwGPOJWbSgQnd0+Iyzs5kk9TqpYYbIxQvc36bY0KWqND1XnJADWWArAigv4EGhE+u3dVqwXJEPq
GBBvbpkNgGynkKb20B3XBg6+zeu7DWfNOgWJnORY+3fmlQ7Gf7ZigI+sXiIQJk4AC14PVRry8KFo
nHSqaA5u6NyqdZKTwVM7ktKGMnlU8JNWa8xFomNoEUUIvMb6+9cQ4i0I7MnzOg/xVQBKiHSBlCFx
OcIs3Wff2jigrNiTqk6mohSKjKswBW0glqIpJww6Qaw8OuUYeofmJBDOt9ZtebAsA9P37iZg6nNZ
8+Ru7dgifEcYLQfzhnv0+qGkpo/QvA/2GHaCgoe6eoXPjMSv7ttanAfon+tX8Bo+Eh3egWsf7PAs
nS4U4oLaQA+HptSmHGX6LITQrjdp/MvhFzYUbZpaOjo7scP3BGM9dovvWDRYnTca2ViWpr5LWFFB
heeFXbFJsS22D++jUEWiekpOwTxuxni9PT74qeIXRIDHLI6QWRQzU9PVxDO4kCzKE0V9fDX+5TFG
tD6FgH0gagv8o6mZHV6PReayoFdjC1+KS2CG4lqurqzW9sbjH5R3iXMQOmo4Xk8OgbmEkZtf9diK
jOBW15vF4PHTn/xuvTAzAK/Rm+bM87Zrau5Ax//NeSUI9RehEiPRRX91n4IzvqJJkFLxCMa23bX5
gSuigTuVO+P241SvrAH0vhQ1zAG7l+G1cMBwYz5Mp7RRLMnxULyoq4XNkY9Fo37fhVo/AsF8uP/M
sd9oOG5p6tDbW1Dk6Tj+6tYZwlrm8GrHApLhC+BOaFf0fgkZybUzrMjSFXUu6Qvv9KP9XGgWd4QP
Od+mAwCcKF9SNchroyhvHWvicNVu4TIp8Vf0ASf1fSlEv2lPjFySn+Imlr/+oQ7CH5O+k0GYJkHW
pPtNGlac6J4Cf420Lpu8kCzqcf+JogCFCDtkGilSK/DxCL+FsHuu1hgkri/8yitY4ebDnQKyPwO1
+jipfO3UI9Cc18Dmi3WKa++ob7wV0fAEG4JzqrJ8H8GcvExebRun+BHFLXzCfZsD6UE3/4VsrXp0
WzqcQvxRgO78tnP3/fJNLoWyhnQ4e5csgnhz2OvlGNOus0/ZLh3WiJT/Vwcz4ZlKd0dY1f1t1WkG
4mD9dRPfYXfmCDILcRWjJIqfLGajzX0QiQwiJVLwtLEbJ6Vr9u1+Te5UQOhi8t/0L41Fkj4QrIfg
4N8QIpfNelNBn7xMuftaJ8uUF+lX93amEso0wYF/VOxMakOG+KlY17uhMcR9QgalUg9+fqbNzx1D
mHbg4BbYnrREsQy8/ZonIAb1knCuRpF4R/8vPoSCkepJSijiaMrXnMSAQLq1Tdu0x+UXXkRjJ8kQ
nwMw4atfzc3HP1X9E5Y7rb4v5nJoVWUW/6re8MPJE5KPjtmfoMl2iEJafZeixKCVY0073FEkKnnt
NGNC7dpPzMi3C8Vj7B8mXhLVLJgCci5D5yh8rSxDSBI+wVjMPbpe3s96T8m39gP9XKuG6O3o9ial
XKN1VpbDSRPCFvXjTNvIvrqm/oQh4BMs7ZByNB3+lLXocCnKATvtZiReF0ScyIWmXlwB+gKAbqNd
NirLMCf2Ssshp9DOewf9jyKutz3X/OltQN0pqb3DD2u/X+lQXpBqCgo2lKzGJYbMFDN0G+t5JIGb
+oH8pMKIiNURmuppaKg3IMm2DHWOCpbmoKYXAVQXRH8LXvGvSJ/c/4MeW9Mc2rdnvt8fNtmVFvyp
FlGHteguzmDKevB5UBl1aD8Ue0HTLqAW+im5HrXsdTi4sqCYCk2qC6lCFSPiIVS1Q1yLLdlTnl/V
xDx+ZzVcsxbVHb5lxKGRU+/g1jWk/kTo04swXAoB/+ZgyBOsXP2vypZE5InTBozxkB5FPTliTEYS
IroICPPjvDnrmYm2kOBtoRli+d6uxUCYPJS6sGjgM1xFuL9rvK5hrlNBgsRrMoSFKcGdNZVTDuad
KzPu74PlkIvmYJC5mp80JvXudBTaNs7LJXYnblkX3WOuAS1VD0r9YaviF4mLIKIYNILBBX2cITz3
Hr9Yt3GQ5f42Q0sZ8X5TLQliHWN4boHiMAAZYqhnyLpMG+n39vDly4B4g4iE6MuHN+Hx88NLvS1U
C7YWhrsbZzyLIkRpnIe/nYQFdl2nPoxs5nJuYGGCnvk6CwYBnO1anA3L2KpFM5IKlD/r+hbO0H6r
s+tJrVYL0KT3T8W+lGOemyLcQr7qhuZWjVPswmyqTETWMFdlh25mvRgvRlgsJHCbVb56r4tkFzvR
RVKY+7zKkarBUCJ94mgufgyPi5hr+y4SWOCmgokBWvTqaBydSun/WGJN5E6fSjlUvh3478sXt0+0
wmz7YSLqZufoLfvP5SwbfRjNR2Ae7sXa6rnlt/cVAWSJ2d8fXLxt49klgp/4FAyxWvlCW6HALyWo
EQP2rNxXyCtvicRHgmdPnZvdiTzt2R/4ljZX1iuEUcOjLB3H5BtdveWNJ1KoKE83bslaGgWyDD/G
kuqarLbpUvDCpZ/JqLoz3oqWDupGRVfhO9s70eQY49Qrcjrc1MAxJfPgjY3yXepU9F5JWDjFL0jI
axvdyDD2kV3bon6tp0KZI7Al37aUpWz6LpN92kZM333QSoEMCTy8/JogbMzRPcb3cSsJmT5yG1/Z
YyJjgKpRxmH7uKEgHOX40CZHP/vNx7dq5PPwhz6/2VlMx1WdVW0BQ467Lio8N6JAMLYWbOlNXahg
NLwHdXz4AxHq2REhreWyubyIdTf+yfBJEOu8h4F5Lq0Q8xbtAOt1Uyqhg9L4H1EWjubbZE9rbRM3
/+7oqepD43K3XyCjZOTEX3+UKhn6fb1J/Xnph5kC5TWh0k+iwYI6LE9/5WZOpETTJMNFKHYz7m6c
fjr5XyxnErgdzCu7SDdDivyvyocUNUTggvK00tFrZPtIek5GFf47+n3BpvqZO2QZOo9haon4xH+8
kwn3SK1+XxQuwR4rMzTeRDJwtszoeRPLvixELYwVhGpPI0fRbeIeaQYwiblHz8STJptx8nNDBHgt
d6IXZcHhHKgjlVEQjq3MEAU1omRR256U9OilN9Pm3yqeQY1VI2iuC2SyMKMwVIjri4jY0mVlHoPL
utoWIJuNZEOZJVsE+fe+zSxX/fHby0K5DJSG5lMadsKHplutSc0sRJhNX2apNsvcIl7PaWlZAGcb
/yiclZUuxipyg7Amo3FvOxWd21FCvjozV6i0sr+gPt/w9/yE9I5Ba+l4yG41bXGN1zIQIRS1/XjZ
9LJO+HqdRf1xyhKeC9R6gNmqWq0HBRHI0KSnAevRTiwyd5ABRUOQ1i2nxVDepbHS1LtdYCUOwIcB
Mh46WKmP/GZAMlAy9oLuamD5hkr62/OPSa2deZhdDXrOPpaJIBvn3CPqw+tRC4SGywpIIHiwS82H
7UF3/LxA5B9oxw05RLDjhefFHem8J2rLKvxHxNA0+8ihqw+wvnNTh5c7K6EgNdFSkJSpnazEnpDq
xI3bXhz4DrNDWq7DfI0YjbCY7XcsQTb2JT6gJzfo1/xkOhVZ5T3aKlmgWT0gnjxmF4uUBWx7xVjf
6fYx62EkUkhYXP+aAKL2x1nEXtPmcUCMYeSdXDus9nB2FdaHELS42kpDE9ndmc3YzfpSXVZTpT/N
El+te1G27WEV8vEwGs/HYg0X107XO45EZzt19Vu5LDLsBPJ7K5hYye1YMxjO70yP3v4Q/UcOLdOO
3dp9gpqmvyllh7hD9AP5tyIeYCIxGaAe25J7SMwfTtZfVjtqaf5wsxguIqwdX9iYOL+KuPb+RIzD
9miqZN/GNETehA7Q5f3gaQ9rTSHcV+jF9vzMiGP94nL+rZ0t8/fEF2ouzJ6Zv85wSr/UC8jKQUlB
zoFtpQfRJ6YBWcwlJNz5/rb3lORTFuytQdzQuPut+Uuiiw21si5vJiWpc0ExLjTzjNTjeeL0zHX1
RxQWGSw8RJZI/XfHxtRuEH0Z4K38FSHilP0y7nGoAl6jqSrjj1BAnmQKTNNs9/biFLFUglLW1DiK
qlbi1EEb7kV8+7JK5qX1C8iK0A57A2ax8CRbfJQRz2lpkOlYVlkIqN+tEiHR46yHlz2gFhdTgPSB
jeiMknre4LW83pws2hGVQLc7grrJFHN8UvLiff5/yZS8k+zq0tjoKJbdFUSrSmvXl61OJP6orDQ0
4f2D20xeCqzb6VmWX5VzoYgUkv4SprYY72cTpETqREP6pxINt2RjCgWjvhD5Da3Hyop6KXeaxRKl
9+lH2gCRlDwFJCATDcQsj2P0PohYIC801DU2gtFOg25KTCas4MONnT13F2VIlQY2wNHf1z/rWg1r
FPgQ0XVACTczECiAU4lQmTE2Bqj/wPcrX36XrUZz+xYuChPcz6w8mF6sY0wMZTZSDvGixTb7/K6W
D5ic8M+tPllacJBvxtNvRvTM5+jG7JU10ZeVDNuy61E9Y9fqvqk5uNJewEhnXmE9ZGXwss5kwThl
hCOZAJMiZ7g2O/QnwuqfBmgzJHHaET4CNi1lRix5xCBIOkBSRKxmWlDMdB1LpibDknGDqHPvXYCF
ncxVq/pCYdWJBxF933BoG9gqep5U/MOd21l6Dx3I+MLQqzolxReA0ex9LalvBtRogTyzxfKISHZw
49/6OYTGLeWlE/O+eBJ2uCN33BMJ5poK5uDnBZpZOyeqpSEpHy1uZANGydB1oe4h2fA1exhL4InY
/XYSdxsz9HAilNWXfp6OvP7xeWG+uf960WtazhWkbALIuipuP/LQcSBJKsalZ7HYVxIrt88QnsV4
ZNvc8zIAPKk6NZAkxWGXHPQR1NAq42oaihHxGd88U2oqpNEnPE8uVEN2kapNKFu7gHw+KDHGUTKk
Odd9S3ddxZh/CiMi+5voReBuKxGbLLgHJFl4cfVbW+YPLA8NtJFIk7ArutIED/4xMm5cRYPn/Zfv
osVRPHj+a+DQ3MkSEQb3kuJxcgPRsylM85WyD+T+wcmtTfh/g7dgSu00B56ZA7sba63gX/DToszK
ibLd1g6ioDrdpe5GrzCp1Q910oaMJx0RDsIU/Vq67lOAvd7keJxumT6N9j4q957ba7ySb5sAX71W
tcKeVTSWJPS+xoII+xRD9whDED4Zx8k9xREoJ0LWofcyGA6BaaEC0t/BvWoqTfGLaQWvZYw/w1eZ
MzpMt3JNxBTqMC3jVb8PNJzp9yqmNVOCjSW4lW7DGhCtU1NQWIGvPB8OcWwrq3dZ30cLX5mNATYh
SSKgApLPKrUBl2V0J7ogocDPRhk4EiyUq7Yly+aXrFwAU301mtc3ASvzwPwEIW+58WxqsfxB/JaU
I+wf3NvmipYgQJmlTqIHK+G3MvRrbVh0c3U8GVdxq++TKNhLlqadedWYqms+8RW1kr2ol47MAw5C
NoKZ/4e3xz6zB4FWKnxvv2BrofnSBAuATm17we+f2IMLWd+FFEyUlKs9vwe5tirKoz1s1ggEemSu
ecJFrmD7yqRjO3pQPvA8yS4RAufkp7UI9j/TTpzJCvX09ewl5GybbDB0cRhZjLFmKCu49Smp0Cct
+OAU3/6WGzNGt7Irj3Y3I51fWuV1K+7+De7Xvao8949TSMCbJbrMCGOXfrD3pTR3sbeNcLJ5zVcp
bCv2e6BJ++AopoOkP0WQ1u8sxn0hsTfjOo+xCF2ZPUs17SDJFiftNDHZrNIjmOU1LfEhH+kCd93Y
SIDHsJC/L7twB0GeuEAlYl0gjKdtnouCm+JAzr1fcpDU1GkEW9iWLyEanEjkS1AtEfnrso7eeaS2
ysl4PUcZicfF47GjlYUoqaHiQPL1Hv2Y1szUTt06T4JSg11VcsG73h7ajyd3M6Gzn/Q07Xj6V+SQ
wuoM0JMb+VVxQPbRKiQ0ZFepSICh3K/wNEZfJM5pu9B/46NTIdmDt9Oe+tVoCgbFwDjrxtOm7nrp
h6uRfRrMqitrePUBHurEZcQDC7Spde5dpMZGiqRERPhSeOsKFodvbgPTKKsloSvvPSNqNSf/NuPl
3igRykR5f2Ic2zLG7kFITJCZkM4BiBAt0gLaWrwLOe0zpXd8Lf7EVuzLghvJJbVq1dU46kFdfDFQ
GnXLJaWHPLGrbZbsZPUuEcQlNTWj3Z9xOSO8I7iUs4GcMRma3TSxHb8LQVAImtbstM+/oxpvH0Te
E314S/8sY+jvjQBnebMPkYqtOHt5BJcPXOZfwdDvejcosoWBV+51DyBtHe8GtmtLORVrrCu8v5xz
uipWIw9E4aK1juKa2P4p5Y40yoU22Xj2Y72/tXrL0MfDM4dfrB2WwRhVwBbXVy5mvzmdCB9VPVvS
n7S7I+afRfWfUdEErAmz+VPi8QHASICEljaiY03c/+QpAhnp6gVNXT6ZJ/Lxv8jU486Z+bOu3Rvw
R12ApoINd+cvy5cZ0nDfd+RJxwuSEWmBO/PTBoXVbC47knEjB7oazmoMSzem75dWCnZOXQ8pnBDG
61q90Ny7W7VQutPMtrTDgCY3kspZbQDD7/YHpyqRc6xJPUdrKdcEnoJgljTCpWU3YJOoYMWRe+0j
gO7+TXBdyGr3afuRl3xtPpmsJUxani1dsxtTYMe0pwnUSby6Q+ef1EYuKmRFme6TDcfjzLOdxKJ6
gXrlDuoFPlUHBy78OPqWxhuk6CRs9V+ggKTw2VfrzJPOvAqNDrzoowK80okVZGvXpCjlCI+ty/aq
4JWJ3horTru8CMK5Ynul77FRNfWkE1EIufqHwnhZ7miiWukUy4PG59CAdRaMAGW2p35ts9hCJjhr
pgR4hvkOo4qf0n6PATL64sNzFROM9mWMSHa/e/9w3VxcOnz5w4OoAEg9/ECuL23zFbtRFyok2zkX
em19QiwS3tHtki59GjSIJUoD8vRSutOtMyc7tESHUgGxSIAA9kd72MpNmNenr7JTb6bpXrHpN+xX
7bTZw/QWEFBMN/DE2p++YSh2hT73zzdgHaWVub2viHb8MRrTQCDRij1L3s+pm/wVmLhCa6B56FNU
y617GY6lIDZ3klH/AtWtFUYeWsqPPZsxvaJuua6pTAmqA4YAXESLKwY8DB/4T/+pW3BwM1V+9ako
Lop3N7Z2GvEVDiNJrlQe56By+OazD11J/WoVC9XJlU40MTyJuGTEZknLidUMBUL2rEBP2SanscPd
qTvGb3JSWA3eTg6kBlSHk72EfzAfpcaZgrzcEKS0fWKapg0W4MgK671xXl91Y6l116uuz/ONzwgG
kT65SWbSvKM8O6/Nupu0FQvT+2pU3w1QkCNaGpKXcjMWx1yj6L+ZsGa8i4piJLqdq2yByzBZQNwJ
G3IqUoPR6WJ/9aI9KTsUJlkkyL85YhoqMPqxyYgprFiQo5r0c99Wew5s1A3YrK9ikTguyRV6m4IM
lUbKO/OjyZg7+AbRQu0INYAcIA3W0IdxWDBJd7kfxYS9erLvSsZmtuQoifb93Vr70niJ240umgh7
C/pHsgDFf/TbY3LBYWOvq5xwkzYGpbwZLRRbsaGBQkef3HdqOEoe4VJ+pcqx2gsT0Ily1r6Cof/x
ZLiAj9osxYTHGpqY3uR4P7T5Fz80HYT4i1jqt2XfzBgw3TisHXEod/yZUyEABtQ0JEnjh85tdFLY
qTESPbBHTM2bPwGN0ApLcBXgsuSfDTeKN5wJ4zTBmHmOH9DlpBg4AP0qstVAh4asXcYlcZZ4qf+F
1BpGeHqeGkkLL/aZW9sQPSq3zEZ/Jja6e0IWBq83FYr9V4QNMNbGvnMZNkRemm+2cSoXNNoQmTNl
gLlDJyB3NFvGk6r6wp0GC3FVdkT64qfYSnN6vsnHJOHFOvx1wYaul/YDjL79Lr61cleF1WRjBvH9
+QqrsTcKDA5UR9ViAYM2zOQdWsalcUfsx8aOXI8lSUc0VAJktzmZV2jeCv83bM4Uy7dns/rzjCxS
PojXEtJrr0bygGGq0o4fRg7eERR0s/n3PI9rGQQNMIiSf7DHmGfnXrDkik0XYb6FV0gY7qPLqaUj
bVa3h0opt3UEAmlZaXTUJjP6Qon4jRwQE0166F8ZDYtZ6hu0X4xhKk5UtSE2Ea+qUt2fc3ATRq5r
Hut0cHW5XS/d1MDDfUMGsxM3Yw+w6iFOpnWuB6WrFuz4G4e3Rev2RjMg5NhgMcRZWBO187BQj+Al
OHCzGsYfKTN2W9en+GKmO9XNgWXPFndkQvAYiRZ3pkbxWCu6AsMwlvSGoGKO/pILthLDS1Qko7rX
tuCZo12KI1EQ+Z5AZU1t8BF2JXzhYdrWvG4Q4kRbtc87Ob2KRuFZJwTkVQMjT2LkdeZdNgyftgv+
98qyg2XozhYF8FTeIrWXNbegVPL2EsbNXejf6QMyRjRPspEBb8C8IvXC+/WqcHYVKxI6J8nowl4N
ioc4jRnwBNxQyORSasrd+ZwBTjD4xNZUuqmJM2xPUncVuqoKt/GoGuJesmYu0sgfNu7QjEn1b7rv
WyHQp0LM3v776ekU5TBY3++Ovg7hBaExypQP+ouOyYWfyBZHk60EjG7+F8UikgS2aOlDTfAHiT0S
PWN3//YvwQjYXGBJra0ZbjFSOfp0R0BQtYCs/cBwuTVs8spaRLqouEd7xMTly3Jp8ierCqP6uwBM
Kn5haaFaLigTb+lPxFNPwYu3aGLqVtxf8dbHqNEikFJfS/uknnm1MuJxvSm3YGcNNYfp718MMAMH
Ck4lOT1ffYLRnVKljxZQsk3zBLHybip66OJgAULON6U9QTCi5zpm4+n0i+bvpwBrLBM8HBK8jimg
Yq939eA2qDvcnWN7YNsmS552aFuwZhAFjXOo+lqaxisB3jYlST3ZltMS07OWIg0eDTSfeKox2JiZ
xPVozaTPLR3RQCDpd2fQpHTlqarvLAjADDj3vSi+hxv8heAxkQ5bUtYqvayvzSINrS4oxeC6D09R
9D3rJRtgogzl9aLc1bO/UyVeetZivRe7kxHnx/RExPWJ/9r6IWvuF5cJYkSS3d3NBEBcGEM17VF7
/2zJFKREzhwqlTJzlqkB9tzFD/jAUXkaropL7Xgf+EsffzTHUpHXkl8Ys031h5OudU3i3NPVmzfS
YJ10onzUENy/rtafsH6EvC25/GOVv88lLv+jI3W7CEtRKm2zbGkAhLUuykhQbVg5yAG85J1fFlNC
V1RRIvX3yhsqLVm1ccesU+980bX9Lb708lB3uLfAsf9GWwDUDlt5Rs8uqgYK2BQqLN3npu7iTJiU
cXEGgh66tc3ZrWDTrUzeC8dBy18IcbH3rDPaR/F5Kd9TkPo3UFn8KH5MjrRiVsLflkm8xxGp/rj+
t/jA/8d5nn/Elrfe0ZPpE9iAbkXlSdcvhAnAiZ5XzL/YcPoFra2MJW8IamNfYirRpH6OExIB7i7V
N87dUX/wnLc6RTMY8h8vZ++x5PHZliOCehT/pavFU4+ydVi0W80ayEBrorgxVP51KVfMCC1Fhxd+
qgC4laIm2DLgsDQtEIzkXT2HldiYb+ncz4zJqfRHpPk+67RyfuwsgJgxAHjpaJ0osX9u6i7udpwD
CZdUzLxE9qW5WIVUO3OkWVZlKdiD6/T1UQpcaGmEERTyU7WppDx0hM46ogdgXZmw6zB1bBtrZyJV
ptkRi06+7P/drOsQ15pJCxMNuCxmmTIN47+JwL2fNPSbCU94vM6+27Ei8TvmwswiA6PnTfL/ssHw
5ZGns9njiRx4VPM4lH5ZpsqVqyWqkwTi9iR/NOUW56e8Rg5AtQeiwkaAa4NKpgla45yQFvM8RPzC
VfJ16YMxZ3fZugywPkZGw+w0OyJa09JsAYPT8xOxO9893J2kYL7gQvLH6kWi3DND6HrzbR/2WjHH
84duWrcmDz5gZP/ltZVTHSl3Bm+BHJJsdk7Ol0YUg2kRaHQvCf/+C5H2I4/08PFYatHxUNOye4HM
sxjQs7sRWsEmpn5nB86JYTjpRrWw0vizBa9aMA+fjOI110h5fvyI1CXqszTs10U5uVuVFAG5MIG+
Y8JY0OLE7CoyRkCTRaZPpaY0SL7VtfYoTUKxph98mw9BWqkclWdbtBUhvn2NwrknoBVPTHkQAL4j
DCSzZszsQTD4XAq5hNhSKsGW9w6+UQEgCZf3iwhzFRauuKFycKIz2deysO5U5azxmRQ12Am7m5Ij
RUpjOxmJ/fuWR6oQ2x94GJQLGom3wrR4J+pNMkgHSYhxEE+HnzepLVT0f0ZXTvkXJj5jWKKUY7mo
xNP5kgYyXsQQftBJy86vCaqSq+I11gunCKeKUnn57Xpb7v+2g6AXXk0OzeiHKKvKFDgwbWCCgb7Q
OmSrGJms1aIOkVOeFg+oU6Q3leRQbSfhQBpoZcXqjX8X1UQUAe1nSj1bTIJjTxUdj72Vcm8caHVs
wRTRYxfI+Q9UudQ1tBcVea0ePZ2NnWyyrRATpYjPf5XSs42DDuLq/ZdcW+e2D4XPtRvl9B+wu6RM
qsusI+FQnOmye501ZgxEdiDgbA7EpfMxRFKoYgDFVb7Q9VEfOJf9LTT+/F4osGN968npRj5YW3uu
JL+n1CfZi9t0s75dm4iVbhoGderZrYltX0UxpjUMJkBifL/9aUFyuDrS6eI2sThRdSZOY1tQkI6g
IsRtoWrX8+YDzB07A4k0B142L/0i8u81J+LmumqXi5dUBmPQyD1s9KWbAHd/uC7zavlgjgeqdiVR
UDUi096psV6uB0d6of47YesMm8Y4t0v9VCiBKG0cnPkNzLndNsrWV/3CAF6u/ROMOMrrcfhRFqC9
Pj+uLymhWy6dqlewAgjwR/8/R6TqC52c6E2m09tFzgbI//WJjiBH9b5/gJjTd+G6UYlHeAWkXxnk
RJU9DhlaeKkunA00E8rxA8M9vmiVMFe7qtQHLP5y4zp5AUa5gLIG3LwOuGm3Q+s7VAf9Xx3vulqu
1AgtwEEKE1jiCYrrGWV47+GXNMlDIx4ER1zbXdGxrzL1StyY+53ozvnmyiLdLlT0kC+qndsfRcK/
SDXy/MmZzJcGHa9zno5hiA/7v1edSEFqw9gcgPeElPjPhRSPWS4XJjFu2q3HW2FNBuwafYixdr5u
lBeINSlZ55xUzx7ltxT0T1/1DNTds3k99V3aG3mRi6v+meyTEASjURwtP1tst+uE7JjwpKsyjzhJ
eBrCTovUEpXqFPG4bXoXyUOZaScMXu6IUarCUL/SJPE94BihoP6Hj8aRUj9F7BEglJJ6Cfd+Zk/+
HBS7i/n1BIBp/HgPYswGpbjYpdL/LiHijrzRxVPLHa7/pim5v4ACUcID6pGUfNPI4yV73L61zHjr
b0aHUuIpdkTLbOUNRbfkacqiQ3tNftQJrcn9jMLM8KXS7VkCuyq5Ws1GVGI34fFhB+on5YpwKfZz
W89+jzsjyUEYVmOdK+wjXrabwua1PQ0M7KDrnKVNpm57776ZhwykM0QJFqCpocahnSvJlI3O7ZiP
OrBVaL2fGtLpDSbjJsELeg6hXib27SVcemNjf6NScL5G+3iE7FYnX09XLpNAkanlEEecJ6xkmjtF
tYshlg9MjYcrM1o75z4b6K/iyD6STpU/GqUCjLDq7uxQ1dH+8YETdfNv9wDCE0kz2qyyZ6Sth1id
TYiOfnKNf5dZiFfzjrbNzPoS32qnnGhzJ4bSORipAb5FLYVUbUdSoyr3Sw/PyMbzr8jQih5gsSxs
MqxEvcXb5iiw3ip1fszrqBNEXFxdiLg648eADzKm0Ifc1ixCqLFy22xOH0vRhSX0DYNMRSq8psIu
dXS+hlkTXrF8J78EY4lNqdZIDdQ5RkiWCkHVqR5fiUNzTFIeOTzQLHzfJ5QTKgwoUJvU6pUM8IKk
4zFgYuavRzIJErVDHLmM7lu4/JU/pZRmwuFumMGK02xcVXhI4SAOCL2pJb6xnAoAcDti0yljFweZ
YXxBUqwf88y5YDbuFA3H7NCajf0M6TluvGhoMcbaqyxI3YsPuyvvZ24v8RLrLpaoteBWezXRDMkb
SBd4oSDb3zo3uu3bAz9EcD01MN7YAJfMAZxQjF1skvvh1r7859zdBLpTJZXAXoa1mIvckuYtdCcW
+58Y+KxN1l1lBXgUD97CMNltS0Hn7cLbUjDfpIbfyx4mKUzTZKTi0DWQejduVd50zVQKs5njrUSS
T40cI9KTsyAqZgrdPBPeAIoSIavdPb/VGoaYZ1IDL5pL8oF97grgyrpXGm8TXOTDstlM98tTX7YA
3VDwO548rk5bXmodIVWEzMQ1Z5sHMixiHJjesh29pnDL/h6GxKS2CIWEfHvmzDkQtiX8z3YmBz1L
WEhMwQ49XgMAaLYYOo8E1CsDbLd++wforfGYdS8TWMeTXnBEDVaMZPgiME93iiCQTLE9TPtTIPuk
1HrRc2a1CQJLkQ5mfM/uvYJyYRPIVQdKHIJpYydPuLFu8xAL2HaEbNNYMlFmi12AF1XZy1r+P34a
yS3bvVn6ZXeWOSZb4oT58nOWWr1ZNnImJsVMd59NumHggU438iUJqt0YZfw89rki1IBHzSDA3Sw0
JEMZ4QLOspdk0zUU4zfaT+9W+Vu+Z0KW3JFrWz58q6Cqj8A6ayuvTBJfH4rFcXNyVWFC1NoEebjq
6nyn6AawswOgP2RcxPkznB2hre4FZ5u/wSC/azBE2f0BIUTaS+AFu9L6Sl/cxDnX7sY4J+AdhJX4
ad4b5PThQsgo+nz8klhZD1gIKvRJEydEZD9/NzlIHb5czyMzjlvAQ7o8p/Kb/KMY1rzqImftzaDD
7zmxg9nTLZY6lB6CIDCNkniXkAvzQ10hi51mu8B5WsF4S6Bkc6ETKBOt4b2XxFiNkPFp1G/uKeSF
2csH1ETHuDzy9txgTASkU+sPGHJMt8u+SQPb7q0bOpVIz1ALHdPvtw+pwknHQiLb43D34IZLwdMK
2N0tyLEDWoKKE0TVfOyWFtVo79etJ+2AH1FuDkq+gBBitstymyfaz9R+J2/EVZtMJX4ETTCAd3YA
zsO69SK1HUlQDKjQchP/v28Di9w6AvDqTzRhm3OfQJTHevDzXmzzlIPfhRZbXEVyurJjZeoLi7+M
kIW9kmd6ajwMDj4gppSdtLiOOAw6etIPiv2kZeWObsn8kDeQMKVZFa65n0Q/Y8RhvnbRk/RzdMnR
DNTVgeNi2AvHsqZTKO54D96JLgq6YDgff5tON9bl8iqwAYCqcMgvQqYESLl4GTL8VldB4uj/RetZ
RrBbO5CuzcKik0/xUSDxegXyhgKiXlkFftyW0eIutnIrXv8YgomHMtqaQfx6ajwlChVUmBP91sqc
mVOA+BANpo17erxeOehoM/+i329p/8r62dteJK4cmp53QIDY/LxEA90C9IQAM4De81MKmVP8oV3x
Ad2lgsj4Ac4dJdm11yDBHb+CFJ8TuEQO97z8hcpIzuYaglKkMQcnhXPBq5ult0u0UpdR3ePOwxD3
CykB7zfBBHmy50rkUBEQLagmozlncRa3+n/JOmAXdu+ULIumr7Nd9JKMVEaUG3wPIGOJwtHCDuOK
Wd5T542VP4zaWcMU39RXEPttHPnqZzR8qpvo7V6gqVHJoNZ5Wmzw62k01XqfGQP0GfO/InlLzh4V
t1ALhhsheG8DdffcnA7+mQOPF6fdoArVzpUaOrqfpzG6E8KIDA4Umn6gLFXAE0InTBMQQGvUP1b6
mKHfKKQED0h2uyTCY8m6eq0Hb3z2Jjpq25t47tkTcQN7mv66L+0oylZZPvXJaP9HZ3qOHHl8DaB+
EcRSnDSeF7qpGnpvvlpBI52gllxxXRjbWRts255a8EWcSQzs9zqKM8cvkobxffmKqo6tS5nlWrmT
dJ2+PTTurzHje3LSZqgfK/N9waK2XfvV2VG3PCeG7XW+Scl9hr1y+tuS0iJbX9eEAfQWMc8DDQ2F
wXZ8Vu5l4nvFQRRRd9noB0UBcbRM+R5fZeYtm2gDTZgXUZ0S3RkLa9Gve9usTsWT5eE/E0thSUGw
PZ77KOq96NN76lv8vvcd4RP0wuRZ3iMpmIJVQkA8at+KSxjVUWeAXeNl5lpKQJ8F5FTClmX5ZO5g
rlQ83kdNpqrMRmpMVPgJ/rah8NuZvmW5QIIzEhAF+L93vvBUIn0LdVbOsAdbER+B1+Cuw4Jf+WHa
y37iAomzUxy3V9i46K7eM1IAdhVi6GXHIl1BaH3q3piSmCasG2D44bLDdoHtSPqdE+Fl/A4F7wuk
G7Ub0CNYhdafPzOnpwCliOV225yDriFtg1iSlDLrgDD4PZ8aazt66ma+9HSPI6K5ij93i1iOMQ8H
jsgXphJOxW0Fl0nnVU/LtNF4kI9SdhA8/31x7WtvMbzZXHmE69NMg9vpHmzhaVb8rLWB0xz7S02z
Br+ZyRecVJU1H4ggb3hDX1sddAaUddyShMR1b1nvixKxMgx85T1sNKiuTdQz+Y70rfFkkggHOy83
i1ZunguFkydZFky+9kHiwJ6BBatBYA9vxFJ7/WJfIw+N3tJJs7W3Z0oi4P+pzlSfy2ufSRrP8ZdO
BlEyX+cfy1+yxijrz+j05vcrZKXHhESSWPRSC2UaV7zHtlcq3y6tVgGbc507zfPItU5o32q9SZhD
K/h+ycth0qTsEOj3aXIT0lB5Al8SRF9XgOwJNVU9UHPfLk7xxsrp/uNjtbJRzQ4xgzHW8Xfc/krT
n+IDpK7TjiwD8VCT+IAFUM6l0JgeT0TZsck4sIizi5jD9BcsPON1VJAfe7x1RpxMqi00JH1sdPTz
F2QOv1hWkcH4vJnzKyXUFbTP99ESmjQJ67egIbP+ycyhdYoiYBx3BpgZi7IN6p3KuRJVYifyTbrU
G4wPUEXI5imjPbMVXfkECTR+SgoyPkEJJqhy6G2FHDsBsqgs2dA2PpkJUK2dX8BPo2rp1G2zbBBK
r308r+0AJc/02ByDkh8TkfvSaqsPb4aOuaE5XB99T9/FPNnDLixJZGzCQ3u+UCYTHXtG9rxv4B7w
D9iKdbzx1/HjST2fmNAgeDxQwquHy9aCJJQtAE1qufkRMuB4p8/6sz19GCILAF/IbHbGG4zoft4U
mftEp2QuSQSYXSeJxFQKm9rim3ZZK1VctXJPDrWTtnxqh6VumWGMzY4MwwAgG1W3AM+67i3UZypb
a6P0+iK46RDSwky9PKH5LUcB4JhU8cOY07EHEyu86U+2qCu7G2Wk+1L+0Y/BExwVPLACPgm7mu1u
9SmFlFT731CVWsKeWWtTvUMUnCY7LFusccx674mDAAknpfo3/PkEXX0i6yZema6EIwsa6vIkv2L4
vHLCF1VjU7p96VktObPf+HtaImdvR4qFgQZoKjR/Fh8noRKpsI4OaLVMz2vcJnqjHogsTGythUW8
9rzegfej2WgBYM4HXUcSXFnE6kMWGD8WMcJAmzV8i11+VmEAxFB4tkMCSi5Q+UBDIyf65ZTYN+Lm
TLDn6YbeVCJ2q92htiCzyyfbCFA8yBJMRjqEZkMfh70BZNq4GsEafNSqpAnlX85o/mdM8+nUutgt
0llVOa7sqG2fVm+OSITPuAnIyoNWhmJHd/69QgJ89Zx82hDrwqKcPYFbY+FO+CSMh6hr79v8OoPO
7tOZJbQ3f+Wz+ThU3Wk9U/1h47qTOrvsM5zs0pWECqLttook1V15U6KM/pO2QLKopzopLwGxYACR
QTItfkgM88COb5zxPlyRQzT6RHGGkUuDyS83tECFCgEVmbvdKQv9DeJV4pShJeyuYbOmeJNtYkbT
+34OLVx3spPLotVGrnKVVhcfyIHoqGWeGO4nfeTMfBkEJhDGE4rDmCuKvqoD4zU8Rw+Gvchs2x2q
kyi2oyQa5ELZ4WZ7knLGuW3+yeVNFGPFfJ2HFO1e+eMX/Dk23weZ3V5PD5nEJ8TTf6lMPMUHOhLb
lL7b2SN1YPYh2sOD2WX8s+jX/TpW1M85l62CEV06CnfemteyWO1AztVScx0zsNDkvGZe9n19kJAy
9jZd3Mgi29sBqdQctn3LTAJ4oHb+1eBOhbd7OBITi21lfBwDY3Lk/JJHLYtLjkMczQ9/AMkfOHcN
eboNF73mQ8bTZZoLF2vRSvsoXZvs+Qgq05cfPrxzuIk9gV1z6eYvb9yLHlPfaK2+suRYMLCChYVM
DlvExk8YN7SjmIWHiG6ca1w7bE4Q/gjA+nGr0tlJ+gH8pCkO4dlVASaGZBrMVx/njOfOqJWk2ArV
1/zJWpuVUBKlcmZEGKUVzDdR+zmsOd+C289boKFqIcFOwjht8ftyDmaMWh/8OoSH7SssVfnMvSY6
6QKpLUGwIrCdKcLb/K0l47hkIjUE6Nu8TG0/wqUuEhEwRnqxta56koBJvez2msSt1khWc5xfszjD
nKk3DknXmBnqGS1roDyaZ0c+cjI7ufwqNajyPn3aANGqWLC/HDjpQ+wHgvA5FGmo6JjOkmTDhs0u
wfdmrQmm6erJjvxAjQ3jRDLyGlOByydHcJjnv/X6bRD9hSX9ZsjujaG8eivrJsBkrdwwq+Ajzv91
kARaibX+z0DVXNl15BISNjRNSp8fncDi8DPhKn1GwQDZVUbkwzfUoDIM/EBnGMrLfanTzZyxeMNx
z8MOpE2aCMUUy28WNllRz8mRw4NyI7Mh+h60cfIulhdpdYzYs8wRofiqoPFAJeHF/+SISMM+oIBt
27ITym3dQZqcZMl6cOlSWDCSkm+cjAagDZEZK7NCxZcBuHiRTDJI8wuW6zjEGoSUcrsMq1SdLyA4
+rpUwDZj5xWVHxrmk+Rqq1pIbzuMx8WHZCOPP7OQM9N+wl/TKmC85CxZVMBt0ZAZH4OgVMd5Tard
l1O7FFw+mVCBJT6rqVnSwr/oj+9epxDJxxw72ut/CPr5Xu6U0Lcodv8tqMX1lf9UCc3/ot6hWZbP
wMQjlJio9Ai1WwKtECOPW5R7kWgEMzNnUy1huA5NEv0/y/PBoUK0LuqqRYbDxAePBmOdw+cLl73t
KnZ0tH6hIkTOY4862YShda5qX5zyyfJKgo4GCBZwKv8WTaNmAu9jHUFimiTdUbvdG5v5YqiFkrUa
hA86DEvek3xHzMoZoaePuC3kWVgqxCbSE5nFXFzHm7sLGbcJxdZCQJhl3Gu+pnR5K0gnwDb6AqFx
d7FgWIYw8PVCoBwXF3tbreV+JlpALZ4rp2LF7ypGLF5YXkMFOQx5hi0o4nMJbvxua4ccMJW3LMB2
Crf5VwAGUG/O8EOmJ7k33UrLU1WLlmU84NgxwiGgD3AunmmOlZixRdASiYolykWX6CeYL577AhnK
ug89vJKMHa+YjKBScuMstKsuxDkjfYWy0UQiqHptqhw+npfhwThtSVes7lPE8uLBb1KUWnanEKVz
c7Y/BJ+V7MTpQB/lQm0pEKSR1s8BJzpE8hRV8fbmIx+8/ZLZ31VF8fJWry74rs8r2c4ZT+p0nR9w
h3/waUy9vgDmVgEjzQM/Rb9N32Bv3DnajJZHdaL1gHDrlQUQkrksag3xPXVLSQhgUeXkc1SWg4SB
nD5ifeeCY+mha8gtPs5BrOoqC4i3GhlAwozGGWoNU2qYTQeOKuGjpvuwzu/7grRXWxIZEdCwKhzY
1k/wdS/iTfrz2QrbSI0++eUmfhF6ITOROeI1mgOtS8Tjpz53lyKhJTTo6nfLZLAAWpov37L/AlX5
itU2vUepiGQJ8qJZ6S9VXvdgY0RpS4/8pqbtF5YHnofQ3xJOoMZIsWxh+VD1+uEH/WOpFi1FDA1Q
wqy1tXbhWFjQ3yVrMPTM/hIwxtFoOVHABNkgB5tSm4mDTmdtmT2psZrHkj6uFBfUl8cqE/4k+s+8
LN+gV0GgkO1DEcX6LQBDRR9I6zJT8zuRrtFn8Hmoz8KJ+07j+iw3nlzO2NMRtoCciUSmfoC8OlvA
SNQm9dCT0bHSeOcSVctf6leNa09SNGiNyLfPJl6UUdDpCIkITpVjkfKtZp8wv31vwkH5ob57XWd4
NSh2mRycwt/SfHit+4ECkK/Ep6O3E7IsIZtg0uDVlrzIVu1J4Ron2sMrTsT22J99gZJ7IxuX68vV
iWVw4WIzi5HeJEz9XeUgN81Gp2wX/0UahkUYVqQNQmYkR3VnolngPszVMq91teZtds7AGSQC7MY3
kaoXfpwATkXrDq+0EK2D6RbPcqi1pOw9mKzCaVCTxgbxtSneSwQt1f5ELY90G7cN3uNJpxvl0prS
u5z9yByQemNo0wO2+li67z1at76ObpiEgnfV3+6JB+Sizj4jFwfDyk5HcFSuL9RM6tUwmfrqGD6d
wkSknVUj5PDgjlMdplPCQ5/M9pyntj09x90XaE5eFZJs3+GB06W+ad4zqItQwZDi8ekjkll3Ydj+
CgQop4R0qm0hgu99diH9SncVepbiKQYIAsia7Myn8Db93hOXUrItlg0A5ZBHPWsxmUSZXfM+YDLk
TmTh1mOKXOGrCy7zev+gVlDJ1P0NxAB7hDWg2XdE3Cbbm9Nuiku9KCZxHqqR9bMJoF4xMHdj+Qrl
0ar825njbijqI8lAlQ2fcfyKqo0tVz48I8hxuJwhPD2yLUko5n9JlDQBk8/iUoXJRicux9ZhL3Br
xfwLi6qbvTLKHjIVX4UXwd7gVLu7h1Nf2TyfZmY87v2o0xFayT0YSq/ujDQqzbe0168gTUeZvVFG
K2jvCcApD6BbCkXOaYyZQtDbD3pIeh7fDwoyiPXj6BXEmYoryLxdGmSn8vjTbij9wUuqTLL3Eld/
/3kY7Zm/iLFi6N+IKdj/2iWNMNDTSsv1BRcOfqkHFDLPV4jnjaclSUyK28+bTJ57crqnCLAcTeqe
QtihKbb39L0Cph+0GlyQ6/xGX+LEzXdW3FygIkIi4kTMUapUOtE+Z7CXdzBbEb4XsfGycHFYtnJ9
3bj4TT/fmqr20q+AEDn0gI9v1b7giNYZ7yjqTngGRWk3Mvl/lkoRP6ie+Nj777h6bIFNm6fkOLKe
l//lbm50kV8FAG78iL1qt1TdPMjFWq0zYxvE5rNOP/Opl6j9H0nKfI8+ZzK/7h/IJmHoBhG1mInF
tQt5CLt6V/EcKJnGrrENEotSVGBhcas6QT2ROdcSp6dCMQKc+je3F40ysdB+QiiSQev7BDmRKf9U
XIbA52QB32JCoynOqnafXM7jFmhAWZDBVXH6B99za1whOp1UAQanYcf8N5f+u4FvZkWZGFYCk6yj
+ZzLS4QBXf3AyKc4hxj/KfzTJyJ8VG2xuQu6kIRFeAKMOKXxjlqlFkObkz1VaFovIc5+LfvZa6EP
iPQQDhNwEG6BL6e/MZVyw4Ju1cq/os91bPE/fUDWqmvm4mG4uEf2FtIwU6misCHTRoFoxNx+G3Vd
OSgRDUKXvYj4CAoaUuyiMDq+ihrgw8fYVKpxBwhqh4f8szu/nyzF6snMRaa+h2zoJV2acjXmDhn9
ddKlqfRZHltzRRshyag0Pvm5Xvdouhvdxu11pwJ4wV8q47CB62+G1VhLOjYIZOkPppzSkThAh59W
D1MdKiNm1Pa0EggZLljqocnSp9AZISjwO4xmmO5i/YBMisozGSppL/qJ7doDLTM6QLCv45H6c3cV
8RqldNaZB6TIBoYfhJdh8CNtnWqk62eBMC6Nn7wnJXASVOv/xHPkwL2FgdgxBHa/DItPgiG/Xq/K
DoG52lQJrhm3UES4Cdeb+S4ih1oEZh1lj0SDG+xiOF56zVDc9PIu7RF3My9QSWtCZjVPuixWxfVv
5zwfIaZCreBGda2Gcj5diL/TjpFxoa/x/l/KibFL/Zejko+4lzMT1EkWCHtkfKS7+R3sBtBmvtCr
R47W/jsSBgF7glYnVXsQnYvbdFbS9dbZgC5FJ/2tVKxW69e2NFCTf/Y8lHqBZtaTnkKsk+80b5fA
oHwKVU5Yib+0IIFmLTzKnOI7+h8NR9FLXISUvYuurdAeWxsJWrWmcKbx/DXkAH7donpgUICmTO+W
6geW3sN93vE9l8Mn16FtLfhMwiKPUTzS5t5vJgw4sMDgNxpXYgbjcbF7YlbzRUuu8rFsXEC3P4rq
JnrSfuGDZoLYJCez1D3r0jdqe1L+3f/spncfJFvS8WuzwZVKOp/nZbuCwVdS/QnWyqYnITRzfwUT
Gy0Lew03G2ipp/6FIG6el351FLF+mOp1cEoW3fmwHRnMoPXTi/by1wSVAn5ojZphgYCwv/wQcpGC
wve6mpx+zcgZXmDmmde5irQD69PY8XPjin7e81u78PR55eqAKn/4JYdXV3+KzsA816A/45r8r3mV
CqdI2lT0T2vvlmOSFtZfF3osA5KjAnyfuArePYa+iI9VW48oBr3DEYLS0thzJWlGMo3lZPUuRDoO
jL5L1mrQERZAWKMHXTvciCEJ21w/oeG2XZsEeflYRuWJpP967Ry1eUZwFA4ca0FK/isMItbXTMFP
DsTDOPKVTr6RXvvSwkjlZifGv1n3/HJ2Rf7AN7ZWiR6gk9xIYJPLCx/zXyhA7N/hfo5ThplqQaqk
zvgSIQl6l8WdPJwDsVZvPN5y/VPBuCM/b8/z4A/oOZ//uWwzmi0ZJkNg5aXzp3PZ4xcIb82vejKw
bli8vRPifSwTP+Jiw8IVymmFiBuCaIH/9oED6nQ74hGi3PAMZgEDx6bENxSLNYgg/mu7lujvp/Jz
R1Ke3Ab0ZDUJo6MY9a6c+z0gmHffpRYhQjPaG+KBdfnO2UELuBZtA5IHW4KcwCnrM/79QPTbOMMf
us4a8VHOqjwrzc6QvTTGOnxM12uaETlEfYMHV2EOH7YjsB9ykGY9DXNq3MTbU50ZR6rnBG7k0mFJ
I88pX4EQNBe82XyNcfEeOHZLLUgY/RTwRTt814xAVJdSt5UMQkR/sTCfrT3Vmz5D5nqCWeM2mkeo
B3IeB2cCeX/T5bC49Cj7faKivu8R+lhQuomEIuM8pWYbOxxW669cbogUzIXOAheSuV9RX7ZP7CfI
b74RbcUWwFuC8mgkxmV71tGxBlPRx60tRGhmosCuomR8R+6z8JM2Yh8l1uQ+XoJtWgk8zwhnn7im
/kZj8v4tdtIttAO55lrJf9s7YE67KLKVYVfxE1qJZDIR9X1lIdGlHnMg2KvYmtri/Mb6AcfJ6ohW
D31dNqVVPQI0uzr37icYnHO4Fm15WLwJrbXrF6WaCIQR6NI4DjFLv2INmvI2VEBtvnp16y5QPrCM
HxQQ+my5w49tQCLg9TEmFj7uwZ3/1KQtTxJ4K4e9Cj/4IfdITMiT6VTtnmydqBKxhPfZEtiOqAxW
7+ar1K1wdpioCnHL8ckD38LAdafEzEePXN6VhgaH3MVvSsGeZETAXHsbqt0Y7SBfreTkbyMwGnRm
K4MQZNA09d4wFuMWhNYvlVkYlW3xy2iEMop1O/0yfgG36Dr0uTnTxY13jsSJ4DHtB6fQ1ZpKsvBi
a1yPdj43uWcjIX5QA+fyFKAjVyvpPBXKD4xe+w03zifKzsZwFcD/GqiHR4JuoV8U1aHDsymsxz3P
mqbFIqL043gCcpZbLw9OFOKBZSnZDwSO/kEBs3y5ugtFIVWS0hvg+jz1azGfvaY+GWQwXyvnYQHq
PPWob44TCHtEQEJVNBXbgnkMBZNDo0ZYDgutwjYDQvvHlmTGMRcC2MJbYow/Zpv6TcCCdXn6KzqP
Ii359Ziw6s3N4UAV3+G8glV8z9gVCfrXexA5Gx+0aagdxGahU1Rm2wCLXqjH09PVkdhUXvIAUUUQ
JNTwUQqiam59tlC4K+hEIy/N6VbSjEn5AHN29d84FpqOrRpP3RmQSH/R4FZisUBzi9xS7sbnP00q
VdGhkIbJOW+V7b2Iso4IBk10cub3KJW9X4sGLXPcoVYCHtmYLcVYLiF1bIOM/9TSlgV/0y0bkuef
SBUhmE2qIARAPcV3sAB6fzWk3qTqoZKZT+9gnpSsTSdLucRDlZCmTo1PrSHQiCvwrMYPwBGtv1Sp
FlNFrIUzKTBb1BCA8cmwO1Uc3piJDf9ExZgFWGDJRAoahhA8Qg8U91w1IkhItpH0mYjdnwyCtqQu
8f/9IeiNYxTrQRxeZuFCYIEFTUtR2AXPOJ7O0FmAHcOXqLxDzqxPzP0sM7I10CsOSDRPk0dvGF45
uKsFNcAhhL2lbApUpkPxDPRDCtQcVK8ZBNnVKFjTHCGu39zmBFG174sGYD7Cp4tjkb8aHbitT4kb
qbwTk6r3kPJeLmHcqbzlujCa8TWtmT2c89WidZX+y/JSF4Eq7cIgT0rO9Lp0F9eCAhjvZ46qHfc3
uMJEe6cwmGuuuuamVgX3PkQ/c1UbnuUIv5YxRwsbnB8Dh4d62QT/3aBQm4BbwSX2vqEy/VUEfaj2
wCyLx5dPdVSS2prwzmNX+g2JL6pvuq8QZNlS1+qp8AzVlUcRv3xSVWdxtlZnYwceV7z97s7WyA2R
Dh5RwpWFa7BC14WpCRiWuTAD/v3LtkxhBond7DCGLJk8XW6aMHNrpDe1zuWDdIVzO2bbGhel1df7
yFo0aQmwwWFMQIJOn5xK/7c7peEfYdOUMww6uT47OqjSb2z4CyJb2iAC6oDkCdsbdB50frBayLYQ
pSzKdD5NbOI1Rk0rCQEFnPphMtH66IQqAd7vlXOz7gcFP+sGCfPebe5E0+n958I9xJFGPuRgFUPU
J/hGeTzUI2+ccgQb6KwsLOXg0xavIdQ8YJFUorfGB1S9OHkxMlRF4xG+0kfJLKhItXYc5GbYsVjr
oEMRlBawhfxgMMI5hGmwi0AO6crj9ZDSrxf0Yc5FNVC8ZnDekz2zDGnQv7HHmw79Zvrguo5EigOD
0DZa5vUqbWLXSAB6VLEtP6Ik+VqDHGkh3czrSdYcFi/qpuX8cFOb7UWlg1jUqggLK3mPOhOS0dqF
xR3bXSA1wzzVvVbqFmE/pfKaZ5JaJSzkyTRMQTpdQ0BuWzNj3SoQOOYckbz3BToy3TPzBBdcyN39
GhPS9IhCNlPASW2HPZIY1Vxiuj1aAflOFYcXqUDA5ekkaT9dzf3fqsqHNo7F7RQeKJXtWlHxAgPq
bTKv6IZWd8T4/G7DmhjQK8wut3T0Rht5XPx2pRdIPmgxZJ4Q46UgVKrrgrNocfPc8I+ermwh9C1P
vn5QkhXx1R+wfPJ44Fg32JbHk8Tzo2bZhJGd7z2vWoVAw4BRu5vzY6r2w0fgGjme5g+9VlbEZttE
vZv/7q59qjpghzVITb5tcupPaci/RHUmcQcPDGtDjf13Zi8e1Y8sFLRhEpP2kXVgPM63e6WC6mF1
xCtPak7f9eUyIwz8fMi+o6EyoVuVkGk2MYwmIInmCp9tQcvwJoPO3HEi5qNUhQPaR0BIGLYXNAxC
scKQIwWdUr/tfcbvX3fUn6A9xKDjVFVyqyNTrYmq8XkpctMgkPKqQ93KqosJuO8RRMrUO1v8zcix
AYSWp2J9fQ5IpADvQbqWlKfd9Z4ful2ENT0iM7xtgl4XvKy95u/i3lvnqp4OZguZL9rluYFhlSXh
9QaFEjsVHyEkZAQyqzC31xiz8Nw8p17T8W3hrqfWJjjQwBemwkSdlj/2I+g7o93p4fk59c+vwviE
gPfR54+EPvo3ovB0QinPrbW1U8xI00ZsVdtAgp/cou2HCoqRf5OQyofcNlQ1I4ZXB7V4iQGE+pQD
E6qhMkUF+UIS1hBZTTC+MMPFJJSow383aEfrEdsJ6t3aG25IPqtYjXikcTXGMKXS5ARNOabJNRae
MVfuHoeu8SdgD3clDKj20iAP7ZjKQgnS6n80D41VzFKFReWRZuVEC2eSsJQslDcPPwX2SZBcSjQ+
Xo7867H2bykBmAM6iLxVkoossxwyNJV5ryYGNhrZkOqvx7mxFOn2gD4Cf3mqKhfTo06GQxe/Hrj+
2C5zJge+wT3CX/LpJhKTvzzkqZJLNuxBo5btbDVorVSlhuueq5Q2VhRpM6F/0lO7wz45LLUdkuyi
Bav6cRaVn7qOxKN0xEC/g7pjk7C6G4eiEqaQbtZtWjp3rtnJnFoI/8A27u0PFrBjayqI3m+Mqaka
+Ocie+apm58KOV4wftYZS5vGi1MhUm4GsLGYzoQ8RIa2wtFCibj75s/IigzE/BpS9nQn2w+yT20d
qdcaDua1atnCyHy8Hah6gJ77Ikr/KbTb+y+0fPcilPbEppIdgUzRv+pCbzWVvtuXKeTLw+CN7SGA
IE3KrbA3SD1fGlTbviadwWzp3Vzd2HMhU2iHvAZPUgYu3eoj6sxVTR2BrfZht9e07cU8zisWT4l8
YUcms5j18ZgMSBplpNLIS3mwpHdcnfP6R4PlySrkw0O1HmBfalW2VRcIoKTlEXzqMd25wdmQ8A46
udlOd6iLkwGauGWH8nD83J1IM+hjn2lHkQr/rL9HMOw0jbhDu2jZIDYkueZVek2r/VBUHXYquiJe
Iku8hLHh84xbr0SYSYyoLKkp9gOe2yrp8jo0p7abp36TB5wRadSPcin9viotl756XNP6rpmw4OBA
RwQdvHObgMlBvTKqlTZ6FatShxbywPkzzQtgHTUE9nvQOjkOP4P6riDc9mLh5lE01T1l6d3CWx88
HQfVEQBsy+SVJyofKUrEOQ3rFvHKOShOpPpgeg3XeC/+WjVrIgQaTiD3GhTPnb99g/9p2XejbaYE
7YvtuOJ0XKq/TuoFkA2AUyk1l7XnyjL+F/p1ysmJ10um4RnaOewB9kKmulGqLI4u0zC/5nOLzZBj
DF8xsg93Fq9GuK6V9ifzawlcqCF87IwlMhgFiknxWjmmpIkAUYCxTtBN47qNqchWzNNrBNv7750C
YC5I3quNeJp95ca3Eem5stg6MtQnJX4axb/LwJpIn2Lj3mY2VSVVSBMKgQET93Ea3cYdlgLrbPXT
ZHSIynTuw8EtEsewCiizup4sDM1YfVHsovG5OjqVHtLjAPZBZ8xcJxYWDSWpfGv0Q1VfmggofIuN
uhY/RqFME2rKTl+7IRnAKQ6EpgHSrJIwCfTgQp/k3Fy36dj+U2JX9kHYHk4YM6O2lFaRS1c/v08f
oZNh1V+CAle8kDo0DtGNqpMtRMDcG5eseKW72hrLVu8oIX0x5utDJs7lqEkk67nqmR0z2Vmu0M0c
5z3FuVQrToRKD+k2HXtnvgDARkUymdRMaiQjnAkilD0e54u+nIdOEmtDuimHXJTQ9mAkguo2xqD4
4iEMaTRDjnQkyQv1S86H3PhvdJ5c8MM9ebUgc4TqKjIjXb83QHSdaU0b8deMSBb9nU7paU97vkDH
fqF1GlDrzTTfGGB9e3UEe+L4Q0LLvH/+HQPXqZhh+8pt5SsDrPfEDeYR08dZ9LExBooStUCjA5LX
NtIUSh4fzLLfcBGGDvgQ4tAdJ5Ov1rpFQS+bXNMwzYGg9Qwj+eQNxBR33KMCNOOYooB7Hth6yOJN
FiGDHIKpfCa65B1Mj6D/dbyLaGad2rWvMxg/b+VT1HvAlZd9ddtw/kP440jFK+/S07XbvV5TUsME
LPjjIe6XtT06JGu/HkGNC+I5gzH+v6fTJh+XK729ih0HkTJ/gWy1pJFuQ2X2ECUVr9+HiTzOtiSI
94eZCh6u8gkH5qmmATVObxBE9glH2Lu7Htn6ze5tpaKHE5vuoz//Iu8qTjb3s83NxfeIZ/kBRRsb
LFcKMPg4vWAy4+tRHMjmdE/BkmNnF+wIGUXbYnT/O9d3MjR2YvCg3fbGUb63kdzWlTjc/zduaJxF
pwIu88HekVUluSPV5nvrpdsYcPSlWp1cPbc4lu3CUL7itbykllDOg23NoCjuUrnuSOyKr4xXuLXK
gQlIp6uASQB0wTtET8TT60ZiGogJE3FGGhqGytitKoI5TXKCHlbVYRxHBeB9nu0zrCxehqasPTlA
iyzqBWmr4dhYPA3D9ZtsM3pp3F3jri/ooPksKItCEeseWPMNBN4MraX95E6MKlZXZU61t6gFBzRV
z2lQJRaeRIqlfbDCZAHgMPIk6g/OrcwbYWVW224KRF+Jn7cDacOtfmIUiMF+VbxX+vlTOg7zf1q6
VkNZ/fePJxPTYnAywmMBMcYh8WKE5KrjziJwpOl87FguKMLT9AoTMUeuqvoxH4yoRSGV8m4Vnk/u
C1yUxoa/hK5mqz3QCSkvICTNDL+PLnQ/r2ttLrbDgHSxS00g85X/7D6T2joD2EacxgnZqdSvxo2P
IBUJL0S7rp2F89lvtppnOKLPB6I8kEolSnBcW30n9kwPKAOwAOLGSKN/3e73+CbytEWh8gIN2tGD
tsziHqBtWABLHXAy0gRAvgPWCBHDWDAY0vjBAg58NlGINxuHTM1gb1Vr89YANq9WS1Kq9n5m1JL3
ShKJx/jvfMGrNeteDqC5DV4Kwrn95w3wy4r0ql4ZTa5nJRXDcIh0TP7GvmwA+d5lJZvx6icYsWoI
zBMU3jSsbmoKXos1tipMoV6+HH0dR6mEeLWvQYoDiI/dg6L78AWt/O0IlLJp8Gtgwq8s41jnqkRy
OS1i4OJbkxu4FMXrjc41YVlAyGIMWhA+GR8OWBqAf3EZEwoTNjG3um8mmv75cr4XHyhTBU/80CfI
v8SAwJD5NfqvFHI8PJKyoQu50lp6hb5GcQLgqSxWPTrVnYxdWJxsK7SrucIxF1+icDN1earmqqNP
IX5a1rAsbdPfZ9cs42hL7BV81KkMQv6UFU+4nQuP9Lj1Z3QnSFc1BCyjYd50PmSdHF+d5AmyCsCx
Trs8GNkpD1Y0U14iWGFA6Hk2xp3BFW5d9CidjO9+dNBH5QTtMHTiLw7JOchYnnXVD9OhveUu51cV
GI3HYBP1jrriNEfDccuf/VORsHZB/VJ0xHMn9S7znMse4BfLralwphD45XCZvgMliCfvPfnHNwBR
mSk7PcwP+S/uAvABzU3oQRamKzZfd+nDFSKeHfZus8b0twIzXdQ1RpDvL+awpKS9h7YUY9tk2kbf
x6UlgEv1g57AZ8d+6F1jzWlObu4JmY5IGQjik+gs1TqmeqW+2Bdu4Gw9+XGt3okdC3+rH0zT3NAH
CkbO8o2T11YV2mY4jYzDcIoE/cXdw5PuoXEvZV0J5Y0Fh9trlXlQbGXaeNqvFDsO+sKPKFY+21DX
Xr/xnKWnqZYXOL54eWrldjj7C9PtBv9CI/7iCda7z7zE5tTCXpzDwez/zXl5Uic/Orse2acDYPJx
6drBMoGjJ+KwdXpkzqswH4GlaQ1mjIUNG0rlVyNGvSTGvVSqO/oYsrhEFl3DaFNATpFm4dhNlF4+
ESXL1VHGq875VCCTVKETWqbRTfvuGeLB5sEaymEPT+GuxP+qRic0mOhf0/oXOKNeIw7walqHJUB9
m8tRyzf5w9wMn7KLLmy+pjsixY34oyWx1u0R63knzNUrRJuWMVIvYyHuJtm03SaAKlUblRTkeK2w
RWfkF6noiPPK1/KWfQPEK4ZcANcHyc1r8uZIHfzGsJW6GjXyTXdadTnMz9Wn84hKafJRxSOb02Y5
4hlyCBydOJX11QWchlVI+/fCqtjmwMcb9z5h9fSg+szzpUb/QZ8xTqnOLUwR4DcY+vxPAD75IWoH
qdxtA14kJz3WoDaYMpyXCo1iyV9VjjZj6g1hE/za3DYsPbGJMca7ANunX6qXJXhuvRO/K9dQXvPg
LVHGaDqJSZ/UNKwFtHOZrpsAYjlBR8SIKq5CSJzVXLuvZqZclpiX50iutw/cLWK/LNsYF4eo4PM0
UHbA146STgrAGswTui+QF49Opd6SyOZ60Ra6h9iOEqIvG7/eoikh9/naeZeKswGLMjrnW4MTq0iB
sFDucLbmIT76VoLMkR9Jef/KtoE0UOMuBAWlv6eb9kTedKW19a7TpKyouH1RNWPS46Tsg4SuBjmB
A7oU+PpRomPDG/ANoTG9l2/05msmAJdTBAc1QBvgKO1Ud1CXfQcU2XpavJauRA/bqWXCILWWv9IC
Y4UEeVhBhikQ/aEDI+9m4k7zX2DBgldwmWHffwjxwZWVatu/4gL+h3u0VP0aP2FG8EfO6RPRPQvq
bwCckg5OOxTr6n0ucGiMs03zLglY2BGFG0Xfri7sk+wCUtWZXm2FKEKGGu0nFSllA5XZ5vKfv0/j
Wlt897PkA7oJnAMrogSiXrx2DnjM7ymwMkr+TE4UyIFj4YySaKca8cSFxc1AK6txYUJi3wAXs5rL
DwVzkr/NwgWS8l+lNMRtyRh5XFnisNhp6jCFesaiS07QNDJLR7Pea+zN7Eva55CDMfxkL2FaPnVa
j3aO8O/Yhs57CzODpNlCxnVeTvTX7YEVRjr8F1EBxeMiesQog5bXOvzolHtYbjamMRahUYcpak+e
pcki2flS340lteK+JsrBIVPrt8PTbjEEaAMDMpLXVGce9kuXncEBEnscefiS8XPogNknRe9APq7c
si1y4EyiQXhTcdcV4hsQSJZGLOSAVXIERluiY6ZcLW1JDS+2cTL4wXr7bhcW8pW5kAsbFjhNOWuh
uOIKnlYixJuDJi3Ka1506keZXneROfHysTVmjjjySi47e28hEltVZhJrsNRA2xQNHmIF25XRI0bG
BgJAXc8CT4EkWRc3TtapN/YP9eMkYSOkL+ptraKaM4oaz8wb+erQMIngcxc37sNgZ5Wj7NHnghOD
BvKeiirkhGw5y1TPaECaZtnIR5GilEwoyI1ekdP7zf2XEiXIv1/gjHh7Gdi7r6pJt8dypwpYD7qe
XPzYHPN5EbD3snFtwfZ8xH8qVcGBtxFBh/5J0Tklfr14aqPDZ2QMdYTP9dwa54DzjkbCD1MP4N2R
N3vcYMzxyWJpObArh73ef/vmnJgYSS3w3JXL6gVB6ulFEDJKGQ99yHm9BsGnLKJnYbtzT7aPJcZy
7dY7U/43ikLIb4Kb5R45yv5eXxAH4db1YwTKP13ZeEANF54viG3KHu8jn21oumLBPfqXCIDHSuh8
JSkimKQT0ls4OGXOKMloXCkxrqrgIj/+m+s/h9NxjtWLH5s4Rdcu+sPCIOkH5Wecpa8B3O0IbqIs
9c38K/LbuJhpgBHuptyaz9qRziA7PtU7z0aME2HkvIWUM5Nv79gcCl/3NINI0mSU+8ck8yF9Uaet
P9yGtmIM3Nxbrjr5pbEWgG+Y37exLp2fqOEIVn0QwxW2B8dBRhYvpmrJvGnEdoPC4Y0TQnW5DM4n
XVAtw4rc38hZ2NendzpBnRrt07u1QeAfseOqN6EjzJsVpjgRmLdSXvNKk3ummyX7IB9g6dAdCoFq
MbbCgGuIrvm9cgpUpPUeW2g8rbXHUgbjNDwJk1vDo1m2XxOz1wc0V8hMWmQLV/mabgvmLV13XI+K
TJhTtMUxH4pvfZRJFVoSAOexJaboQlDuN0dZaAumYioGCLY2EZtaLit2fsF549yq2gVkaO/SPu9t
2NXEL+HzcKyp9OE8zZfuZzruWaRvyxeOj5J3WHRpe5dhRgLXhHGQKWQhKTwLSgL1Ehs9iurg+RDC
ueT3r7KDOsvddrL4lNnvwyEcRAtnpPsicuhKMTJ8ZLrAM5PXDJNRBTDkWkQaj6mjMFiRVUk0thox
MHqir1A7QVSaCHvbL3jwC5JZ6MXQKX8cDfckoF4oaF1GAOMAzlQWHeKt+HI0pnSSaM9xC8ktT8I0
MAi6TkA1LoiQjiGvpKKX/sBZujlbVBOChvwg+IGpi2apBC8teZLabPs8jua8o4Qf+IhgIzb7pTIr
adlX1TOZKxs/OCBRTYIAA4JBQ/R7kxkCNT8PxP5UMOTth7zCvyIJrBLmKxobWC1W3hmrLL4+7RgP
UjxEanPwKdDEBGKgFek6Zk49BcLDRGwt6fFrohgeHhhN4EwGZTZFfWC5+RYLPAVeqCGA2mm7a4TG
WAoEEaMjFAq441OTIX3PSXIwVypnE+qV3kgHPz1LSSFhYeFD6Sux5mWFH5zBLHg+LnUgPfizkm7n
HNwo7d5aq1hlu1tSRQp4v6m4iMzYB8FSyKru+bu+cLM87j/YJVPoy9nQhyjPiOuwYicxGVfM70lf
FTaU/QsBo0eg+Y/vAYRZGsBRw2TupJgoHqczDrE7QbCWUzJGHFx7N8/Ja1HNMRAxW8o0j1Bd+66l
k9j8dlaOTRESYUHF/dIGVuHZD1Wj0xLq93E4j1LmxG9XrluYLbtbN/2/FYbXmwvUdpDyvbCKptbS
qxoI9KDHhFwETpBX0undvORpr2IW8/TfmmveouGjHjKCqSXN8nMDMeKviplbsaqyXdNltd4klN+1
Hvx/6iGfDMW/lmZf75XPFiO0Qb+bRiuIxidrjC7M9SxKDNd7AUCwQKpM7ZTx07KqED5JuGLfoMz8
wUFg/6SLLtu2P8LqShRCqFToiVsGp9MtB80J7qWNQArT/b2hxW5S94vc+08VgK1BBZzOILjfIcso
wIv46dQYdfxiB0n9SNhxL0uppn4OjmC/df2R9jrLFQJ8HsvNmoCniaiLlqV960bpS0qbY5yX7/F+
sEnwVfXUAc3GNJJipr1bX55dMv2755AlLelAXanm/L/6eocy4pTyspN0Yl8ObHzvlntex0oW1oyr
GvWuWdptmUyklhJ39NBCdaDp0hXDJfyEPgre29oKDxzPtai+NGwfspxtPBa8FVBoFkScpFITs/aC
nkZ65QwVbWwVtN/doZxbu6JK3ZAuaP9cyjy9vdWudjcPAe9DJ/7w9815c6eEmZsOFzX5perENlha
RMPUN8E0MrRPZ2LafRv4FlIiBGP8PnTENfrns0fzQTsQz5CSLJqRcLBdy1HXkxjWACkYz2iUO5zT
BtxT3HHiZPbwY5eOxyBwa06I2Y/mMkWmQZNdlXJqwRPU60QBsnO0ME3cteu4irGQ638+tdFQ8GVD
Tua45dSlwaWythjVtOhDtJ091lgcjY8DamDNOlNHcvr4rsJ9d0g/XR6EZ1rbjQuHbJYV8dJ/LOGq
tfCc76h7VUNuuLQqd3NHUNbkV4ntOX2114Zs8eFUx07qPp63NrWBf0GRQZ9fPICx5GGSy0r8TllP
cT3BMYOfdZ6ZtZHYuPYe3XYTc9NjqYgo+RoNqsHqNrDTdVsW4qCGAIurBt7UoONm9/8drnp3pdBq
EVslxlbEUDLlmWuTRQAOZKNolE9J3M1X++iG8+AJ4j38lOiYI22M1ooJOuiXI6zsCLtquZI1O9vz
bjpaqfVPsoQJeo3tfzKMUrP9cFZUQYwdDC41nQlPqQO9k00Dk4Y151mrwpAEMokI0WSpYfasj/A9
nyrSJ2vPHzUMC6XSx7k+UahJ4DPKYLirbJ21HFJelTjBmL0H0nGJc0Qlh5WlPnE7DTj+/BSYdA/K
+NDhOFa4/lrliVVkqSolApkUdCyidLlF1OS2iCLct6MpB6PkiDi3kCttGk9yuCMHw4yGeb27ePnR
6xHUa709YKHmDtpm3HLNcOkCTVvhnPIE2KAYhD4tC+YFQrNLFeWFJ6VXQIY72mXtZIQ8sMRFSUM5
SVXT8WGvAj+SfVNqTr1md3MUurzzgye9eoRbUXvEQID+i34TDB7lN4eBOhMyGXS4oGQss9qP7G9g
RP3ndMbLk8gzavzACcBDQ405EbFECXab6xIf0pdJz33sHSZJ1yR9feOCW78Hp+nnScYVDTuVLnAC
9vuojiNUJxVQ/Fx6suVdy7BaXsOUHLnB7kVyBd5rqFs8r0melZVtTO3yFBFu+q6k40BVonsJvzKd
jZqBFiC32Oibp0+Xl0NFXYIzF29MskCOn97im5w9c0STm+Jlhz6MlRym0Wj/+0OA6bpFzp9tnLwZ
34El7N6twf/mlasJfs0DRERnTCbz/rsuxDwCEQmQa6mAuJzktOV0wEjLYZ7H1XoIfvy09aJiyPQY
mp+TkCXBTE2TGM3qU9WtTB+5n0WIk++uk72RZJQPhxiUd22VqKYe0VdqJthuwOQhYSC4w40ZIxrH
OTvlLoHoVHvkQ45dXNRmepg4c2k5eo93iySzFw/EGRmiDjx0dw0dklJOY9BYnjWCoyOC7yfJSQgO
On0mMiHaZLi9Ylxkk0Lp5ZYPUMXvnzLX9EorR+ILtrafrIR7ZRfLj5ykGsIw/iRb9+RnlUETLCn2
WkywEqRF8gymg6ucU2423O0xLidHA+4wABna4yfBFBsCt2MHhHj0L1ctxxAUeL1uOxC0apPvamgM
ctFlhSwUzgZC9/WQq/u4ZxvBZ8SoD5O83XfwxklfllnU6cKeqSf8z5+3HT2mT6rlW8SMKvss5ur/
0uEDDRtNxymb13acKt+3i8Eguq2iyQAxT8pOJG1sapAxSxp6G7m0Cx3zpDBHlUZSHJHi2FOUR623
NRCIgwxlCh0t8YqwrTwRUn6qyu+xOqdwpUsVxTyDPVbL5d2mLu8EuqcQ3P+6p2aljzD0z+3Dsl40
4dJw8OGyIIvIHKFt51gYqyqK0FLAPDoVPxRRKBuTt97HTHnI+KPYacI2rwrSm47GDLavP4NQxVBQ
9kybNluwGI8SUGxCesV9emQA0K2H7tgRD4/HvMhCeBfJ3g8vT3ttlCmWzRo+kGlaYLKUAyTtMOol
CnlzJ/5VKkjdLBSUuGJBwtrDPcmKiHmusdF0FD8tB/QYjo3vHW8QLsbwIiNN8i8QqwsWPxvoKSfD
vb86m9zzAhfUgct+l54PcvsNUMJZq2dtY7QjUPoNmPYkRI3DRdKyQxmswePd7qc9azePfNz5ZEGy
eZ3YTxzE+2mc3lXIc8ZoFHotrqb6BkQPv0ea4YrqqILiNFawlbg7d7QYdbNmCGIqaygBSq4XIfjY
qBAOM6q14uye4inR2dcIJORvMLBww4KZUpFWCwZwlkJ/zbPUIhOC55+9I9G0BbX0Qd7SFRELlxI/
Nmo+kYjDuvRIkHP2jQBobgsb/6GMTzOscYJSz9mcNIqWe51onOP18R/wc2aS0Ro8Grfok54dyJWe
VddVrj8OojcXroWb3ipk4nMR2U6C2I1rUN2XHhQImEMZDckPflOLwHDdPca0lex/acSXMhwR7FQV
2PYBmmZaIC+pBKVu1BvHQNj6ZKPh8sw30RUsiU5D50OhVP0jDUBg+MTk37UJmT8RjdlSK6xrcIZu
aW9RpZ4lXayHCp3PLP9946JrNkemq/4WtZzJ00wEXmBLi7j3j/K1Bi7GNx4zFapghI0NIevOiDmY
mfaT15edBIEIe9ZKTT/exjeran00EEP1jmyAsW/A/Xn0atjUbgencG8OYeDnUaRk6ysv3Re+BM4K
S5ZROullQHdLFYMnoWQr8cSGVp4lQgV1D2m2ZGmC0H1lhXNUNrdLHzzmFJLysAx6yHoB+VQH/Qwd
2dS9MEgQGbQB6d44l5qNgNV/Q5cJsYxAif5sx+liO9rFn/RD/nxm0xh44QQYQUZSaemAk8W4Rnox
rkzAxSKKcIRJgUyXe2FGNsq8+RXJPV6Bb7vQabGwRJPCS1DV88R/+pyvNgnX1wj1z5+migfyl0lm
LfqEnE0L2A8KlixTkYPIrCA78TANclQYfmAr94+zq+pp/WGkI68x3UCNPSIfaBJTWabV/73d1Zck
DNd5psBgyv8dYCho5l0NVzCzZa4425eWCEWX3G5PHMfQf/Ia3+8zgXhfFRtbCP+/LkoiK2cCjLTx
g5hYDZEUnmiQpx6uh4yeNesuON/wnlYbEK4rblJZpBazqRwTRYxE7Udm7N4FUXotiYtYsAeICZqQ
DG9wM3uvODXIdqadJ9GpEuHBYGYXq9HPQcEZiCkJ6iqwYWUOh1ZqbhhEjTheafguaJS3qtRCb55I
iK8H5uJQxqJfNUTHyLqUTqmNArkXUt+DigC4Ek31GnGQAFfMAaZyziyOpnYpWtFaRg/1y9Qew+2q
P3wgQyhhVZE/E+iabfPqkla07LmY7N9qcbBBMAe0sANZPl2I8vmwoK2VvqLvTLZabCMTEnTuhh19
rsdT+6ipPQeUPZHqxYgt8HwN4hduvnvbbJzoIAY1tze6Zdoyd5qL6fFBiQ9ynMHYfG7eQYEMR4TX
NFIgDnDrMS8nv2TrFkmk4onsc8byiqBIppkWhK85J6XaO7uFJXE6r4Vyp4tKFO5gXnIkYVkSJyMj
mdPi7f/4RTmNMPttSYY+Y7jx8q7UAVr7QT2r/htOaVhQKiG1zE4VWLToYej6T7oeTSPUvi7VZWYU
e6+ZgrCQDYZw06/Oc2xuqkDOoQZ8b6BpuWa/UCnM1AFynpJrzL3o5PkhPau1Q0tw5xF7sQSfp+ar
SiKU+DJgcg6ODY0YIfRmZYny1p7aHh9bqHZiXlEds59sgU5oW4OlKPmb+OLuIGKDr+ATSYHufvcv
+es2MMjEKJ3IdGvyq3swOM8evwqCHPQuPzuzcoepvCJJqoEK4hwglomKI+mLMXy+emLTUM0wnekF
R9gOKt8M9NxPegNFCVRSLnNub+8+KQBarDsZ5u5DhDkw0Yx7J9o9BVH33YeBZjHzJqE4qRP4PrUm
is1IhOUb8sy+ESuLcrPBk10DGQsuh9jQmkxK59RUl+s/m0c8vG3esgLfzg8yrjIg0JQ4Rqk3m42J
lVLTbXdZNLWG7ucV3hoviUJAbvYtHXlct7ueQjLOl5wW855W8aFYwP9cN3u0H2YjbhaltsHakKZ7
UNPFkCnZjVJrCB1Zs8emUq5e2rwhprtPrqwXlVcQpiR5I6FTGP5qyR/ARx2Oo1Ock+AhbFbSwAu0
StIIycJsjz1CfuSUHU1KbNA770EfgsFPd1/O4DZXPh5LlXpSG617PEV911PYsdLPGdH48GluBMPN
uLOUmsMxe2X1nkyYzqKxzdh71bqrDVg4TiZRARLu7RdHK3pqfc1REvdu3vOTV0GXK/1EZvfeejyf
CzW+YTTIlezuyScKvEYIzd/vdK10NqOkbjF8VymX3CUyNSUYL3TT7xa23TGcwD9g51UShrCXXXJX
fDs/M7Rts1l0d8mawBTGGRNx4+pqpf0rc30b1u7UCz/g8qkGCPIPWK4TgAewZ8DVWrFQo7C5FDHe
OntdVgtpecLgCk0Y/n0ouDx396UH11PRqvtsZXbiPVv9GzwL7Dv5Ap8D/y+aTFtYKoIbhLT4+kzA
DRYgBdCYcGzOBiKZb8yuIqEKhAPdKr/KJphQEsxiE1MmGgUWjjtmE8LW04FOvDFVkdr3oh42UvPp
M+IMLYl7ELT7h2MfY9XHU62eCLROfzPYtf1q15KhJ7X6O453hKEVsyCLMhMTQ4ZdFCgPzYgQ4tuD
ygeGNbwUMBuwhhrlp/yzAQbLQg2FDAhBGLlP3d55NUiObnV2k689DXJjdefkyVGNfgU2biGH1mr0
LSfP3mjYBZmXvxJA4/8FkZZj/8RJmxKwXX23Vb6WQ7xBqKWe3CdX5474NJ30KBTXBOLc57MBHDQA
dr20K8GuB24L8UWKSsA+/aKFtN+wIMWeKr0D1BDSJLVSTpgDy/lCQ03SUPHvOquZHO4ucAgEH1p/
iDJgOhML7NfDJ43ngKhDeb1aT6ocRgr34PIi11MJDLVfPuMA/oqF79C52PtDWpzQgZdjq76U0AaB
PjalZTdaXVryu0mtpcYMoi259OAva4RWCKxfDmmughGRaTTNSD0Dl2qoqARJYtLrJ84kdGrH8KjO
UaFhTeYcnahPd4A2OvWyl4UK+yNMxojInNrwnBDHPz7qt4ApKYpRNGPtGHxHUTNmiVhGi2WXo7Sp
SQDgeM88dRmsGudISk89jdWIzKIyNVy2rmg+OZ0ffNBSFSs4WQTpSITML9I7d/RKuDIJ/CevNHPC
ncG5lWjAPZ+dX0pDQMoYlOynvhIeqaE1JXdpErd2zR3jkLHqFNT8eZK5SUE6jE43pVhsF5PiDHNu
Yrn2Q9gG/n/Xk8ojUCg52ptYdGQ7mjNph4Q+OJa1e9h5bGELtc7plnHyj2NxcfKzS+c2s3jQ38s3
XtAsCB2ghpRujtZRl3VgUc5wyXvhr+awBzqJT3VJDkjb/5W/yoAsmXMu0c/PI6Rtn8znsgqA5euv
BYBVESqlNXBql+PDKJr+1As+zbWFkMtrMYm2g9+VvTLnRqKXx525EqjUpO9kMM4uNAnOKlHWb5AS
kprsd1AhTQpKQ+a67qCj9r21qKwXWGViD8pekp0QxYI39BaS4As60Vjfkp3v251TtU7qDw838myH
U0HkAi1vIZBYRmtYXyi+OuSEP+o3N1RMMyZPniM+7DbjD1rKsTN7oorx7iY24y3mZKF0NPoJH3zp
uvdt42QZTvG25Ah77M/kAIvlP4RqeuKWsirUZnhtwooj+gYZUe1swspzGQUVh3BOu+B3uwa6JAsY
HLrUgcJoBhfx8LwfC1X9g61dKrnfLhCG1fmm6Anm412KKAVGZffsW9mRcRVTrFyY0ZgwSmVN8IrL
qxb3XRUMQCELMd1kyVI2IDlJ1DsOAhOKvlGrmBywvBzZXKGRnWK/ey0FyqhDzYsmU/OcBNq7Y546
JHttr1C0l3acOi1vfXs+fFX69qkMTrpbXT9ZfsJDj96vaR3/fSXx1cAFMR4AZBeRB7OGLtA7j99H
KQrnbo2eEntPfIGs78YcnpMS8UkqtSFUiqBPekDZzFQKmK+No5pOyrLIzcon0L3AE8Uhh4TBidvV
J1RkvjSVeZhQTMDdSNV5/hBgiA2WlBkSgUz0BlMs4Q6gBEsfsbjb9O0KB/gUTTcqXSi/RrN1JqV+
6o5cUTZgOUmXVHWt9cY0P8OhpXEyRNP7m8oigs1c7E359si1weBPi9OkbKQCZ1uGTb0lVnekHT3O
5L8WGuzeaI6RBuynEReq8ZIujcTX8vM0HT05tKH7l1CFH7NHmsfue7Nhsclegbi+bDmc7YsyPC6/
ky8tDJ+w+rVHDH+4Dlfxt5UMcapa0oF8QVnfigk7tPC6ZCgavPMIUk6ZxI2jpBmEOQblJQ6rAPpy
sV6b4h+zSL2pNcCoPcPfEAB6DTJf0hO9zlQ+vl0uZ+enIopPQgYUWXXFbxWU3tfGFLI8lHJ5OvT4
gh4hQQGQGCG8avxDqflS3BFbiU1F+B8DTUYB48f+XYihELq3mAXCrlJfHHLmfA4tZ80AKHEIuxkZ
hdx0o1I9GF5hREJ7pzVfRInsqLvoyqsjHAzOwOsGhdCJoFC5GjfA8CtygU467cFxgYqxgoQKnXfo
0LXX+t0TZig118Ty70bzqGSYkvKypp3Zj8ll9WVih/PEqCQZ4EbUcPHpzu6Xu6RXoDg9uAnlKSVX
9dPvSu/QgsuqodP9qA0lMwtuYPUzWksUt9KAjRaXEfMCR7nBQt6K63VrezBMmWMWTQYPepiw1A25
QZvmPl5VTP4+jCxfcpjLW/QsQvg6ixzWUXEGDle7TJh/kiMFKEHNlPdyRCPvy+1l0j33y3GtIyv8
Qu34RVNqaBoZLhyinu2yLvUJ3xtMPb1hwAcRLXgduUXCadZ1B79jkmAunsq6skFoFzlWxSUasQtD
ZUwwgZFFjND95MTsX+Hx3++BQoKYivhLmFBGqe8uzN4rreLU8nRpH5IFX1vbBUPQhxxeRBNVhWv/
EPsSluc+1MLzzN+vYstv6hW2NNENy2oBclW0fBso/DZ8BEEebEZTCtXv/x3zibJUy9B5PlG+13ZP
jO8uzjy6v9OfOGBg7mWi/LAcLghFGEFCOu/fZjlDp5pbE8LWWc1pGIM0Il0CKJ9cqyrmVn6bWitf
wFI++oxJu0yZZaz9CysRYupOrNb/F/oBfKfpPYahq1p0yqWHBweY4/U9LSqP2Dq/YiH6g3rcMUHU
GLDV1rplBagOM2SctxqD5bEWOFEi9sJoBOb7gcWgNgZ8I7dbbLmKwMy36IgmkfJXiwmaV/XANGV2
aObfXyAYC/GVIosE/FnrCP9ZE9tm3DHLbN8QailFyevzANYKSNFPNMHNK3OxnWzJ+BMfNrqNYqLs
c0Q8a3XHeql0zrEk7oOAb9Qlb5pSuMnsahSPlgwbEJcy/a5VPUiLizGImGVYcurNPRarc649Dc8K
3avg9Xq/Vqq0SNyswdLtIHaNuiLwoSPvu5THli8FjgpoeD1tsyRuxPLNFh5Sr1bMT+lcXpQnRurG
XPBlNmBO828mzFV7439S3AZsbpizvAehBtj5O0c4Y9t8dSx5IbeSjBQpPozk+H1EeALXL2DbuXYj
em+rNV7Zkj/VY4WCuiqDj6T7MRSZtQsvyiRvTj7xHXGqY3VjOq644Ez5Fc8CTx/g3XL2ldhS5kne
wJhOeG+H6VRHQme2IQ/nmMCBs7d9JnlSZIjtrpk7afS+6ogU8P0Z3llnjSxH9eQISyHNayVJCeUh
+r2mnaOmYwUqDIIHMlL2BanheHF+xMBL5k8euooSl4KVm9iFmykSKOF6GXzNbB3QcLENKwmkmfZY
cZZSLs6zHG8lyu2SSXHghXjkxbeZeMBBpc2V2h8cKt/3Az33MQ70XE4mOZMkdbO1tCMFsAtKOEsZ
2rr7W2mp4QSIDKQr/ZeRV1P/4xtEiPE6wQpWikbHF6N0/DYSSa81UhUXObbTLi4rJ5yf6evHssB4
9GvvqFfrmSLxhgY+G0T8rU1cA5yeJqZIykjg0SIsD7vs/+OgafghX7XO/gtXzFh8NVJtHrpRSTgL
cVQgT0qOo5J41o+9GF9rD6PWkT+wFU+fnTiKKnFauazLdZ3bl25CmBPog8XTrRx/37LOnJwVTo0M
36k+arPOpzvZjFAG3dzyIdvTirpWWgm+vl9l5FD+Q6Sq2MlA9IwDJfAwa5sMlTmWbmWLxCsIBFuS
WdKJfZSgfR4nOF2kQBhDWsS1o8VXPuFrhuAUkplCtAR23KSBHNoQ+OlMdC3R7VsZHFX0D+rPe+LL
k0JySps43j7uqVgFt+M1Q2N69WCx35INhQNys+xK/0xblyhuWDN92wOazPp0xu5jH6p1ojee9vpi
bfpwkJ4LLbduL9aE+7wVoCNoRCi0I+4wH/Gn6v8qFuPvyJ1lGBJfD3xm9AuWRoy9Aq28PzZPejhH
kEwpGMvnLKrbmsidJDnP5bwtD/Ttx9pZttOk3wg05BsS2GRJxYED9J12WOL0ZbVoKbVbLXb9dKjK
D+5j1D7lyQh+luFBMGTzlk8hn0TEZtPXWQjMNp3XyZvzR/sqqxAltlgdW/kHQifOmfUNDmhe0cYc
tQG6lzknQTC8I1WGjJZAzqLkO2wnEiZVfamU8vYG3ZuK7QwiFkW0BiTPinCfhEYWNGkTzh87Zby/
DRbsNq3gdaecxe0kU3DkxoD+mb0l10iPlgCgbYWMLY5axSw81wusGgtE9c6rkZsPTFsbn2tCRpxg
QbbAsS6TscCw5uNpNLfe7boBabCIsAgK3jgy89D7+mLmgAemxFq/xeAHOg/7tF7FJnBQBSYRsKu8
qSW9plBodKh1OdZ8AmOMd339wGoccpU49mMFqQStijHWbGc8geuORoEuYeztNvNUSl9ETfbGQ4Ek
1eMt9oWci6YNk1dIV0EoEiJdHi3fGXvfxinSqxvHq+Av5tBhoNN01PFiNVcJraXYCVPE1bQ9N+Rl
/CAx/kTZ0mh4WZVHjfZR5QrMN1fP44YlkqFCoRgCdLKPtL01oMd/iAgC7j54NI5Gk3fI+pyH3a18
A6NxKee7e+C53P7kbqCvZI4aN6+eVRzaG5dLjN6OSIXRbRpGtZHPhMry/huZ6O9H0aipVhSnA2qG
OjsnqoGOmykcyWbBcVhVXUIwxhkDOGxS6xf2Xn4hBHmC3Uuk0Ttr3QahMjyu1n+L2P9uHHNl30Ea
XQTQTpB5osbrTkv/ri16ZUhWtMZac2szYmEO6Q6xrh4xMiXBY0XP0sVSd9TMbDUlrQ6/ZrUsg6my
Lw69y2HncAnZjMLIQyCXJIG3mZEZ2l0PZ92WJCgtbhMFYWM2TaKVXHNGgvvz7cSrtr9aouoJTy8r
LWQK0keEXDQbAkVlMM0isemOU+3oIVhC0uSoFWALnaDe+M4Yo9JmWLi9xp6Br0w8YO0lFGTCKi4/
hluFCOIplvwqZphpHTvC1jQTpMY2eFb+Nk3xpLiWj+JfFghT6qaH1MyPBaAr7NnxBZBNSDz0jvLX
fTkkTlpwglfXuD8IN94D1PUotRkzunmXjfr7NDhYpGkcfX+7+3zt1lnY/90yBXtOl2C7xrUQ1eh8
6YT3+necYRc6lFwW7CL0cUXxP0SCaTAaH4bwkosu3zKjr0PS/SS1ECWig25+mPp6Y/K0i8aKTNq9
sSwLIP/apU9FN2YqT9Q7Qm/7xxz8AXcXadXIS/tzp1pRdWg6ExDnv2KDDR066aUzV4m24SKPpOJN
fplvnulW2+mBVR8yxQKU426j7QwiKz/yN3PWS8ukWvTfuJa+8e1cnX0iMEv6ZWlppH8+LgX2Foty
70hRku+N5q+mhYzHNmH54WRFTUBAj8BwgM+rCYvkyeQL4tCNHrHgV6fMqFh1v1FiBTqoMytTvbg0
0oPaSlRlfmqoX3ZgvlrFvlkGnHaXmCFOnoPEH8ftVUcyZx6TEmUsctbNol7k3ztcGkjQlUbx1kE4
28UNTyJ177NpUhSCt9JwLP15tXU2RN7C7aZp4OqKWWrx1C9tFMxBi3PWrglk19TbHCyoH2tUCFbA
xbIOUd2yjVPL1L34HeV3Z8Cd+KTHZ5jaJbqYH9koWrnuDAt1aiFGHDpEK4ygOYHp1vu21v++mSwx
DoOeP0iQ13hdtkdBD16JaHHjByEWNQqn9tIYJbEogAM/9h3tF6JLwDfNlxKbCtj+vlop809Fi84V
rLlI29nJcwEN5qbRMV8U+d/A1vW8oE2WP51BaHYSriS7tD5wpsyOEPV2MrGz+KOTLIKCpg3feBrd
9XoiYdGUItqnrGtsXUh0fjuXNxnvvbIH5DZYC5fcvfnrKB8lk/U+7X3g7tFA+S4ws1rTYIuDXPzi
QJbPaHo3G+2vcCfgA8QQj03xsV9HI9y0/q1IkemIsEbLPCPvEP2oua17CsLHiB8AyzCqtRb3JRNI
4O54Q+rtu6v6q9CBqZXQBdk2RcqHhuaz9BeqdjEsCxn34qCuBf5woTbMjJPbaL9XPpXzNaVOcP6C
oJgFBCK3FwyBM6TbNrSzt/VVKG7K4cy1B+g1y9uXJWg0wEQg+9j1ilB9Et9vOgWuPMAtyDEYjPNT
9rJmPTBP+o1nM2rNOKPS7Ue0vXSgbMoBCl4LKkKtaG8MJwAJqUZfFAwSv9vUB3szs1QTKeyze1op
bkUOloCii9W8iQ7a4iLmi/4T5z4WUU3Hpfq6q0Nvb0Lx4hYX6I22ovBubaSbYNPC25y2MU24ykz+
f8dRsykGU10iwTKIGTVY5c98SPZ9axz6bcPP7MzecaQlWaY5xPDuIV3NUk+nKmS8fOO/IRy4GtJv
RSxJAJMu603v4VoyQOmJDToe05vQtEmyz7NnRV/5ZS4M0fQc20kvOlfKOnSaw8efp8O9X0G8nB+P
gv9dxat3Da6PNOk6OJrMLW12NAt4zyVDg3yQb85ymDTb80lu1Tnz5NA9AL4pX8vLgToPcBkvW5a4
Cf9M943NCF6rfyNM1GSAeLua+RqyKAVK9MlM1I0RqNNUEvY0h6KR4GChm5heU7d0ZTeel4RHcA5O
Cz+/qDNKaRFpe84G57pT/lW4vARMVrFfn27KV2ftqBbPOw6VW6eSJ/ulBH+tMiKF+iFzEeT0aO31
KTxDKQgb7wDPWX4M/ErbWCQwSou5WmbCZRgb5tftf9yamS+G2pUODhjiSsWw8b4pqsjk2oZcDjJ+
ZhuJ9xqCjhcCu9WYaijQdaQ3Qt5tGXlhpNktsBqWOtqZi+BNeDHdBkRF8QklUIRC7snNy+0LZySz
8UmXsbGrPDnCMEF9Ge0X0F+PfZ5SbiD3McFz0D6Shq+QgUhxIg0662+TXR0lFPGXQymlJT7J2mtd
BtozAKkEPDV0SdB0yBPtqnwS9DR763HD/v0WqA60J+OtWZuZkz0X4mzr3JdWbTm06twVt5AOh65M
J6yubormyp0oK9Pb5/Hx+DHcXCu2LmaToEO7m5R4hYYeAp32MXF/7q7ItbQQfZgs2fqJFmPzlevo
ywLxAa1cHQtbLz2gU/gjTGjNld97CUwQDRtfbfF2qfM6B8z2DkQ0ffUQ3AYKzCSj1/x5KZQ4H5Gu
rluWspEFYvxferGQ6oesDVgbTcPaPgE9TdcQp5RNJ7MZQKL3d3b2c4nmShLU6WuNNSdD1YLXJCvv
iFNdOXXJUHj3dmP7VGx1EI+d7ZD1t2Bmu8yDyCRafnj/BBJ2AC6oqzXeZQklygKoBSFGkXQndsjL
1Epd21csTIpA8nTBIZhhuc2YCOrzN650VEtQaO7vr5O8yvBM09lO0HD3a77ZmPwmG+gCwyMHizOq
3qsC5Hi12grQYoU1sQvVVOb5uAy51401keiJIGnK6R8AAPBpmn278LJsBGjY54/Z5zodSAR/FgBK
XMhuLt0BMTQig0s4RyA63lit1NR7OVsRlMdrNa8o84kILlWsikQFovVatBS0Cw7hFBodvZUlRh2F
qwDTMPj1h+KUany4iljKdkKhqT/7TJ4UrLCGuYAUvA9w24vZgnhGEDt8RzR2DTwc5iHfYgY5ueg2
C/aaWf1GYgYW3qMbRMg9Fh4F24uDM4iHe2/R6ObqNEj2tW5/ipI9QoN7dsv6vk5pwt2wOQA3KBrh
KYLLt8tuW/lPV1ByejmwZtSLh8T8kTZuXX/P7hStoVU04hDIIFi3Hn/ACngtZNLuLL80BJnhFEko
QR+iLusVqY4mLF2UgeDHdbcwluZhwBqIJ0bM5uhbo+SA2JEEQeyKvGoq9nKLVl5H9Cv+CfC4eZxK
kw3mbDETubBb9zhe2DpX7nmPWAUhDw+eMV2MQAPd5SG5150U9+7H4UJyMAiq5aW/xBak24qlQ4w7
5vmWv+q6kGXxIDPKkRd9oYdIH5HagYrtWAHqcfYVdEbP20c0Mt0/coc+qke+UBeRx1CcPvIoo4tM
cuL0zL+p/qzvzyAkkkXrXZQFnS1IrY/zJRZ3sOvKDsnOfxQ3R6FHsPp8q6hweCJ0EgSFW1/kARO6
8qJ8uvUa3KBNEKrrkfKkxR3GYI2gz9DNwfRDwm4OfqpTN2FleWW3pNmtMs/9zVtFLAh7ebYZf8ic
gAOLSrVsTMFkICrYuS59xq5ZHIghugVQVJUZzwxKJTa2SpY6i7sfh/NoexZ7r3E0YAWr7Htct+PR
JU+qvG4sc50vgTRbu63j8yKLeUFJRpbdQuJiTkoRNqNU3jEpvgHeq919T3Ch9qbHGGGrTc+kaRIO
8e2lsISpe64W6e3izgG2A2OcPQjBVYL1hpmTt0SkCDoySO7pcSE2FfwZwjkb/Z3L5Ah2n6zWUcP+
aMutzYEHrJjbm49XqKNDzfrZns1d+Bczyvrv+BQefmlIssHYwIgm5Qgu5FCw0eDDi7lN7mUYsVrN
wseegGZdTYaFEATSETdTPkn6sr5DxeJgYYlITuZZ4nyN/8C/RZXRZVlx5MLHuMLChXnKKNmb8qhD
j03sgvz+nrH1Uo2X6q8qWQcRKfU/i/HRoHl9/dVyXlybxFR40PnEencylQqeMrRFYuJjhTGdIbFR
re02c1mrgIO9sQb4deKiTeNY9SDwbaeuNwCPTN987eL13ix2ma6pAwvoEkeCbtymimD5nBNiT2oe
zGvDAiqgI/9MqOEcxiA1NMQdAsujKa5nm4J7bfZ/ngUk6V4a9HKk776yubnxhDj/JhDU1VAu3Fy1
wQRocKTzT2Otl6Nv92T/MVjLIJDT6jkd/mwnPQdmvs4tmPE7F9qCWoQpmnfggHB6tgDSJo4c1bP9
9NTIujIibDr/wZAt/yC43GCFgYE972oZRu2tCKBYf12V7ZRiuoGei7ZOfsSH7UnBrIsN1H2h2z+f
oyPT1fDQtjNWrDAwsGl4eG3dAfM5uLoQh/D1TL0FeQkDNR096PEoyJiLdY+xPH3IkXB8GFJPd/9J
3YP593s+xVSVTkFb1lVImsWGVvfbsHL/jX6RMG7sOgfNPhEAIPEF5ZZK3wjtEypjBIjG1gFfy5nY
WEH2JIAlk8Xdqk5gkbF1usWZYrd+DoUPs5hg5HDKJeAI8Kg3HbR3Q9JpUariWq9qKhrYHwYIYW0Q
hOiLhmPEE++8TzcKjk/DqHblI4a92HFEt9IfzdWwl9y4atUyuWp1P986ECBRaTAPhAMsbEncMYXV
XmG7IMGn//gE85ENF98OKH/t7eCTHOrcJr+weUKSqV0ian/02bPih0cMIOcOCheRmZ0UEeW285jF
KyVx66oSAZcBxIHwJdzs1kGj3OSRvCzQQekLg863gW2IIU1WQdV+1WsNXvyzVhoMRAqp7tro0OYd
2ICjbx3zgeGvlKP49HK3Lh4cpPBJ0neQx+clk76jD46ulxlD4/mdVo+ysiJ920K8Em29eUhuGpZZ
YSE+pC5VIF0+CGdzQy+RN7fimQR4UtemL+wohjpVsOgdNNfAI/ssEtLomoUhe4FIaXv8ICAV7cky
5DN2jyJ42UQJrjSVzXjrEUw4ZuzZMbo+nOMoXeqedI7YelCk+byR+iLRlAo2a/bXybwvomLXZLvl
ctCURWfcogPG+utAtel48O2OnO0waUhoFVAfI9AivpNbMKhCzv3JdGp0hzRr9czVUOhm/m1ojM9V
jbG3QHE3FF58LlFrcC5l1cVrEFYZ9PA5iUGh7Y70JZNU3emsndGv8bIKEx9AQOg8PpHX1Wu5+r0K
POW8fEp4xBfw3wfiPt1088POdZRPcN4hJ4nnK75oZHV1ebyOXQ6JSdTrGMBEN4dqmbuZhys8YU2R
IHp/x/T1/8jk4Vy4jS/6tYsZgNSIUoFNSH+osyiwXSRIEnziP86u4FUzGu7Y/d9QYee0oo+Y542L
uNxFxqJzxInrf3gEAfT+6pnduC7BwWWCKAVceK8HXlMs9t7nT/beQlYDa47eYyGxuAQwYnLzN+ec
UKZ1wqS+NyK3rMlEqsnEkhns2RRH2N5rbdZ/KrjYxxa1DUnFecLI3C5kX+5vFNxbdkos4woCa65j
N+qraoBrWOPjwCpTzoeZtWRR5+/zzgbVQVV1zrgg41zYE+p+/m3PfsipggXyyHfErhhgEKQiSW30
ra0STSj+bxvZRxwMzwSlXM54jjPfoDt8NvBgojEQbumrLsQtSafVlrRR7wsV3R/reMZEzAEbqyBY
a7NxQCsuSpxlAANsiOO9PuK6dK52Bs3SNk5qBdjNOa1n/937tBvLMXAEjznvHgV3zOGduW+mKAx7
b5TqjIQF0vyg4JSsKixid0rXkTNEIyW6VtvNJi+9TP3A9EQYJQjcqf6jzRIUw5DDn3R6UZy308ou
y8i3F9Cz5AErPM27lDKJpc0uDEFljVrTpUO5GXkpSc4h11V2LBQBMxElwACJ7ix62gHMhICwFAaT
UdJbLPkZ3sRjEtb6T2G0gGkq6WU3UgiiMFmH24y8iEulwvk/4Esx8OH8uxQRn/KbXipKJX0b5tGe
VqbPbn4n3unuq/PRA6KCi9ja35O/hzIzlI/9whOndzhuaE7OqOgcxjojAPzYHkqqV71n2l2UWzh0
HB2kXXsdubppy88oT9QCXRqcEUrsOUe52a7TUgAFnDwrAbGzi2KVxzIRnoddDfd3+heEu09zcfWw
MFfzyxG5NDTkMmnV7+hvqAgm7WT9X5R/qGu8FKvvno8CUKDPisVIKugLaS59Q1Mj2VF0XsuKV57a
mA5xG7/oNaLR7Ak8hJYPDFJ8F3H9FFrlOV8Jykwh03+UuD4338enhw+BE3Cg0w5EBFWSSGJUTm6O
QV3ap/u3YAsn27HTXczNHLP8Eg+oFkCUkZz/8PLvZ8Ar2kXL190wB3FUL/IfSfzjQGMpe245m9vj
SJgF+dReO+5cb51Q7KXoWq63LieInfc/5XsUZo1P7qUtsdMZskLQWQutFhcD+1T4MtZrVWpIkvOl
YiDyFlyQkkfFTsljLANFrMXEkhoXlGo2HsfDsG7v2ilAMdN61mIIopSXLbPYVWPC+HFOEmHbNzHb
nLqr00ohqcvL33VWrtmsJ2MW3Tsq0+anPE7MNwgFu+ZKwkIo/IvdKb2bN8p6dZeiyUcMYa/0lWPc
EzsQnrDJkZy3URAV37xyp7J4rMkx1/iqejxH7JdoMdw3xR5Os286dXRBkc0ICBQFgE0XWfVEm/Lh
4TLorOy01o5VGg6wfdueJ/PWt4MjJMvnd9DGBxp3KyCp7Aj/lAJKhSdr7N8ByEDiHcxsyh66kMVd
gUIMfB9c6tkNwGrOAOz2WE4nyenlzyWv7E5qAHhm9lAiat/C873R0XnD+81t+uFybVGrN4GYS1KN
W0hp9I8Rep/g4OhiRR2DVqNOZFwYTuUuYkxGhP9GQT22a3jG2soaK4zDOZ9bz3kyR+Zk8vk5slMw
Xu3SFvxacvsvt8DV5dtzGNhTTDPYKciSJUC06oWHHlXfpKMM9ecHCsneCWvJV5QUzITyg3T4q4Fd
K6KdVAYZn607xXykxMxod9AmdXjoTfdOPLzD7QSv1nyfCKwtE8yKqJkoESvXAIW+pMQ0TFhINguk
14bsQWmzJy6dvExVD7poS77WIPKY+rP9YHohb8FfX2igWT6zj03lt2wBq25TlMFIXaJ6kGJLHB9v
87eXrWEl5rlbNO5Ybgp/MDiXyzG0VkNntgPPiKIEHFAFyr/ekI9WSr9aVznWVC6IFiHhGovVE2bg
5wm/jTY4ncmFbysW6E/grbG24zh9is4lfNcDH6+TJFCGuykWrHjsFy6DhlN038QjoGGyaAEFIL5u
/0qJI0oeGlfRSsTJpSQoNla3r37HCcm47REJEcADpMvMKWGuqPRWMxyvenw8pVsnw8hgD7+i+uuc
SHwnmsM4AMShpBNaeYPA9Ld/VYQ2JBu4nxTZlmCwdIcm9dlUO7UifRWrwP+hShJa2yWy/1YB6PZr
COq9kgeHDAFAdM0Dqap+GTYhFx9LK72zN3OSo+BJEyvuzRlOkDMpSS6rMGzTKgUP2M+iU7wWcpCo
9LbNdp1WqWrIkP1qtjOsTQ4krHhOT+enksm2zc6nOZ0m08C7al0A7AYsYWC5r49/FHhnPdfoUJfY
vwhgVeS2aCnVXfl0tvzy8JTdNvHtg7IhvyUgbCFk5T6ZECkfmIVGT8Rm5Jqyi9a2Y8OT4+mb7UMr
rcX/o2T/bJPmmjZSd/gdFXDTOiNMCtDNumHzBu8lb8ouUMO7Qt5Hlh2jGALVHggkY1p4MjVrmlNE
d6unWzNtbXOmvpg1vEglpI3bChplnKq/niX2nH2W184udFhoVH9YRtKSt1MJmWqYIykEZgyx6qfI
VH6TEzUcrZCVQ0vbCXx0QOesj53J0JN8agHfOeh6UJUQIdCzKWkZT6EAetWkhRwRVexwm76jHgU6
OSjMpmpc9RGe9MqJLFFPKlvD4kQI8VpzRrXWhDEJs4DUmRMqwlAUU/81YQK4kftpXsWQ4NWs/Sqi
hBJ/L8tMvmVLVC9szvISU7U6avdZqkMAshbGzKqxCKoT9jpomWAdF3i83FRyfwR39pRVSpEYD60q
Z5JkNmblSlTnXWpFU4lsNLmOdN+jQFx4T0b8LYdcCmhGAgglhKkf8AKWzLS0XwLAwLFs17p6fFwv
kiLHn+4kDninERwodrrvdpMCYVOYZUFPKKlMYVlVOLwhlTfFSmXtlZlSGWoO7RMw6209rEOsqWIW
8WS76csPQkjjTYTkAnk/4D7v/+wpR8bW/1//t8WapTKY9lXu1ozYgUhRh1aRa0tSuE4Pc35lmER3
oU0IOlMY/diqA+j6SuFsFm3muZAgUkpBRO1CzwqPIGu3NJwc8Si6faYrZDq850+uGfqaOr7AnKoo
Dhg70Ke7hJ8HZe6M+eNIxvl+l0RwPC2a661cKr5NTeVN1Sa8D8VCT1P5rND8Cyy2my9UDFg2mC4k
u6PGoZxFd2I0DalW7gYDwZ5vPr9ihjyn7+bUGlJarcPpH9fEP16jtpBXNNbY7i7mY8a7VEBObAiL
4I3C423NAC8vxzlsN+4IwNOrYpHT4QLVWyN6gX0DYfpVtfd0Vw/BxJSYEb1AJiuL+pTgGOwhufwx
MvzBP2pTEfNMk2beAk4GltGpmgkmUoG4xRvTQ9kuAT2aPIp7LJ4d1kuC3CPGqNrC1uu9rtRsE+Vp
R3fjAk7OdMGjU7wfaF7uXE55i82IvVQ7HCMtYBSzxUD/9iFsf77eePX5gyD9ysHtN40KAJr/jqc6
RWkOkXpTiw0NW7cqac5qdxVQypxraBebYgulKcKsN0uPRhk7OhZw+kO5VDiUQoXnUw5Twcd+EJtv
MNP8VhPWAkqJT3NU7X08tiZgo7zEsNhoPka60FGrknjruyf+ddeQRL6XGhKD+6ryn8uA4+zidL+9
NK2VvxPIkh0ZgkusCGk7MovY1wHCk77arTG/pUpMMiWMOZW1sWNWTPVAvaOZipeRATrk5XDOw1q/
IUXtlaHhgFY+tiA9GLjqJ42RWXBqTVh9WxiyOK9FKwipQE/k9zZ0K5nV1dEdr1aAnKrZnfz0N1yt
8MZ5G7gT0Qd16nTgjwAGioIhEZpsAmueghmtts1gxyfzvNFI1n/pFI79dVfBaECoH/f60FMb5sAH
0F6/PbALd1xpy/m/OoVLyvwcW1R7eUkpAafXRpdHZlpB5+Xraho23+0dFf8Ue9tNG5JSVWOT1m/0
QL9KwgA6ev6aCJPNafgsYODncH+eetFeNz3Cb1ncVGPs5ak3HBoYv4hIfp6fKW73UH2+1O5QNCDT
mcQI/cbfEVGGXox6/FJolIW9mDRi6WgWHWienkH+84oHQsZZvuhKZGPKYmBY0lagcavjL5vvu+QW
JL30Po6EaqxOexAVDr8j608Xy4uIzETdZv+wYNImbbp29neJyMmzIgEd6QJWUnPR+x4Lni6eIxPH
FTD0rLoVdWDDkOMCIF0x2G/cPo1uQd/PKPHRLoZujiBvU5Qbcl6DUcDVwxzRStuynpl2o6T5GpQJ
i9G0uRQm39uJF4fJJIWwcEQxh/hXIa011Q9SP7gvUVY3WzSRRANpxBWioeHKKLhn7kRBnkqIrQny
D/3t8bSomBD+yANThijqLJlW31qLbzU2jobDSDOJouVXVcugW1eL2RYA7CR/18hcqd1qghrKnGt1
skBEYqZpxBBCRvFS1Gl6FYdn9Y8uSei14hd/ql09UCKKkOmtcNk9YGZBPb+XjOpYC8sgV8m9uX8Q
l9nRhAvHd2QU6ioucD21+DsHPaHitEsyed1F1/5xVONz6Uyf48OxNcn+qLzwktYZfQrVDCDk1ZX3
Kx3NjURHk3H8Dh8bcGV4928N+2p3nVQ0SdXe8kSxowF9JPyRinncyoJ2NNnqnwIfYCoCBh0S8d/U
iw1v841C2SmUslNCm5tBGiBkVTtRy399oGIdH+KgDD5MT6ziaIaRBsFvyeGtnExTOsjZTNnxRGYC
ckZWumCu91BfcsGoneqKejDiUrHCfE0J1TeGHGmFZO2WKuDOLkHauA/Ir2B35hclGWoqcYxdoRvP
WJN90vFtRhX/5yKZHcVpH8D2Z+GZKaCIJXF5uA53TOQi5MEJddmzPndipAb+kbvWeFhfr3VWQN4p
ZFeygjswLj/W/K5o7vQwrZeJdvhiDa72s7h9yMv+1Hd+GjcqptW28uKHRDaJKe4XND62dhSy1XGh
9a+JHGg0Wxz1ha9CU5vbn+/qsKIxq7/mj7459opaVjTRbkoXQAPqMV6Tv/tIiswG3mj4k5FdTILS
Q5RiOsAXO254Z/SzK7nc1OA9SAAiRAocIISHWtfYmsjVFjsYKzh8wBuBEhM5by5d+JH7lXoHWRel
Xs9FM0/IJ6uEL5pPsdLi3eiSbatzsoXOIQHyno8I+VwoHLO44sVpBsdiqOgBDH0kuJ6rgx04AZ7P
E0IhcmSBLtgiGqkjX7NwkZ9z6kReVHANjsbzvRiXE0zeuPUNu+RY4FRYy9lUMo8vPEYSYCNb0ueY
SgaZ0yvp/khe+1x7HXs1FOswT1bfoLkodEhfKHLSt72aAiE+W/W6LsrBcygBuKthbU53NEE1UbjD
AGshpA2+UaXEUa6JHEGu69v/T6YIU2CLtTVfitJy7L6n1pFju7nqyHTXZvNiY/Ada2aqM6BpwqyL
YPjfirXG+X+qA9YbR182W/zQT/EZPxOJmtH5+KHjVAKKhH19ZaLWMIPWm3saMIuQRrvd60BG+S//
na4NuIBnJjtIx9xbvcOVhuHJJChz+CrnJJONa0YWirdTuhJVhTiFyUanaphE31sT9lRGHXPoJzck
EAbHrKDAjf7WTS5+TJcil7Xc5H4YN8pP6mnAjf8z46FGdRIrznmqdgFvgV8llOZwByXlpOHBull1
998EdHMhYNzOR7OzRrK6wFc6TtrRfvVtiH1ZT76HyrA2H27Qu9G5w91+0VdpRlyI66aDm1InXcRS
aoVd9Gtf9K4TSypDi0PURomG+h3EBrfb3JCiN6uCVnggP2mUEpBRiSk3py+zZs5rXPagbhBK6Fjr
ckbg8SnbE8FcD6XH2CAnQeZ/OQPIMauj3fSMSUQub7B3Bb28PGfaEJJwHnyX02UIJLYOg4yEaHbm
Obn7mbzKEMMjlQh39/B8jQSht1HKBkVCDIWeXlOPamPgk8BMceuiuGrU+yMkY56+DjCddvVBpJAN
CFDFIClj2jx5s25EIchHOlm1QMsFbN81n9+NoSzlxpj/M2n6dIZD5U+AO/3tIlNMYweXPqLhjbIf
6Aw9pwDp7dqzeb03Q/Aq5WW53QSMpmCx1uZ9mxo5OoOPoeOqNVX1p2a5hOI+Tz+ivtMdshQaV5+z
xyuYxK6xmQJfGioIlYi07ieRs6QJ00dksITuNnQVRfCvrDY9RAGP5C/YBNGkdZypfmU5JLWLMJmR
sC0EicdxAEAF4jhP4lakFUX5Vu5zuZlP765OsXtd3k0V5TCyLmLYd8JY+FBJe30Iw0YOjBpAXmLT
lzHPscAsbych0X6BJ+NlfDK1aWNo6w+ImoSL/S7allo8Z/VMJIrv0n1I1cHrEB5//l6789zvoIps
TMnt8eSW0i+TAFZeDb76ofG6UjTBGmtUtJrJj815YVwwRKLb2c0c/sti6f7kxKkK6q7rP8UPnqPS
plgz1DLXsDE7ShoRV+SPN2kiRm6iIUjiM66259MsQPkmU1SQsaUsPBEHeNjq4pLYgosnaxJywz7r
CrSe4+zcE9zWHKJraNBsQYrSiWt4lGYNUN8nTCZV7wgMxlenJxyjSRFxSm4Kbbi2P0i2Mydvgwy3
ZdnIDKek8u2Yd7sJvQ6JagzFearfhf0UpiVdUESF4PhrwsTJ9bIOlqJ/1Y71T5gRkiMwe3XmpKR9
yr0tQ+u3lHaFnNGsaiVN3e4N6xnTZEdEz4EUTCig9Vm4B3nrby8AoK98om3fYbZwYQ+tr+6YT+of
LdBBD81VD36aHgy9ikaBX5bf/7A0nQUDZuaqAAPu6bJYH+9/BBD67LGRRhsOKl4FyuapcaBoA8K7
XQO2T5S9XpbOkKa0CbeHC1DsPb8T7gXaSHJL0zxStMiFL1sxajUZ8374rhJdh5D5EQI23qziA5K7
BZLElquoUuhQmwjf2X8ZjIGi/mn0/9h/Q+mco6oKoxhEmx8Q8L/PoivYfXy9r0cifvkiBfVDlsKJ
8mw/apngGv0x5xk/B7wyv/YDQ6i5z/VQZN/hU7KCW7Ag01xGt+MH6Z6pRLD7zBT+BykOwYlEdT4+
co2tIjyUPYH/dlxQxlYLYwh5A+cZB8cqndSTpy+jmVCPxO/PlzuJkD8Pc/1JhKIt11Te+hHcvqVF
EQQd8uUI6bIZPfKUYr3jZfqicgHXN1KhA7+ysu0c1kQxrmQr3PRPyHrWwNccGOAxCIVkpntbIVwG
AWRTDbXekVfpORHMGy+y3f7iCU2dIHFSVgGiaYrj9+5Oei3VgdI7kOQ0M+O/q6O5+EQcd1Os5w6a
Y8H1lrjbuAkoOd6kL0wTEa5V/fTRdQGoa/PLb/1jdv/T9BBjKAnekIf5IdFxYjBrlrDM6NxJlNPP
MTkfDV+c+jDKCZX7Y0FBa1Dkwl1LYtrIJqgR0DkvPR2gyg+SXNg64ze3LnOYjJcafJN9Coiyf/6E
VUvSRHg1IHzZfNdZ9wL3x8IppVJtfvCtKKt7Qn9N2p0aSUld99Pd2E1zRS0MJKN6gsKjadftnbUK
LQo5I/w7mPHSbwGyG87g8XSl9n45wktWXLCgyAebmalO6yIxWPrcMmDNEVrpuXjYNDWxa4N8SIVg
Ablix+nFTCsB/px8/150+abG+dj2c9Tqb21SRfj0odNte/WiptnaQZsI0MXF7R6CMz0EZ055Vp0x
u1JmwAxN93EmuYUFsZPrwSMSTunTltEjX7/B9iPD13rBscST+aYp1MikVOOSjj63OZB4RhSQjEwx
aCwfdPEDkUOms3K9uyx7eDYgvNmegg6YABGyyalgUUkvoDZGxHt8Jo8yKncpaWPNOTXGqrgB+wUu
IePDgPXByNuM6nHohixleuNIx/uWjzQRzxH/oaqNRmstoDLTVEZNby00lxDBZNyDa6JTZJWwqnNz
OArdtvEVhZg/eH8wVpgF/fpO/ltZbS6gCG7fwUXpM8AhBVy3CARJ5vs9IZD7eWF24VADKC825Qpm
3eRFyrGd6q6G62bqBcBYyREQsYwWGf8SvtRVE1M3hvOqruNqIaHS5h+kD/OI299NoXb4w/5vFQAG
TrWf0bGOYLaLYZ1K/8zJPGsaV2WoXozCPO+7GQz4jUgZz+hb5sQI6uHLbiULeHMF7nnesR+z4Byk
LdIqa6N3NSm4xe4rHctJyeDIbQnfO599iFQveGgjGZiqRJ9l9N6wXBozTp74tCayByumbtztbsGR
XbANjXcZCrkaJJQcNvACI9fA+lkCzOylNgkwcikQHmb1dX/F8IzLDPeMqds6ZzUJl2k8qNA5JYC9
75T29wR/GEM+myYUU80AkZxFh8SgUXVxakM4bUlfiViiWhH32tSd5qCTYy0Wtzw8pnyRLzAXcyQJ
Lgy0wGt+wgOqR/EgIErUKBb8YhYPvB8zm6eWli2OQOnsOkUswYjmXZi2sgSEkGThFiPUa6lmG4fS
aGOyM4axumcm3VkiwWhKNveVjdx8zEB2xvmbnL6l6SSWpF09uyNDYSU9rPUFpp2epzKtD7GL3DhR
NQVGDtQjgXED3kpXqYUMCXDYe+D0eA1i0HgCQz1qNLBXk7iM//zpgaSLwZNfO1LtLO5mR4OUydbt
nclDI+ddqctryQJtbKLNHDFLUHjesroq8Q37Y1aewZ1/0BxvU9YJ3EZdsN7dC0sGMfbuAEE06omT
Dq3V2v4yUpiJXvHS0XONO9R51La1XODnLHnFppLtzgVtPunzNWGWW+rh8TvzPbvMFfP6Md6Kqt8B
LqD2XISLSvicCZ1zvyOpIHSVKXpzkmzTPdbMNvVDKXmAAU03gkj1HpgoYAy/73liETxYt6Bodziz
bE8oGSvI6AaB+lYleaMV6dfoHx7wr44DtYKS4pgfYwL2xQ/T7rBkzqzVEJ8SaTfM62VENg7VXGZA
Hw2sS4PB1OmNvQzN6Q6Rv/k7Ie1rDGI8+6OJ/WFpk1ZF2Dg653/8s9te9BlrKrDMTnGvDiU/GsKe
SLhtqjMPl6X4Yb1HyI815IFrS3VwNJkcH2jwW4uEwFaa0nE+0FoI9j+AVypcxoS2g2Svbt15lOQB
7w34zOpOLzu5m8iLPJDtSbfZ92HrNs815zrhNUsqrEzpEMw1xV9Z2p3Pg6urOApoZTfaIqdrtr4p
Yke281fdphFBP7vvqsgHnj9mVOpElIQjMtSDiyvPxgzrCl+U4GO9Bn2NPrzqVIGNSozJu7zPFtBO
lgY5swEf1yy/iPPXiYZ9MEVletOaF8ae6Wcxe8o740lN7QxbwS7EGbNRMWeBLWDczx/Lf+8eoD/L
7LfiwJe8aBamSxEqaR+YxeDLwx0ltyEJT8ryzvvLv0Y4w4lWArXiVW0L54rjx8vDOsUX6GnnIznc
o25JTXj39aIdqM83+BMQQhPJyavdn3WYB95h9xmY3lv7P0A815loNM9VA4dSKkaXBe23I9rjjcgm
nsbSBhptiUZ2AGA2snCQDRfNxFCW2Xb8vJnItTexE6f+1mV5zGWpEb3zMrZB8iPFYCqj5Q5lM3ok
hLbc1aFTh5atFtVeLf5hPJ77gbUOLRv63h1/7cEHEKuzvzJtIqEcDSI2CAYBDOfgsWCFEfb82RhI
h4L+jy/XN6ct4cwa2dX2Ku2fZQ4mKIELIhLe0SQtEDVx5kyZHcOFsbjAqbskeiq9f3gSTYvUV+Xy
bpWiPSVgbZp2nFT4R9Lj2vw+LSEcujbHgAhdVdJVpj87pNJm+xsLe4RKSZZXjM8pnkoohrBjt0C6
NsBEgBu/4CmPY1kuxeLncJ2LvsLGU4jqTPmQl81aXimv1c0cR7vXe5VQfFlkaH5+uWp3BYv3sOXO
AlCx0kqtJ7XRUrf21juX7qNBlTj4FHAdOLIVuvP/tfBAoLUBpuDfHxYoyVX4DD7Xl73JsIzKOk/H
nktlkJxNSRGiUibzmcxBsdFvYMIhmM0F5YkFXQJ/WvqztNUr7XUIgySZb4m+KX8efWyLI0PKDKQD
319tXyEHl73Scfl9T9wJ/aaiF/blEc9U5HYnDxQ2aNcZ0tNSauFOU6pM/bxDbF8xZAvn/Y7SrFoN
6ZY1nprKN6bjcSiIAw7PAuTKfqjbyVQc9SnQBuhhwu1migtMfAUJ+tkdtGSTpW2SkuJOb4a0UbW7
0yPjskMnwlbclssvbgOKTrhxTET5f2fGqrx41uYaELsCgxkyEWHWFCYjuKEmyrkns+UumkQzBYHc
Uq5jP6WORq6lvoX6elIEOlmXuPnDHZo8RgeqE+LXX95cVHJ1CbomeZ8jDkJP6Yp/Q7+2m6i4a1bL
DnXQoDNkEJtHLoGnFUu06DXem8kqQDE/MrE+E0pX15RH2Rj0tpv3KN94VYkHyjvUk48zl9FYB+FX
BYypNpzS64OcGG0NbbwA3Fjf6jnq6yf0JSo+UzcVCfQwi2L9ekmcpBLoXOeAF7kgS3lmoKK/vWtn
YetPBibRfUNXEcaaC1CfWWej6pxdhTY/hwUs1I1ygIMWp2cfByAkUtiZ6Zyvf/x92rRfqPeTFAV+
DjGbd98R3rv1mMIwUCSs1sTVewNce9+cAAeuto6IlLU3GQzAmy69O6jJXoHua1utLpVmMFPSGUAL
VAKlZzdjPDRIGXEuAuuqps6Lm9sbw5C1CSQiEPkeL7V9bYywOz4GTJoaPlWGdD3gedfxrUKU1E57
fO30ZxPOyz0vIRZDb559q9SYU/L9uoUfm0qubnkygOISLZ2A/yW3EZ9JVgSDEb3Ua+mSHUtue8pg
nbQQ+coAiVdtwi7cWvl4YbijVfQVGCZSj2QNhZUCrphEBdwTD086e06S3kf0uvvYmJA9hOXw5FSl
OA/gNIjOqzZG+1UWfAB1gllJgef4TY3GMTtp/eX0J2qmXpcOZsb0cT3j6tcx10XzTmuqHTHKWqFU
C3ahzhdGXAOuXZCjunzK+8DCdB2+bom+9Bl8bUIlgs/UktJ55jnxW3hBWAbeBJD2Pl6UeDWnlZAa
yP+e/Nw1DHP/dCvgNgK6P6Ujs2km3zKL+hJAroEIbX1HFHCiwRLnmJk1kKw7HJhRSWyqSrOimh6v
LkUMM5eaboRG64fGP5FvCXw9naEGpBRyfGohI9D/E/NLf6pIBFLn+La+aJ/O0ijo8qoAvXki7M3f
B/9yut/nclylc2qH61ROGwPKp2tYJeM3b6OIswj45BkV2GQOjq/TbGcgvgcD3AL66mlOwAxtqQkw
xUlMMP+G/yqJAzp2KA8ej5woS0GxHEdJeP5AS9KgVhWq6Li8mxd+3qLLfDYsn9829uUY/1R55ZfM
45QQus+XzcqnSGE/V9Fc7e+Ulg1wwd/aeuNCktu2awnLwqzcpvM07loGtmcxiA830K4SJYGwBRpv
HuWl0DuKpKENSGSOm77xMHMGfKkC9S3ITfbl4tkfc+bdRIH6L0Jr8UrDrabkkBtynJ8wPyKHyy9b
DyC24d/1EpLM/2FpeLdg+5gyY4vGsljylIJ/4RvK49dMuEdFVz7Bj7R32qUh438byLHz0HK5tjxm
NSXQwuygbv/Vv2iK/smDlGGeRy/p/VxOcy0+DQu0TAWED1WUKk7RTmWdJSE2F/+PNcZq1HZ79Uj4
kgycZB1lHvGaw2zD7ALSnNuxibka14tWClIcYwW9zldqgXQKi2sYP4mSG2RN7qimEV2t/oo84Y1u
SkRN2KZvOeBTagarJ+USC7q64kOZslq72SMam3rscR/8+9OESecX1seDoPLXKDhNy4YAarLCSJd1
gIf0nq6IztfcyCsKoZsAoI8ZlqBK6Ujo0Oc1alyEjvbkkd8Ms3Z1Z9awEaiR8at7Bs7Ko4GPYEzX
qvfzwa+jxuFNlNUGJe7DWFaK5tWfSdVBKY+ZUYKybmWCTZbJNr0r1d7CzlagFare0lsDisv5cml4
asowGr6DTrK266WhsCtwPNJSJBpZ96c48A4Wv0uDrA+1vEd5WaXYT1PzOI26Ux2V9Ser9gPmifQl
R2ZLBHvSPa6Wpf+RJP9XkK42vyWRd4i3jUTT2PdRLjxoW6CVW+0B4y6jkZm77C6fvALHUjNFwuRG
LkyKS/+SCK+swMhvlGuxMreOLMTQoZSYVkv7HLWDkn2YPGS4oBpqwUzAJtBd3CTCIDU5jFgYSXu1
u5+zNV1swGWF6nLoAXsdX0q2TQHd8vsdX7q8D8Iy1KmnBzoMTRb1Ys9cKvZEku1OlQBgNn2RYjR3
PEZWqKBbvwFVoazDMzS4m3quovyxIrbQm3VCmhp+wsV+ytbdQSoJDiW0BNyTjKCFtTUx7sTEZKx/
2AZyfZuRGATYIPqTgUFu0oESfJkLxh39SMhQBsiS68rNg9ZsXXDm22QwlxllYQbShCvXaKPu0V+M
XU0WiPJU2g131IY76p1ayzS6m1/9Yi5Cj0NrimCP7c7T9iReTD9ydCtjID+St7hBJf3Z95WWE0Jq
LWM4qlDWd2iAe2+KP5xb0TWV/O/WIrM5YxVc1cRcaQCxW258fGgyj8Djfip5nnls/UswjeutZap9
jI663B+UY//Nq0fBGkn0pAAwhANlR1aa6uECY4PiACDOgVgOi4pag84IBNj5k53Uh/U4M/op2Qsg
Nam/YA9FE6RcrRMwk/QUZ+4ddI7516qO0+oU1T6ZXeEhrVo045WHdVLw3tIIGhDAV2ZA1qgKLmDS
dG7d2RnYYVqGJ7lH3c7cmn5gQY5gcsPcKUsSvTUR73PNTb+itvx4rktGQCgaMNEcsbSLq7oPeXVk
SnLLUvZe67e9t9aA+d9nzOOUoNJxBHVlrgDSWzqmkxBIH1Suo9qgtIam0VAl8cyBrcR4orwCNa9S
kMkn5KVtVxSuF267hF3gWHJDOsE336G/1JkXwpHDs4RYiPk+KnoOcX+2boaheXywGk5Pcnoz6p4j
bPR1D3vGfDEaU4WZDam2diyXNnsytm5NaqIJOTR3okxGURWrCnw911mYnDxBzXMJJiN4QHnKdTj/
AHYJOk253TLnYnnmdKL6XdmdosIboYOscROpKgJKw4sYgFONW1+Fy/jIoLW74OHqp0c4gyo8OVHw
5Rcrc+xOieTQj24iG97j9DtIP2P8DYfBcCj3HPiXRK8fHixPsiH3kAUhIddUVsIvYlscNIVjykDP
rnK7nCQz4aII+HqhtufgFFleQeUekcuKyTNKXTE+AeJyMbHHGK+Pjdbk6Ao2sJu4Wvz6GKhUwtTk
qBjPUurcHGkjsWgk8gtGIQt4JuaiFUUznNgtRXh1au2aJVOdg7DZT324Dz+MD0/GiHAemdReC6wI
0r0l/D0xRx002e2yX3GErbGzrqaO5Ejc/D+d4QJG6Haas7Bn8FIgUJktv8NMbtOoYXo7dFIV47+l
hh0ffFCwgaz81GYpEWwxuE9akmRTqqhZyC6AhXHqj0K6JLtQuicc1tOGvZhFMkHvMefqqsiaAToS
xKFk3bCSJhs+Rm/1Pbjuq+rYtt1EyqtUwdTKyc5qYpHq+HzNCUC7ah0x9FH/6f4sLSqftZTgeolD
7cJZszPFBQbsgbwtGH9OSSVYt8aJmF/84YdHXJWmU80OYuZE/agdRVJ69vySCuQKGOwhFDi4cQeA
H/7cZafaBJTylQlPZKRNp4YKdJAYZP5NWf0Jm1GQZDtJeM0OD5jEplbukBCGsfIV8FJmKDCG4QVv
7OF7wk4loIoIEFARnEAKoC2/U2SVeh14DlRI6alsSjHe9CDbjp/TkBCI7IbOVAWlS5ORPBRA2ENE
YWrrGgI6gRN0tVaQw9QClEXN57/sb2Js7nsnE36ZJLzbnoNRD+Rc2VUuGhGrHVQa7uI0RdTgIwl4
fNOe8YparlMbq2N90TAXxQykcywFSBtvnKswwWd2DrHXlGLjJyloQaVHnWQjeQuAk7o2kIjMDZ98
KlY7P6v/JpR/3RG3rGrXZLjQUj3WMAAPsGj9fi9gG4ex+izW8gOvtkIPMrj9aIeNRZWi4BMPRYhe
vlDPYGeHcSqEzqNtZpvD58zE9L840apXzCRm9UDpfyX4PGt9iGAHg+gNlb4HweTvdBnyY6rAbpIY
lrtr+UsJnFY/h6TGWzTX8+p1SXXXkn+XDl4xNkERzsKHGX26VGo0dWoQ1khWF9sj9OXjOf58tEcG
vSBUB5pZ6lXefsCFE1Vs47TKDnWQkfwIRocSL6p+teciV5YhO7Q7guMcwqp3ggf1++bj7PIwV82P
KIUSsjeJvGTnKpIKnn1Z4m83T+ETbKSXzVqD0JddOzIpLHIhKHaJXptqz3mapLG9KZY3ae6n+caP
cIYHm3AcOtD7t69jxniC+K2xXb8mo3tNJb5WH1IZ8wrveecWvwh5/qa0v8AJVUln2OSo9CoZa02d
2r6s7PHXlwnYdbBnuE1mH9DAibjo/X22dJbKi4LOk8ZGL435kVg6u3JNIjA+U2StAFUmCJuHMXG1
pm/7K6ej4QZgEeOzOke5uaBKK8/dmxNHMz/cO8V5AsnV/+2UUoZBetNXEawRPyHggFlbPFycYpEq
7xsBl7Gc6KePF+hHGf8ZrgaXvn53o4LX/1IWr+lYlYdl65moX/IYQEq3b/UAli/hwFR8TPad8riH
Rpva3qv9uxe7Vz0bQjO53bCWsueQjx4kkqPCdWp0wk9VQc5p/4IuHk2FXFNbrrG1jXonaZIes5xM
VNTuBTdBiIN7W4m8SdUOPwaMEosrUH1kMykenXFVREwQ10tIXffwjp5wV+bnyKZ0vVjO5lYH9uBT
zGm1jw2tO8X+hiimk3fx1J8SUD4BywOzZm6Nzs6h+XVXi+OjcecYen8GU12KrIWB/oAhkJtDYz+6
gXK7+tfDBqSUdNbEqXpYW+5UNXVQ06Ypr3X00lz+J26ZwvNOiXkchaX9Agsy5R1yMUJpmIcdJAuS
sUQphmIP70/npj5Lbp708fzW1Tu354vzQHhPYry8t7zVnAEV4DxoBRrsW6VuTKkA/51qmH9FOvpI
33sLx/r5tI5HTJkMerqxOlyT4RQC11sZX2GHPYFkKO5NtAD5deldGnQJcQVvrLhYVYUy5DB+RnMQ
G8xYhE9maBOSgUASaDxdbsfpVEJEbMUSFMd+gajTJjueYLG1NRErKuPAz+tdizCVt0ug8SV+vCbm
ZB8dpQAas8n0YJ+grmdiXGdPfrjNI++2un17a2jxzAu2mERUar4mGnq+o/VvLrmDEzBnoAUP/4wm
hhhzla+oy5cB0BNCBK/TsCIMo+Tf2kuH4bc4Mh6cFIFIE/pBoRYr0D4QFCte3UsMH+C8tIXbjCFo
qsbXeRSjZ/QsL9rfwVDm4B/McXh/dz5DKi8h2affsYuvKF+Zgo2Eek6NQ3GLoyBNXRYskut3A+lj
5BdUse9QD+zQng6RFcCCMZ/Qd+sap4uEU1kC+riaULxgMVYxfYXm9dtbLxFGZMoK9yQ/DgadhtZx
JmQrf5WEQcp+ZPcCPdrcX71kgqJxPa/uz5wKKiQyBkx4jJW4JQhZK/4lcikAmjmlvxoeaqkzIBDX
buSJav79SSkZn/bV6v4czpPn3mzYGY1qv9F6qW2cYKGjlSISw7SKN+Aem2z1DZAJ4EEK/gfsA19l
jAmDkk3IY+pEbjFRifwPW4JD0nhqsU2DMdrm6YyZBJn3kJtOtUj0KoflctF5uqCN4qotd+YucFX2
1/J4xO7+NugDE8XrKaBC2t9uPbMvcz8YomlmuPV+nj1Z2CGtO0Kulzl7x0qZ4OJ9Ls3iU/v3ZQXB
+9jKjeKqTyi8ZtkOQbaiXNG5VeIW85X4LgmkUTYiu4/kp+lf6sIp5ibeZcz7vsQgMen2UD5seKXc
sZfCmLaB56XkIEyHSXIrUo4P232yBgDTnNNd4MaZVgivrx/shre4Ul6KvyCS0tU/ZDqr62njZGre
39j9iwekGZtLt1jEE5PkpFoMSVq5rgM0DB6GBE+zZfpP/LiTNbJTNqvuk4J5tqxHsKijhUpeI3et
Ggn6UuEg+hDj8fQmZr08onNXiiGlyZ595+/C9DGlwtuF8dveJNthrio6gYGjgwNzlphzN1BgCB8X
YeQ4bObta9ejfeEYdcTH+xnUaeuq9ME77ZhnuM1fvgauemuboe8+wmG+4PoPaC3ZLUM7XEd8XasD
lBkAZMfcfs0psXYjURkAikuDAz94lwRjupHv0FGwxTo8C/gWpNm9ot43ugQMkdSie/m5D9Gr0Lp/
Q9z4Y1j7aXPoi4rl8KpwARSjEMZ8TLyK8KG77IfXNfWK+vEHSEYfFLqtbFYeEHx6tD9lqdHyfo2c
YH5YT+KKMTh0+FgqK7+ja/d25jijg0pC4gOJpscvZt5cB+NAMlHD7fYB1GVxk+17XeVeCD8oz3FR
vN3zJb8PcGkhU2B2vr6FDvjuHp+JTE9hfZHj2M1+AVqcGGthAST550HhPLzvGIMh7Nt4WG9qv3vl
xLIGqruPTimH5aDDy7aF/POWm8M+UuhYjqFWkLjfioWu1A3/DX3jcqTfyXr4Kc14O+7CdZpI6QSC
cLC+G+B/UgxGpdUARSTDT08EiPf5/gzILqB/tlEW6XFy5CZWK6KShikSYvNhE7JJ3PxhNAekHtND
j2nXNlAUvTsBOMJxc6jFZ1GN9AaonFmK7jCmA3hT0AKa63YP2B0Ny3TFbuNcZhLcIazOtAgSrLvd
wArSsxYq4l/nSPQwz82WfLN3EgmZM8XjJi5h9ePULiOOSYo9nLyzX9iIZIaxNh70Y/A/ms+MhpMB
pTcSFD50d56EW5zu6acGbttGjgGNpDwDsAv07Tatt1r7U0Aeh3SC4Y+6y9pv9lZJdKTBcwdOtV80
3Ku/jvjWN8juIyLjabCxa75Ac2PqDv7himiyaQTtEXXSgV1U6G5zIOSEqsb+XxQv7QMiMC2jZS2D
+xdPGtSxR26MG2rjJ4WrJwfzZd+qLFen7He+vl4hFR20yPjV1SDW/6PcH90CuhUq/ZPJRcj1cx7i
Ao8urJSlEtaF+MHvM/WcizEwDvhHJrm/HD1oaa2H/FBFWtHjqJCcJRkUuo+MlTE4YMk194MvLrGR
i2GBevg4lBl+4E7IFCdgFS5TCc6Ooom954Faa0TnzQ90UPCEOOmMFd9RJSVYry+4+Ovr3sP9yZsc
FPmppMv5x0HalY7gpdpxm8ZRXZRjBC/5oohMac/iV03Fl93Y8FzEnPDkYBc/d0Z8MufKOMQ9G+lv
ohuw8B1FoGQVW6J3zK4s69H0IIm1ERQb081q/Z7XpZHFv9A8Ea1hGeaDXleUFingBoYTX2drLDBt
3mVZAk9I6EbuzHeFInYPcCbzx9BDMcEBZYZsI8gXQjY7VOuIGiODQuSEGMJSyOJWdRdbwA4NCKvQ
flq1LueY5+8BPs8R5EuDhU1VsOlE1N1ibeYMNDnkO5cymvOBskHrFl1Onu9NXeWGF8gAw2Ve+aYJ
SnOllZf22PYnZNsxTuKk48do93QtGtbX50YbgPVC2tYDjOJ9YecNo8KqJBPHKdQEeU5VdjyU7QhZ
QBtfDbCFHO4gmmVYRuz/D1i0XTPiT7NwdqIQvLXwFnrF4a0Ku0woiHCJnjAdG7GJXGELy4uKicNi
ZponIQ0dV7B1wzLpk0O8RTizwsR8XKrnf0JA+yP8ybyMCHkNFpUBTbmqYyGiBZXKtt8vKg1X38oJ
u5Qiydbk57PYYGWiN9j703fmvIBsLjgzxX3esgwBuh9wd/uPaQCOmFdgJ/zKOamjheOlG2bdZLET
BmDfukR0J2+hZOyCn6M9eP6/ikI+mmhslbBJnmU8sRSmD0NjwjC3Rgt9P3UFAoyF+fQxyEGTkqUH
Cfv+c9YPDTxk00/5saRAf8QyH78WtNSOpRrH2GVzpdGgG3W28/wGsnRbG4KeWe9//MdGNGzkUhuI
Rf0/s9YBHf7BHNp58ZucBM3SHUX85ozGZpW3pz9OA4aqRxg3MCOe+mQtL8mB5WCTT8ooc149jTwj
YufIdL1XJalnItTIbe9MyNbloT1WAMHDm2g/dcJyDbA4pOWeRME++S/8G7zXPco5KMbxh1ZS9tLh
K66Og2uZD8EiZ/XDpGQfJHqwsMTJ7k61UD1qcInj7QgE1A+u1e2uj41pAzjzAs/Lj9D7nXki0GXV
5PhlgLRwixP27Lo6DxlOFROuC/339xzvISHWplhsyPKL+1thNzVOVFm286PwfI6wohkdfUk4Vsbn
vVLW87aNTe8jk2t1LRuC2M5JXS8KRb3VuloQprQpVplSnd7HapQliuincWQr0RQUtwe2HNUICMZo
X9YUfgrVq1bP9CqfP9tnx6hyG9LZaB5R0gu1eh1ZrR2PSfWRvjNqmwObSDgNYyG+K5C9V/bTtoCV
i+HlNWvB5HEnaFU3lDnZhdx4Ffl+wMJXB3T2UOCxXcM7r0SPdrg6QAZLVzs02CDelTQ2/Kxs+3yV
A26VWnK+6wIRSSnA/Z/li5n56qP0kfgZsvgyePGa506EE4OvulCuwFr3buwopc1OSSJy+ZOKyuAe
6/+iIBr5c1n4xJVOBqNjvjhMPQAyYO87ovy0zG4rorv5vWBi1Cfdm8SKzNWqttWQAEBdm3Y6Msrx
68ixtUlqGijYA/KxhMEUgAT6uLp/xou0DiJrdPalIov4d+TtSn+PE9TbpVcyi6kIsBruZ1d/QEXY
pSSKpVTvN8v6Rg3fri+GOHSfS/eYh3fbNNma+n8drVnq0zA8W82EU77sbzvAw9OJFbhISfHdyLyx
CP63xmjN3rlnJRnK70BHcjOcA3BTT959trWQGQXQXcSpHtV2a62MvTWZnItbkQtTkc90LJMduPeM
lw7Q+tJ3fmBnF7gFYHuV6y892YMQ4URVIaDYte3NgPKKrMfC+uQp828Lnxu3923+VcD9ZMwRn1xk
a8uZM7Jbe5XSQawi5oMKRYSO3/a+HWD5+yBLSzK/0UJPPdEXW6TRFZAQYr3DmHGdNbbmfXSV1R+T
TsuYiQcw6WLxcDf1zG5ptrs6eVSTib2zetkpnSpQsnAn2skzQxbH6MyrridbQfDmcnK6uf69j43C
UJZaOaWySuLMxfECw9D6tugzjxiyKt35PvOpRaHw0+FmF4IDKR71MHGa01paAKte3rniCLA1Pcb5
lzFipOuLTscXBSfP0IQRVzgt7Nxj9ad9FZPVWtXtjiauUC4/IucWieyz1R8xo9tUXWaQAHjhsJP8
N+WY6j2xGlgdXdjA1VGbxajjrhYAhr+vR0nRX9SioOfphZV/chpq+gQfbKNUS6bEW4v/Gg1KmEA0
JVfNrcmd2x8MOSYUwgrJurwGKHNjs4nA/Pzt63UyMdB+j84nyHc1PR1qEV+cMPEPhWYrwOKZtX7j
3KVy0eswuBYKrXw8BxN9iCbYBWvrOmvQGt+Gus0o4tsfySBVM6T3yxhHKPuq+cu+64Ca7eYHiwow
F+2fmoyaGASuhMUsZJxbAbop4TfBXFpwxh1PxmiL3nOkZTOV7zbWOY6nEWSlv3N78g/bjNMzhBeC
RcI89t0UK8tY2rjFwPqPms1oWqy/lRV/o3B1JAGjSm0x2rdKXdIRRBEl5dvRyFGMGXxsKLkfkLwq
5cw89kHFo5mzd1iJefGVmj746JGOWHPS3WywAOizj7Ix9E7IlBOAH6MGkiS+wdrNFs+L5aLwQStD
T/5t4X7C+VfWlj6faXl8mYZLggTnAi9FYJS/SBY/R+NBEba8PtnowqusZ2BtYbkcgvfp1eUjWatu
f6o82h0v27LS6y5YrHr4M117blb9rGksFRZynVvHYvBaH8mZ5NByC+uajd0qpyCeQqLKHBsFmb05
9JwmKSn9saiDvfbiJz0keIlZK0RmKgWfsFMqBO3VSyD/Lc6U6OcRsxA4CSvywVnhmnanJFX5/jVG
H04WC9XsfCNlCbIGvfSKDxC6I0dxiN67QUtVZeHTjCsYVgn559lVQ4A/zLdbaAgL3XU5o40rNE4+
FgnckyEPJMoDBxJtbyXP0xWUkMfiUSUr+mear4dONvZjKOu7lLVj+HxY5RlaQL37bOb054k0mslS
kd4XJ12zTfbhuSi8Vk3T52Sm0wNuubF90KGk7KrrSt5wPHKaX8WIkQpQZ6TEfmS+0Jk2zQQlOZNb
/wQ61peLeTzdHS7RlNi9uQmUtB3Tq6Rum6k5Gfif2Jts5DF+mWXbfOWjWY7Qo4hy7V26YJKMGd+5
xg+5o3UQtpMgSEcFkk/pZS5q7os4y1MSL1aEM8fbIEabJ13G0xrM9lna7f01kmjV0CMfmxncGpmj
ivkfAXGjG4yzts6X3cUaFofoaezSHwHxcT6sHM+YtKk5lZK2bnC0DjGO8DWWMtRmrjrIxFatzx3c
/Yr7/oOBVHqziZ5DH5o7hAU8G4mtMRWV+qZZZUcAuFoylb066xpuckWwrCTCcS8XdpLXc7+MnDaM
3m8I8jI+zDpAWE/r/Hg8iWJCJNkgfVqMc2k23uJAmeYyZ5YsjmRxV6FfyMnOG3KE8EBqICj9BWC4
x7RvqllLoBqJwaMh4ZU8qxDg/ivbnBOkSV2NbDtKTAI7+hWneUStubz81siqew2OshFIJXrUDRyW
rfo9MZh3+B79nipjjGc2zONYVx9aD7Z4k5T5Uyuxd28Xg5kCXIvETSHRZXvJNbX88XKiapQqqSDV
bRWvEWwY1oanSM4zraIyWvC7BheMisWmxakBqfebD7cR1qNPxCYkWSUMmZMjq17RphGenZ/xOxjo
blXIHSf2U3W1b7sSgaskMFbhDdugyASahb75Aecm+z4caWvjvBnvElt102oIMGWwOehAydmecflV
ZCXU9ng8D63ARPBfe46Q9ne8cXv+T4wrCtiGpM9iTgfALBSf3uraWFuOuSGdl8dhxsG+N+Szd+Ta
Vc8Py5zfumjLFT+e7Os7a/TnY+kaDSXcrtDvyGB+gkIS2YiiFPugVtfriRnpZgsrafqclM8zs5wh
vTTpmP6F3N07KP9LcuKTmIsfT9+Mfe0Cpv5wgMJRI57DE7jwiX76m729ZhGnTcZ/7MaVTY/fT9/D
hrt4mfVBZ/KjNOfgs75Eo4F3KQ3mfOL/uB7wwZd98o/+gqiyE/0NKzg/1mybNHIpvAA+zs38SH28
vpMUv2TGCX159t756S2VPqnElewjIUSR2pbrYQD9luRtmwyMyD9T4tA1rZHgOMbILXyOWjzkNRpo
zPGCySwftuo/CUSZoV2Tuw8OvkXAqk/NkgDUeDopMyzwUo9m7ZBFpmpxIZorvCHXFHFBtwZ04yNK
Z7289bvQjiEk2XKhIdedUzi2by5jqmIxQaJCoxhWDcgc13DDGJGsYWeuNwUKADUT405s9S8mO2zR
fw54/gmUPj37VqzDHVqkA8etIDfGzfo4wC9nHVm0059MuflHH+TDEVDOG210ESSR019RVCIj62gH
jX6NSCTJV/0ZiTTqcHlJ5z4w+0rcrV/Yj3LGgoqfsvm3r45vKK4z/t7OrE4fkH2xaVNamzS0gTo/
lzeji8RyUKpqc0av1Ftc75wPhLfn6+NfioLO9GtsR0K7vRrrpdIRqy5UWn+yzqadrkzom+gwc1NV
aRHRmZreXsrN+odT8IX7Aznnq/MKymqUe/73ldKAfW+B1r5ceu1ryUfUKgHTgqn4b8mXDjiUno2U
RWs5LeZ7iEqCbUcBPv/9TnOBM6QXYOOWxRHSJqYGSIZEKBfFUmBeC17vXYzd0QhcWQYjT9SUCote
yUkWFez9pwTi4WDcs1SIy2SU4+7/sTODiAo3ok/04vGToUs7zefbtnn4kgJtGaxaVtFf0NwhBHAT
3KTKQHI10SzL0A4jhJTHObI94FRRzTJmqJT89ImJKeyzfAWMzPXQuWKgUISgeBwZpfCOeILrrKLW
BPZJqCGEzo67FNsItx5XT9qdV9+nm8EfDj18e0uklSFZVVaoBFB7x6Pk24QP/bYaTb7SiugWJS9B
vxcOz6fXtAXO5p+1ev3dpfbUfcB8CPgiI/8Ak4Fy9QfgGWF6DAvU6mwS+stHfqHf0MFtUcEubfw8
cwlawzj8llgRvm6M2jvA3SgHjMwAXge/SIRsVtOzxDPCGQq495o4yIyVwm+08139Vn3+ZO8Nt79v
/HqMGX9/JvolP0KypCEA5zRs482gbVHB1wUeVQlJm+uTHyf11W7QoYFuhbH8MJ6VO532cPGtOAWC
AqV1/QKDeuoPo+AqacPseWPrWsRVPQUrR1OAZMCwe3KNwqywb6Plm95RA/5F0xu4ZZpGk17RMb8U
WyxVl7QZh5iLpp2YurE4hoaz0Eju89h2rTZLuCcP0CtiOk/sV9kkjYvIATtUaPD1bJiT4OQjLQ80
XZ8Kqt+EcOiwyamT/zoUdJ+kdjm6FsOGZhrg4ktDq9pi/K1NHuHZs6iUx3x0mq9twfjcfjY0hrRJ
4BodWzHS1OkittUqTVzKV2Wfss59LsuwEaiKBj9XHir3Mt1dyBH/RkjcXdsf9T2LH8jQzR7WdH/U
XTWDF1aDKBMq5j3dRF0Q0NzvOGbXP9piTPAbfpEPQiscV3x+O6/3sX8fz1YPPbSXK9GDgmv+TvwP
M+KK9W32EigPFfy1SbpxeYxXed/wo3qfNsIfProPU9hpuDeKb20vQfQ1rNEo0r3T5VuvJdDoOSjW
3tv1pJt/WlVfF5klzZrTgWcEyVxg7tNdHnEBnDZKAb17jrqzrvMpXZY4e8hD1htWwna05uSO6Vkf
CcC0+S18ZtNDs6L+A5C3UQAYALwQuNXU09aAg4/XFpQO/aTwE6I719aAO3HKaiHdnrsZEZqFuvsB
/KpPlsb0+7GKGa2/SROnSq5XMUN2Wkmjy31DrscfbuqRdNi3HCqrPmC6NCcE9B2Jh+xH1ZnficMG
bna4Vm9+THX2JTGQJe08pGBMqmtO8kmK0bJ6OnM8s1/Dkn73XACR+az3H1eisHNTYblnFd7PGroD
I0wghj13nakNlT9pP9etQ7Mu2v+xEzX3Rs725hWtMWE+rduHKy56L2TUYmP3doULmUM4CgJmqohI
E2GYRAwCh1QVSsNxFgVZQyjphQkAHvEgyWKPH7abszbAGs457In+NMw9M1vxxcw1T5/1ql6LOdxg
hhZ0r6wO+mxIvIT8GJStuVCVoS6yYcuVBBKcqyoZSJMZtvrZPMnNA1PiE0fyDFvrHbo4JTF9cBzC
Z1+BewK7LU6RRTzQQ7CTjJfT+Mgq9I0gtFbTNqo0lPzsgFuFq09kkiEeJFKuMi97+tU6c1t+qzzO
A7rfmdgys9CuxZPB2SHO8Cp1r4m2/yiNdevDVgbRsAZuIKLXcw/1tGJ5/hwM6crDDOZfq9FjCm5S
NGpNIJeIiuWsYIULDzwkHMR/E8alypROMeGUsID56Yc5fPp5H+ef3w4nncFXO8ItGfeQqHvzPdFf
SJWvvvcippiNTN/Fjd0Vu6yz3mD+Evw58gukPZfKZCbVFkPhy2uE+UycUIEzXXNVCSXBUvuQv3ne
2oDN36yGv7nonr6usV4K6TBMya9DF5kK/oVRXeodQJuNWBfJk4AYtSaPwarsl48A9iaTtUsGE0px
ZvEmpMxkWZK0TuDwGfHH+FfSmvb+fwJJo8t1OU13gVtxJNM8htF8TYWyo/JQzxlz6UI9BYColT58
6LMq0Hb9bPQXomil0IwJuv9QWmSH6QiiHf1ZjzFq/d6kRRkfN0rKQ9L6XtzYgS3gMrecepBBReK0
oXeCROnQBl2Tuanue9POsOWy6lnBAwJxTsUe7xLR0dJ+49oaCufF3AYPSicf6hC3/pgosSMznWx8
fiL31DNqHx1ohmtK630OsbX06JwTzo+Jmc2XhHw4L4TwXQEmYIC0xWf0uJlBc/Lac5TJVAJmF9TW
fac7DoRIu/SsuRkKGkaPLTAfxz/RGVGJJ+NjY5Eud4oxeWZ1RDx9yxkNusduGvxv6qQ4vUpyR+Mm
U/hUVQi/0Z7CsluBmZY0WqGt6tIAWKJYKPDVwl/iAjcgVTNG0cAjhVq2XupZrqnovXfAzfPFWTgI
Jxeme25NtRVrdicwkKJPKrEfEZ+rQPGAZEDrN98hybL/VcKNyIe4HCVOAxMwsCZiB6p0byAP/4v1
+Ftj2lSvWjOdMCiQYdCBbqDfCEl0M+PdOTIvN/f0HWcYTKDdCQzw6ItuGtjQmNLNhL+OhO2ATIM3
R/a4/XU1GN2gQBPRUsC4lT8DmQrsFgl6qAGVMg/dW4gxVrRkMHu+ct+Tk3veV3nrS4VpUXBo93HT
jQpiQ8F1aoOrGszLnVFZjb9rMIdBpX0PJAiaRboisbtF2IeV8oEPKHpnbMCNmTSg6VmsvdAQR+fF
+w1zY6eUeVvQoxrutEfzenJz2RGL6fbDBXZQnSkVfqQxktLN3Wy9ATC7cw5yFTa7f/5cFnMgQLyy
Fh43cC3r2ZEKnhsubKr1AxX3rSDDpgW5GDDNIVL6AAOxXRM0Chj8Apj5pG+7JFpmwNcMSGy3kcu1
kx3JsQho14Kq4frEV+5jedWsAqWTzIH16iLZZFxpgVodk7rZA8tDqhaplZmzgO2Hrp6/0CKKcMkK
lmoAnZBtQp/tkXMudw5eT2bmuYhkPReXQ2zZS6wAEPPtP8hT5rFZgUAb7Jdjzlv5W3VDOXr6MNiR
dVojAOnnjYiM9RXudyomwdKDzBPdVV+Wpf/CEEG6yfOwv3Jr4AxAsKDYTXlTIB2Rb140ZBVTaSL/
Z/q7L4VVPLyyZlnbgxfIr8bwyKfEysDAvi16glsJQVWh80REWidxRvgGtQ4SMeutSNADqfc/hDiT
7y8eSaE9mTQ19f/oyQRBCFu8np2FLHdygbHc1ToByZESJm6PMcJ0ow2bk36YuT21Xw++tSiG2J/P
t56u4mT3DcvzGSYOnaEjPjweTUUKFi5MWKxvyYSt2EOCibM8bN2JA4gdGegx+MHy7DsBjw12v83T
wLeFlGaS2hfcjwh1MOv5vrPnE4xHEBFZMHjSUz+dVBhop/UBR/FwG7npHA1MDLgO0WFxpIcTKXSc
S7unKPpRWHiiC5gGtAAE5AWgOBKSMpexzwq15Nzu1xlmNCi8f8039yBA0u7Jk6bGfLaMNqqaVXPD
GpNH2JTqPZoAk6GClbnCCM8pYo9XRomNoIQVnW1jijllf/cYjDbEhYhK177qRWbz3pwhtDyMpfQw
WoNtqEOJsr5yUdvVyH5CFXIu1KG/RYdMP8qy7I0rRh9060d5ZNBpTfpGdlVz23rIAg4/ciJf9tp+
/Z2qhlnozwDiKgBEZGCAOhrXDH1pwux/nh87blPQAzYJMIHc7VYXnaPnXjE7vRsJ0OfVBvY97ri0
8zCXBYBeQVxMCdGAH/arU8RWmLxIEz5IQbiUqzA6YCrZvSDRBTDWrrSvWWHrg2oVe9/+A8Fneapp
l9A/vzlzAh0bu9drKZt0ABiN/bYD6vSoX34qy+QP1FfITVFcXgxrzjynWyCkoMtQ/J5XjaPULRGR
yHQBKxeCYkGqkLngB+lSN3+O5SYYRcpbPG6accvfEafPMUKfXjrYhO10inJH5JVcGcf9XjSK/Ext
X0Qf326ppJAYYcC2NTfj+llJD08tb12Snoo4+ke6d/X828qUqGiVNwHMHXHwtXc8B1kTLSwSJ6Dl
MQZ2e5OYoLY6ruRkSf2o/zRgeB19DeWVRWSKeE7AYUQtD1+OLRwSQD3YuwV4MxDQ128yADTfFU5e
UeiXfLoM4/mzgDdqo5VCpAQhpKaJU+eoYIxhIsQHNh0Bi25JepPkR/B2DKKN9ygLmBTkzBqgcEw4
+WPfwqAiBiTKti+bBQUa6dnStdh3bI5mdzn3TavMWqIaMsOnjtBPPw95ea5/AslO/xwom9hGSGvn
KahbGpapkm4YQSuH7Prmc06f8Ti4uwjqg221GT8W0bJFFeBDWw+fIz+WWx5PrG8k5rWqEFqeUivq
10d7kAQBj+H5SNdZbroZJ1wP6+IbDtq/tUa1XGu2h30N5Jx7z3qug8ksJHam3mTewvSIQ7pzUT/m
sMFTw6JAvlglQm5/vL1dH8piElB6k12WnyXTuBc5gh0JWi6M6YgwPi4N3t+2YRHn+gu9nAWhEEvR
qFwZZfY1EJTekHfxyl6cNRyHApZ0rzhrWwlbxiiYWdGA0HAsm6OP22+9LvjLnTp+VY45WKyOKCbF
hM044AvqbyDGLh1eC8CuRTbZlojQcdimesedp+jNP11LrJQ+cIEmX2cYKU2B2wbFNd20qM0Kx2Aw
mQBssYM3YcRRUkFzyp9dUwmKXPErqL/R6js/oaqbTPPNlcmH9SZ8AecRSeNyDr6kdN0Nehejw24b
GSMs5aV7J52NRxlCnAOCDIA4Z6TuPxVK+RFLQgkhldDOp90H36qKGr955Qdx2mt0Dj7kFJyRQtgc
/vNCT2G9ZL60C2lGPK7G23BUC5wQTPN+HrU42Hq2FByO+n2vfUQ/OfHk6fcY001xOm20zWkpmvmv
9fuwAZj/qs7feBhBQhG7mEFwJQ0sXMA1+jGmzsJUsRN51pMHdUbNtPbfXex1iy/WucGmo7HhsFQF
Md6B6TPNdK1Lfxz4YvQVApx3tZPtpYMCYhG8anCrN2NlfKx7eldjh7Ctbl8cCY0ea6mr1ObznIKL
cwq/H+iTiK3F6f0asKNYysZWJiDOUb/qlya3B84ZcErEOzbvxq+Ln7TcvnfVGco79isEJLT0xdAn
DLg29KSk66HYP7+ZpRo7UepxfNi57voNNcYyR1+evhwJ+rjJR0mj+++5bwdjrXy+2FZ58SfqH3R8
lX3q8cdSxlnWFy9jRoxRy+F3AArwBXb1FA9/GXyg7OXP61KCpcu8qH1qwqNEH6zCrbQkh+f8gfiU
qCWxp5gTtPSTeIzdFed/VVwA7x03ygSeAo2bqoCea4YuPoZROuKWAZDA9B0ZhwZ55e7rWbc4kijK
JqGGVo1IabXnQLbB2DAPMa3fLhJ2+Lk/BQ9vCSrfkhJ43BU3OL1ldpn3kH+cNeTtR/pPK6fLDY6D
eJYrqLBzdL93/yr+Su2dOdjz0UzD/yDMp+/2GMyKMzq1k3aynFje4fDxEnoZkjfC7BvCFSynyWOj
8SsMb6DUtyUbNlTT9dtt4xDM/PNaVdklvfbvHfD7ThA1WFaI4iAUi47Obo5kTCNpsWhBjAgt0gmx
eapoydX1dLrJs405I94UftHFKhKQ8LBNOnPu+Af3D2MlQbKp0Ye19p/y9CAaoyRNZyQz2x86Z09V
jE6DU+zjhvO6GpvJQKIW9QdQBrlu4h7Hmt2HI9OHGJqirkiqjH4xHRS1Z+cZT8Rn+xAujMxNgy2Z
LZavoFcG7Vb4mSTyU3W4l/2rL1+n02iGSJH5HoVGVF5qjSFijrjbpGob9OrYhd37eO2M20cMcnQx
/jrzSwLGZwK1uRz6ljuf81wStXRqHQLjfZv1WHnpDfnRdbbErCV46Rof8nMEWU+aNhLrwWZfeja9
MCDv49HrSw7DUX+PLu6yccFT3C4Q3vOzGuGkjSvJBZHPekz+27RBtdDAXKtjrFTLCA5YPGizgHOE
zS8as2XooeYtwGgbhQy1dcF69wiRtZTfnUGr5faW3+EcBMaIVv6wTLxL7Ap7hp4gmTBmkHjRBtNj
wGhxuuo/n3X5xZBUoSw3EB4O/KYlE/OLwGChMIwUryAs9LXNpOMXGIf4csS9qpsAtDvNVLrYYqRj
nmriOYw1w3UvE8f/SbPif5QwLS4H9j0Y9HEocaXeCKGOHeq7YOwW039jNcCrJ0ZRcGiMjcdKip/3
1PNAs+9v+JcqBXK012pGi0TjTi9IQYxxBmErU5iYRdRP6KgF4H64I681Q4ITA8CApZHn+QrC0tt9
YdXj3ORkzbA8pf7ZT+O1QKrTXAzwPidnMlnE7aTnSSE3e3I28EeQ9mqnEO3WcKrXhrvUb3/wcN1x
1uRUHDTtusDzDH08GN07O32e9Q4a2hqIUQO8GBUrYkXceS1Kr8+piT7g57Nskr93mJBO1F4Qt2Bm
Mlglsgzavgfzo4kkOhkYG9oLhxwFxR1gGeuQ9gS02/MdBb5rNcp9yZTK2Mha89COIj3daS0eD45z
yhsk570pPMpjXLId/XsZBUPlfUBrJm5iWv+0fWa3q9M2vQ5ZdxQvPluf/1UmIi2lvM/6w0cv/rse
01F2vVwYyIA5nnDuD/OYX6Wb0IZySps95/G1fTRdeT+tfktA/7WuZxzDb0BoAWXdYi4UmlM0+KO9
qaQi4oBeS5YrHlOmqXQzuyBbF7e32kF1YEXwB/wAXXJVQYQVxmp1BeikviusIqfAY43n0yXn9CHC
tjLwtwuODWiqWCtQpOhJk8UJajbvenMnQD7wU//FFuQrN3L3ZRTkN3o3Np0hFwEG+mygEcEel7K8
HlFXfB9IAPRgZQW/KdPU62/IThlC7OmIPi8R44T+QY4JDi+BRZFbP6gVTJdsfW0BakGMvYsvT16M
Zt3DrvUwFiznpaiG2riB/E/nvSGYglHjMWJmsr48Pi+iy2RFDzPF/+Mul+XZ5AhOaDu2REs3yGjU
NPaKskVAIjwtjA5Tz3K/jSUWapTzgbZyPKsevhrfX7+jpwWy0DXJWRjlNdacWou2+1VC9UG4iEVl
Xut9Mkn/9p7RVVYTxGuvxyp2vBGBfcl+zhtmiMUSd81QArTGZrc6BTcphXlpdUFNmqGLqDjSAsIQ
wDx4uZZci6Un9ix/yHwg6B7qFSCTDep7P1VQZJ87b3xQfDFKxmLx1zVXSS3FkxhA18DbAMp/GJI0
52tMg/XeXH5F/GpL7tyl412V8SlvrTUSqRcLpPkqRdBidbLMoi447i2ejDQpg3QnGXdLAh5fJzaB
eElEjkyqvpXqCoIGy+OhCjFL9zgx4/AMOILDxm2+qSwaq72B5UyjXKNuZr1X32RFVCGtcjVIx6hv
0Yl9nWMqWUnJFyXtxT628CNhb+grGWARL3N+slEZvREhpD5s0WqQdW1M8R2/7ZpSs7d8Ny3wh+2v
9RKC8s23krhcrwgIwre4YvPywLmHotLoxZzpdyEu/K8Fdt+ngWj0WZq77FMB2RfkhpinEJQu8ulL
cziHwPwZ6CAapArfjSIFtcNOojpbcqy9knz0Orz+DzUfAwmVrFVC7zJKbE0rW6VKUs+GPawBBA6X
idTm7QBRD3GKGLaSJhB+2S6Z+Jr6ONXj5TZHI3PC7eGLrMGuwN5/h3XFw0mEBuefPqIiUnE7oN6q
T2D8SEkgE3tZKD+yQULkIO8LOtQSZOrez6Sdz70rOd4hhiMaoXE+euorjQY0RnjkbW3siL0SHtiX
+rcz4cWa/llUWAD5y7jF2uYeS7yZZ10CbFv2YsCQ3YJMFX3cERwO9RcXKpDiW3SpHMy7MM+uB4eM
gVaPfvWyQkjpJNmlP6rhYBahmFZi3d/XZYgWVmZUkoKm2Sy3YRSJBstzJZONunPG1ZJHhnxtNmcp
mj4wkHa7W/GY4IlG1zRwho5jeQcng/YPhrxh4aKyTzEkaZn5+kyw7RSbFs+j2ggl20RRbW35UNDL
bl6T3tRGBgB8OytNYzPd+RHiq5Qd+IkoxJCBXWF+Vvja7imsoWUJxRtX0OSCkeb+fZwfDF0Sbcev
rs+MgR/ZAFbA5Wb9F9BG2l27WnhVJ1QUtcAo1gYVXHbBKFy/0w3+1yfi6EHacXtk99srvsAwk2yN
XuuxrIs55TLqg3NpinHArBcJUR0L4mMRIAQMbo7K4gkb/ZqvgVDujzREz1iKmFjWnx5afOh1OPS6
wwpc/xGYCfffoclEVhH5CjJ0JHSBn+NTJhC3cBlcWZDiC4qh9mXHeBS9wgBVq3xwUV2TiosiXFHf
oUOP10BiotbToiy1f+fOLU6Bp0OD8o+0519Tx5/KLSzPYg7o8C+j0TCW6ngnvScQspw2ht1hg/qz
Y9nMxV18APPytPzYo9uLEV7El/dQxnSdEo0MsQb5uTw+IKTFnHzTjpwNGKYNf+R3THqgYlVkATDT
ErJCK1KRQaXyh1aVhD+ZDT9ykPZPJrHYIylTpdoJN9bBgEH2cPiGMkpAc8OcTQmr4vkBnRttwL78
J1z0qRT8jh6IEqSyTl3W/VQRYdJo9M7aYLYjntRbk3z1dUJJVrYa0dg1R3MVkC7NpmOUiy4rWWKZ
3VnNFKSo2saq0Ff0qe6OnMioJDpY1u4cm9pBjvbffv/a4drqQS229xPykOrBwIDUycXeav+bkA+c
7XSeN1Y2BO6qJ/gh7no4EgKsn+vijFl6xiHHYCAEeXe5oBy2FjAhwgSkjPj1730cALWOHziY16w+
LG5sJPkNfb9pZ83VfrhXWSkHGX0nVEk+z1CRBdWu3TN//CNaX6SR0u6XDlWMHF2Xfix/ALkP6cBJ
KuwzdWQluE3WQw6whA2nnBzy/c809waU5XAFF3A2duINgX64BcpbkXf38qG7igQfNRoIz4lmp2uE
tjIGiDTkmWdaIEXVWIHPPMPhFE7bAtzfU6GFp4ToylD/4SLGMhdaIaKblbsAqWij06l68iEssnCT
Gci6VX2z+0Zq1IbM5URdzuvN8F6CH2CRSEiDsvz9XvKbME/AePgNlpWWnFXjz1dgaPNM5N3/syQA
R1gULg0oRMFM0Xud+VJldKTntCxv47VFHpiWWndyqkpEi+HQ4S/ZyLjEmRB6FtOxAn/ud9Yvn8ZG
IgDguqA0isE8eTptEB6aJHeJ2zyCf1ld4jrynSKrkYG7MPEZw7htN102Oi56lYZvmzdeKA/gwW3g
3gfEcDiNWqrQMramduBL8CNI6seEgCdXsx8B4n7SR1jUmyKdHpcVmt1brm5nBsNSOnfVt4MUAfkb
lu7vT5RV8susHRoU0gDGNu1YSLLuKBnZXZvUovOLs0IBKvCUUKLUBTFOkw9dkFJsRoUb8IgNLA9X
fxJ9yfgZPhBSDQfANsHPj7rich4oUjjZR8GFn/aEZGLQSWd5XIHqPRdmsO4YzZgFJEd3lh3eZU4r
39smpbatZiSFol/Iwr4bNluETevJ+sYsAvIoV5U6Lr/Qg+6GtSG4AU4zndFKadOnTH24clDzB0gJ
b2Ph4fwWIVMm2NGyk9etRqyc2xilxTkT8x/20lJQcVUUCd1o1vpF8SmjnJJa2vhpstXP7fhinlfN
CL6yBNh9K3CHenVI4Q7UnCSouWPZQ5+gPkoTdpYGc4R5CFOCVNcsSUzoszeORGy32nmn4UOT/6hb
iWOzgDtFaP08grM4M2yoSptz+00c65im3UEk1vuEVroH1smBmCfbgGwcEwxeVtZTTX3J4r9aGmSV
3ZikEvk4oCKCy3UXuq0la4Bdfh4WFTz2TWB/XlI7p946GARZCXSjYqxQ2PtAzy2VaE1wDHSlog7S
8VZV6eT6UgGfVcVFhHpY0qw2917MBPYqDVPjFUZh2CfzH+pOopDO6qvIqIgp6SwbzBU5P1fNgOeC
RtgZrIPBO1jkn1/VhY00NozcK9kQusM5hypcNTV7uKsnaDWOh3VDhonv7jveLBaEUAcdvDySROqW
daDrZE52QzhC8fEfzIc1baEW/1IsV9Uw/6so5z0NMWiS+e89ZhvYuKMmxdBMqtJN6toX7XmcyFg8
kgeuO8uZd0eaDyHyzdTDTUnfZVRlR+8Da1BLkUaSF+6emw/Ed1Qdm9wlaKqTbVlqW7b6MQiXLMG+
NNEG145hi3JK79sd1SR8xJXTMH6Us8HJXpXSkko9dG0uarmAET04sOnzS15Ebwqa1/I+N7i2N6bO
YIYJRiXGKKjDBtagmIHSkf6r6XvHHmZ/ube8VzjE/p15q2VdJwsJ6JbbUaWQQhdf0GPWRQy1bVDt
YrEFA6smxWE3qZyRAJUrG4myKYkxlzrQkuPRn0tUktr0IkqMAzDS4ojXgh+JW/Pb8lEq8L33c4wm
8awEnJMM3LVeGC1L/F/R0yklRTTfcIg4zM5eXtgRqGNMFanZkocoROvb19rsbRrg49T/etfOsCd3
tbjCulKfiKCcAeVX7Zk+H0pt78r4wCyBFE+aGH/1qXRijRVHchQ0cgqaAb3W1vx/xG2WIqfJQbsO
r1w+VF6mgUTytewN33Z8pRaRDUP2CmkIrK4K7oGyG45XVslOVqW6ttLWK8v6k4GfpUo8NjOwoh+q
CU1XvE4Pq29ojv0DjyIifZUbeBBU9OC87lCazlH3OOgt4yItdwLlf1x3XSAH9um8Haoz9yneOcXN
SJYM39hMGcJGqB3lkfwBkfgw8yPj1iMZCpnBzoltvyohUWbrA9Yy7XKgksWaPd+lQunlwP26spQj
0C6LsKfs/3J44L6UE8mgMoNFFt6XT1+lIlrI6fTNJ7TCgs8o87NjmTa2AsDR5euOlasMGceuv7Qz
GfqcCJ53Q6f+rLFSWC9qYF+1rlE1ko0TVS2p0/UwgDc3CUCBEvUEg99rzNkmzyGRnmjcBTfQjPNx
MybhgvMGlEGv3ynixOFf29M9NdXlq7j0o35gEM0lh/kJ3JBfSlnXWzwHmPiIg1OzO5nBCe8yxr28
3wScaZN1CbuIiNOc1OV3sQa/tN6U4qhq/w/Juig4jxo2g/cZRRd+3PFvME4QubKr4nuDTzojTnO6
v+nOpYBW0sD4wjib96kB7zLO2Iu1nHs6HATe8pkOMqFI+cSQJA8rdEKhFQIZRk8bz3RpFqsyNKD9
cy43zDvoKPTFNFZ6YwwBascBIj2V6W6dlMvXpO0NFLkwNcRIyI6CHWKE+Kt5yC91rLXsUbaPfuZ9
eyxGRfWT/HvJBuDmvFxQpg/pOpQuUMuHH9QgECPdzVYbG3K/nJtJjUAj06vtzSYN+IByYr7nu97l
xLzkGk3KpRpjl3MoKxyijRONhUpWkd4y7hU8lS9E2AzL2sA6znMJmKWyrLzBNb/WIktDQrJxXePE
etZTv4lD3g1yC+AdaMnwLLgiT268qILUjrpMumQAlBws0wkOaCok4vq/isDkAxi8kRZ3EOKa7hKV
BDv/t/8REN1+98HlWav03+u77JQQCdYFIa0QudYEdolX6kLVoogWes8B/cLpXvqZQKzgyQEpGXXk
Rn61dcfWO2w0h6WvYkoHbpHi8TMr+yq+2knKbDLb+PRVGvUdf6JZqSURfczxs8I64iptlQTljIO9
ovNgWUryd9jWyu107Hg1GTvgOrM8TVaNUimK63o1ohvLOtIdx9+OZrmWgu8NIL2jjnQWN/c0LdZZ
lSjU6r5PHuAljjaq3tAgBNrenfPe4GSdeA5svQv9nnu5FZCe9fnKjhjuhorWeS2GUaPr035RmZ6i
gj56+b+918CT6xahao4+xX21JOlA9y9oRSYgaQaiS+CmR+uPPuUfRYCap/Gp2qx/qy0d/VD/SFXY
CgMNdQoYftkiQ9Ylq2jMsRgjrjbCufpO+UnaDEtNPD4Bo2b+pIxrHvPxOr+TX9yhefmF1LlGjz6+
BY8r/ms/oA9Nno36dsLG5hx16LwiFT6zMdIcZaUjnIXaIufN9RwRm+EuZjzU0NoDvAzbdgFFYMf4
JtroxSTcjH7IJDv1Qohka6oFmA7X0v6rVsCOS5cYMkEmv1atpe1Y2L5fCQAhszj7rgKFGhl6Uh+a
5kJYgWhxEZoyB3Jv5kkoWs2dnr9fBlQtfEAgzuu3OiMTp1pZlnd8dDhVjti4b86mh7Tl1gwi9VxA
xONRcZ18ucrLRU/2yytH4zRZI3D3TG6T+yFHDNh5I1rOnIG4ayHHJqzOwGCVu9HpXoT6PMqJ7YwY
MVg8tzmv0ud0PoLQv11NcowQeKCxIWHwFLprXjKUZSTWpEGaYYv5WBgJR9d6DjB/HvKN6ua891Y8
sf464QNJ1oGCFkNdJKSQgrVca7A3tt3jec0thDrpwwpxSJ4MwmMrXnvUH9vMQScH03GgXjX0U1Hf
csDWAnm5sApOA+lX/KLZLdE1ROoacseZA8UR04zmQXUzwsJ7NPNhOUK7sWFFVPzShHb7SqYmw6dn
4XDgkG78bssRfYZ4nVsh7B6Q8TdP/V5++4XA9rJYQROGjWENb91fE4FaU39oppJMz4lyXp+2CJwR
LxhELIp3ZvA3+ayibESQoI5f6QJZA11lm2+WmmmLnvKzCJaNrnh2eK9xvlWBPK/pH8Y4Bf/QuNSI
Sc/pBSzmffQOqugxpMuymk3eTnQrZe20LtFxOnqUPEwZ7ESuomYypui7bILbOxMFTSO5Xt4FYrKy
88Jqsdwpka/HqUYdQx7ZVknarQLpAYK5l49jPrhA8Dvg+Rt+CwqEkFZMJfW3yT5N7JbXHwKH5nki
ay1YZxzWXTZawvyIF9bGfyFj08ChnXaLwWhIpcGa+2VRwYQ4+U2U6iIa5OicxMuWKzm7TN8sypUE
/3YEDFPcd0CrMoVidi6WImJ11Njr+9g5GNzsVPOc2irG9xEezGfb26XhXxINzK7hBI2H/r027+eQ
I0QNbLjBght281Dh2p2b6DEZvcAAsQRGpYPnffnsxlL7/I+CyTpi0wOG/pjlXagSPraW09m8ID/+
D+Lwpa4BwKmT4iz1DpSZARKhhWHwXB6dFfjziEYoaJRHNSsAps5gnYhsdVNea+/bmNpGO7lh6/ap
NWLjY2M9oQlJDoJeOpfUeIG7QCXurF4OFnKcdKJLzHTa1wvfq5kbF1RI4DvHsRCTusQgZfkTiXn/
LI/pz3nFPxEzoZs7w5jLN1jgUmhRIfOMQYMeOR7zmeG94CIqjh74e5KOtZkt7GS2lSKH/NXG89ci
ECFC5MtHGEMuUGmLc0Kr9Pu/8fUpK5kdhNlXT6sW3I44qdMD7Tt9xuoe1UMW7htfZByK1ipyE6WI
Z95mplaS0UFqBeGtJ+a3u6Rg0HPUTptn5bLIeEw0n7F4BwDXF6RP9OMwGLvOAyX0f+g0bLGMdLA1
7k0h6HJWlGw+k+g6A45YWlTa3f2tiGYLi4xvE+ElwnQ3WHiksB9gWEpxBigTNTVcpBI8ejY/QQv9
AsU6j9cIcAxQ4L2q0ww345TxePF5E9tflkUWTR7ej3x/Z0WbhTOy1SiOMadiTVgwHPqVqBp0X+Nj
41O1WOPVS6MXImrfVlRh+wFJwe271l68o0nUETcgr8Semx2Kyc1XjkB7n3/ENwOgS3/eWeC/TR1X
ZfFj6scO5fxukMin53taYwdWN3IsmJtf3/Fky5vyuzSEXarQZcUxImzHwCdjXSvSbdfHBmsb0iYX
CSlucYSdtrpLkBIaZPyFt3xFrX+MfSisihdbbbZmVzO8nWYpAXcQOF/tg1HowjVAQ24nDZA31Hv+
b8ZIZkuZScdTsM/huga7b1HcjTkBvHTbrpDUC208ERVU+KcoKkA6xXP6aZPzYbZLFz6X9IOmVeXr
zLYuSvfEO6NeoHf1ApE6RJGk2z1/dyMq/SXqPRPfp3rFazgAGzA2cuhME+PbK3yLfNe5mzWG9XXY
20CxmlULJ1YuWuW4QxXK7hTeMNK/0BgI+LMDn6aBhOp1NlFwRsMApHVAJpckcOUAalAyWDi/r/C9
16Ix+yQpYVt6Zznw2mq6hg6jN84D727qI++5qDBVrZB9H0YQk28KMOAgRmwzt73iWNK7iOi2rWl1
/VWxSYxrpzyrOxDfd/R6JF7rRFFG6As1m/0cuINR0wbX9twQ1imm8jRtxBRDz0x3KVHUljicCcSs
mNM5u4aIb/6reDPCaHBi9KHJ+YrmAkvZ0+Ug9cVV1JUEE+JwedLD/GKlOg67qQWJqR1vejAdKN9a
gAqdAg4lWDyB8JTi6qczT8tgpz0jRuZQKtUPKYxZ6XIPHhNWvAQzH4PTT8WJDj4g2JEq/DYCFWzD
johABSVee8P2i+9mxXlkkJvKuoXmOYnrNCi5r3IUJGarlOY7p+QHm3sucXqVnyrdPRJpNtEwUliJ
6TV1WfRayImE+JosemGbi/AWYeJDJUFVJ6T/wpW1I7a1rlugv1qsooUHjWtJzXY0ADyoCMLGp7C0
OV1kVFu4nIblRc0sJOy6Qtbi3D5rOwjeoGFfQp9dTOG1m2q8Ph6nIT2wqp78lxloC7DbhU6Kwea+
vvbsS69JkOh5m4BcWdSTvC8j1InJktzEQTx2Ws51O9tqOIWZ1FzEYAXHxNJlwowaI24tjgQTlfVK
qE1zYdFpbhjjVjzRkbIR1vo471zzBlgRJXv+qoCyK1mBR179eAlx1bZMuctD5sBoCq4KMT0NWt1r
sxoDkUJ4MPW3owfJgoTfcJtUQfZymTjmzeEsE8FY4diXMl1gCN09FfblZvNhpDNAv3zqBYIaDFhc
DvPO1e0wrLXKPDwP+ZCoBvKYKWQoaj1o7LfeECARVGAl+pIS5uBTckEp2FSlfcho0SkRbr9evF4+
tP8FZ3ZsAaLoQQoznU47ilULkrAlRTE3vidXB5cdfnmTacRleQxwgUaFrDyoVaLVWMrxz7N54yXt
wUFQedWMCGVad8+WViRmqjcxiby659KvesvxqmRaWF3Y8gQOLxBrHAnYFTl1MKcj4wWHB/8kZCxO
ySMCKsPQ3yyfrs+WJ3WPd9Ss8IO0p/4sxH1nr+KNk99IBXk5AFQg3KBHtZnMg9wsOwpehMJxUU6V
zljmwPYkrbpot7RW30Qtpwi6yHkmWOuIB9xhebNDLQsOJkSaMBGoGQm10UipEQsQrZ91a2TgLsKB
6NHFoVE9z/ddNDoaYOQaD+zCQDDtrvCSceCYS4+GCtZWQpfMUREhmcS3ZwSN0TCBDIk+fZ+/puv/
+WMfxkr9T+FWtFNDhqHe1KbAUZ0+DwcFCmquaI2dfTp+Z4VET4be+M+7qOhSE2At/ax/S5GRQKKI
r1srCN00dxDZdGklq0pRVeNdvALiwfLGfTynx1qrqI1qGLSsOLO1n+2WjLS75/bMDRnozq3QHKDV
zNs0GJc9m3ijFvti47UAb3MFp7zOykiAbxgXCN6X4girHJX2mPnKy0qI8DSU09Rv0+I9eP72VnDL
gpctwujJJ0Vac2za2REA2PxLCsu/LI1IVVJfRCI0UwQyULR9m1vAntUSAX4bEKlp9UFW1/XpamQd
NJUOQ0Jk6JswQrJ4s/eOL0ytxDIFZGLf2/oLRW5Te9zwDgr8VDi97s3f98Le+zIy1AUbPIn5de3C
DwqAOAOIctfdqgY5fZRY14+JkfFVdf8cAIvLrfq+IZSaK4OmS3HwQqyWe2HdWzK/3UU0ubmLbpSt
e6GWSyKEBghRMSZQtks+flFIqMpiSsXcGQvMKEJaau2RaiiX7VCnE+9OChuBcBDbl2sGHqaHUDgd
Xx2s2iq2wXaYbnknKfebm4DZq/L9+blAirscKyRhN+eusFWsh2brO5tOZCKEMWZCn6XgleIH9STJ
uaYUc2wBpjC6CSk7k0XVVLZHV9EnoKY7rVagTf6VS4gTSPXdzyAgRhV0QWATElpBkD+DnYSnDV5q
cadqNJ2f1nHUsZoV9wV8oZpF8aYgQvMvKLeN1N6s1nU8br9OmEuQxCqyBypWW4WDeEU30hm52gFx
csY+8XVtontQuFcPSeVTj0S4JQwW7MqXsfnXmabGJevAEdVlyPrM6CKmMj+8FnLjxTWRIz2g5bNx
1gipt7UR2Io1KqX0+aDe+ssSTy3QcMLW0LIFZkRkBZCPploEPzji2h0voJW7EKJS5/6Vu4XDcime
EDAr6XllMk8SscJy3x728VO/FCXBKcblu9s+dNI7Mqb3K5cJZ2U65zhpOtCL5E7kU//ZrM6mWRaM
CGkHVJFzwaavRVobbZ3W8i9ERO92NYIpnqrLHZlG0gcfcWY4oBY6frza0eXxx8lZuyVUa0xerlEB
PsEFS5hzz00iYyRkpLxXtVaAS4Jk8sVKhI1C2a9JTWKSaJx409I4rprUmMWvFsBBjhYoL8lq5qWx
iBi4+7xMT85JgI8r0eFUUZKDDG0kO8hdCGIRlWpraZpS+IkkhlzEFdzOtTtC9XZyP2ZGl1O0D5Hr
o8f59bB9oQ0Dk8hzun9Orrcy2A/6ugQ1p4YyEPn2i+RybG9NCgkl6wzEjvpj+AyyzCAF/1v13Rie
R+hwBFq7IuJYZ1h+LPjmVEusQK+4N6Is8wFjxZi+zTLQHLJ1TPH5h3KREA7MiOE1T7TGG7RmU4xv
uCQV87cHc/NejVocLQH1ByhdNmQoZRoIcNj0CXft9QaV/BNA+MbsDmXf036Trlz9Jib8DR9kcAfs
zUEyKVvJX7gz9iWpDKLxT8bnPJwavuJxJ2OBAXVtj5NsUgL8Oa3RhS1BjT3Au/oT/W5BULro29O2
x7m32yKnW2CDFthigDwMGtbkPrs8nrLNy2NBlsbdOyw5eA3RRzxCjPmvzGR2CCgpgg6s4xgQrRat
hqO64qMQ0OoXfK8mraeCF3BfvU94W7Nuz65b/8Ssi/hmC7sYg6pI2P8OLqIpBtanxLN1PwWTSKX/
fTNZPuOs/YH7ALROT6bStq7tveWOL2B0tFIf/tCmEIl/Js65zXSQllmRIXm9xG3R9qWoqznORIN7
zyisAFpctVqneeoU4dAi3xpg09PzEJYjDLOIp7mixzxCDuRo+rFnqm79xM2bhItfl/aiFMSOQl/P
v+QZqaA2ODnjg8+hr/qu9UlQ2EKky85Aq0THW94YBJq9mtYWXCwieT3UEuABy4Ylneqgo12002w1
/RPktHXB1zGCfvd7HSt8rR1KGVA4Ot7ExSKBmAqPXf+NkSKyurW4I5+9mtnx5/tc3vsFcpSxamFx
SDyF2dDdfXiKrdbbHl+ZxUWrDeaI82BTUI1tHfBMaM4SqrCE+//w47AuEj9s/YdsvjCqbqrE9mSO
9tJPc34Oz6nHOWy5KHTe3/dQwn4ijJCqkkJIWi6A2rCQFN6JeZIt0EtEMA0UVxo6f2wsZlL7Cgv5
QqvjVgoUzeg18UzIVmXm9Mh+8i+6Oln5LwygAoco/5cMTpCnJz8qdqxa6kuNt8Ydz/5FCMxtq5eR
KnB+31AKBcKAAkbnNoNQd0y+Qu8pxRzl5BPdVOo/OT0S1xmDBe+nkLSH3JoXjRp5WiKa5lRt4JJ7
p56Lj+C2cq6Pz4E8yoeNfyzpHactYlGTdZPYztkTzVfyvZALz0NWtb24MEnhEFDJMdySHcd9V8V8
iWLjYxc3y/WjR4SvDwNedWYhpVZZiaLSR+viB05qg1i1LyDQ5LHdETgbQ2+ZSFe3TvUNwGwC8Qso
UYOyAFcm3Ud33j00NSbj9H1eur688m/FFUoH+dyN91qcNoosdyogiKtQlsyt6s/ActcoR0O821Wx
dIocpB8ayn2Ux3F5ctJ0uotbfY+6Xi1Fr++nChWZWqBcDcBljC4/7QsHWHp6XCyCluHXCT78Hx2g
UDkzstLPeGwKdqXJPG6wjXfntoVYFz5nUNo6nWdfSFCVF+RIShBdfSfF9BRfZUUQusZGI56oQPvc
+YcP4T1Iy6vuE+pi7mFt8m34gRghIsXINb5ifoa2u8PunUtqTrr/HIezGj+vWOkv/vKjvn06Awci
XVCLj8TvpMpALhgcS3BhXh/2b+GuyvXCkS2G3GO/mjOspzQAbLHnfthniSrFfzEf+NI7YK+kldoC
TAvxy8cCf3ZA1zqQ8CnNQ9UkeW5XLDoHKuFafFNwvu3lnN16+yUcZ02BilhEigiJmbmAy0VbvWNU
DaQZCHRToZ7dOemERDpKFwEPm3yo2gFgDggei3Hufnnuncl2ULsfoLbzknaIUXnhM2wwxG1fVYL4
/AZW44iAH51nkFWUKJb2pqRwr/5TEoN42skyd3Q5SrxGiyPyYShaexLljPipFgD903WKcrMQvBog
yhcSK0C6WgkaTuA8PnE+RXBWoWWuW4SOsCF0pQgFq0uUBtz0IHLsT4sWLBhA6NPcLlyPTqS5Qe8l
Y7Z7ELpRWka0hobZUWJyDyU50ra/FU3M7xqghTOE0qNC921OArlfEfIMUSWPh2mw20LvSoD/EKot
D25sdFl2B78ri2cq7uItBthFOkwNuOCnQCZnmp96feryzWgXJtL5kG5sQGz6Vy+ZXPjp9eKPHT5O
8AQ7lSHKHvGZj51Od6lTJqwLgb35hvRwZ2kM0FWx9XjTaLb+BhGCswDzlu+hxuQ9NM+joj96IPGu
61uptsU7ajKL4qIJsJLuN4ENacz3m3t4jmcQG3aV315//apH3khPo+zjKXj2hYN0VxLgu22ZdhJn
x19NDqhdUXCXfxKk0kTrBfNNPsDIrEDXX4iTQBclkeC/dKtC+y6dPSGWxBdS2NBa5/wiFXIml5G0
lqoJ4P6y25Wg6fjrVdrDqa4ueMYUW5yThOypEfXkK8MMGPoHqGuDZGjnE4/guqQ3+VDgEXU3TvEI
nyQICgaund93LNbzTS7bEgph0XhzRnoDpJl2SmiJyil0kMeoyesSgKuLBAaumdWMFGrNmjjIxOgt
SDyj8MH4/BRlfzICDwr+QBBBWnWLSGPzut8ArYzYI2noXlcnHCjVXwyqs05Osdda7srHiG85OkTe
J/wK3VUD2uAKkHXFVuM50shFSBAi3xnqizgXAdnQg1pKfi2HYBE6fAWrijNkzLXMInynOLYXXuL5
gppzUYOypLSivoRBXcDwckckKg4sav4sA6pqrpkXh5IPuYgS0B9IgdvwQquZ3O3h95x92BhjMAMD
dieq3fxokWyIC2nAzBji7wiLuRlsd7QFYwFbYG5jMTdZl5TaP7hk5ez0GsxuAXcv37ds6A7+tCZN
6Kr8gizGRbZx/lGShJ7zgEULpbTBZvFHkfSFOTDT8NbazIvatkjPiusv4ulC4ZxivdtNeLPfhrWf
JaQiKj2lwSM/E2d18vcSnQgvsZ6lkWFQj59AxpppcGv9oiwcZuc/6FgoK7nrQuDfvY9OMNfDSv8z
kqnYPqdCQpQi0C9+p2tEYj8LCOj4nVE9L9M5p0N2idIqm3lilv1yLsAK2r8NKh+FZ6Cm770Jk2LP
n6wuxjFNpYv4PbWDhd6jqnF60WqgpF1K7mvb5fEwbJUsMK5IZ4ABNwu9lGgzeQU2NIKGQI/U02jb
fYtRXGE/Mv/vN8QjwpScRZLIsFWg/211Ut/jNHcZCpoD71SkMfJVOxlnD4GKmhO7I8G5p/ldKoqr
gdXjyJPfsi3B4KtOBoxVEAbKkOck0HCiEbtanKWN5vFJvy4RbBBa20TzgKe1uUta/OEqXEVkNzpX
ey0o3Pyc2VP5PsZVU+uW8zhd/5KQ3eXoDuo07TgVsBmBfSr9CHVC+Hf/3IQbA2u/XV7Y3tfESiak
8C3s2OM55mhhh8aTXmStGtYeRPZhdnA7hWeWYKANDgV0htuYNuN3grNbz4MrRWVrJ5gK1lDLmInt
T9y4YPji3ZKYxm6syv0IaWIkfw9J84rkaGbLurXftaG6XufrpwAVzSSd5MbE8NsdM3xWJCxELLl0
JOSRcoOfadpchjsPVw4LDOxSFftpv7yTlPyO75aUW/GO+SwmBPlpCny+Y8UKAJ+hwbrBLScEi1O5
z3YzILsMBrrvw8N/41aIWIqyk6TjkYj9VBv5/sZEr2CgcEMP0eeNzp4j87fQbMPhQar3IqS/foEd
BkJQGQE4NRkMTC6pxowSrynyoE8J4xclMMmCkNNP2zIjUV0k9f0ueJcaGGOGrR+1X5zRurYJfPOS
ACUFxxlFqiRuGYzPTZOEi01eTgDMGGMDz8IWdHJLn8xv00NZy2UlPvJeFdQMj2h/HOjfJPl/Viqy
JM9EQRCKthu5kitehJnUJKAWKcb+zHE78BjJ5fwYX7fJX3Bb4Xy/vjZ6O12qx90X+U8q0DWQ5dr5
Ow9VvTDwG7BfSrqrhqQnV5AwMTTMYgxhsSuNEMI1wk49eaiChSPVyahhXkJyIegebHyWmRSsqAun
tpcKgfwI9SatGyVxFCO1Arro/FVkhpawpgqV9IYWUnfzFrg1Tjwzrdh0zAufiX5Rys4+ZnkZzldH
9jkBBfK5TGaaS+qtVhf+0UWXo1gqlzYwpfcEU/RTqwUKUE/F6YOa1QEw0eFcHWflLQ8u3RBw5Q2m
yJN4o0FCpulFA3geUEhw0bXmWxgfpJncz66ueNywZyVds8vPsPWYJqlZEa7iKbECpc1ku2vc0kY0
JjZ9EdghTgjYNtzB9Iq1FjsUw8yVUf+L+XqYc59z+mw3xNjf/UbeyeFdLe690JcWaPDqTPDw9T/8
c0p2zFV6m62GpMH7+9Hf+PSoP94o1rVBQKhKPEBAjU4lNZVJ4GrgalZIld5vwhfGTF1vZ4vB5HTj
AHfoDMHy6m4dwY+CX5MoZ3W6NlMsBqSVLD+LWOjYEDFAmMA0tV5eO5yjmqwry13PPAP1Zd4qBhZa
MZvL/TEEjebbwFLmdcM0vt8fqLGWdYx21opwXifjjVSnFp+3t1b1k/W6yWtqpsQzm4MyqLHHCH2H
2COWHzSrXrCAILwRZt+XGR44Yj24ZawbmsOIrOs3yr6GhilIKyj0+csVX1Kdyr4UqphdjemYtE/X
8BoJ2NRM5NqvFVSDnlGyRGl3jS5Ll1HpCTRqgHmEHjOUqmRZX7ecg6dhr/XXJvo9d5MIvrlOiA0y
UIMjoSV9GMU2bzOZx81kdztprSYzpPgZefHr/yWSuCUWH0M9+IuGxq0gM+NF0bN6AoPLhkD+HL57
UnUuWrIEANltPfTiY3TtFSa4CFVfo0IFl7moVNrY95kyP6paGziTf+ZbcRq9PRvbnPck8+zheCKL
zIuYs6aQUV0tKXcXw0bNSytcEvyfNOVdEcU/gy68uLrf8ekzUTZ7g/P5L64OSYtlY80c0eSuWJiH
NlQLRYUoJRGNr4TNrste1B2Kp8ZxfrKMPIDNVVeGn6PU0jRwizeTSvLPffGU0Rpn/c9vJGlEcg1V
uGEoFkosOfvBwU6hVqPsyAC0PDWzb7bDD3knGb1VhPCbs5dixbZbgODB8+hIPc+Ea9GZuz5yvZW9
zG42Cot8k1B42p9nOKYM5HVBBGdmmxYd9ZLDNJUNj5gApHR7sczjThpTX4GZvS2GjESQ5JhpOppA
hnhf9+FM+1VRntf5pn1QScVvGOWppyMq4gO3IB0YbAcMj35sJgMqmQEC+DOJE936nK4mp1l3yCfy
0IOZyU3dlktL7EvyIjLuqoVO7w5KwKOdqWsbJH4J8FpyHfYja0FdTEvWcV8ZR+QDnOcagdq1vpJX
0JjYA7OGeLwQG0ryQobb/WVGGTZZ+Y0pL3PneIRa313DXHe3INNHlTRs9oF384EFhm0zc6pZBk4l
XZYGiglJZVeEoWZEDj4zflliXnYapuvtwP+Me5EEQMZIgUgnLzzCJ3opInK0ySGO7xZnpGZQiXOn
M6SN+imE2AAJ5iX2Sg5eUmiyyRpZaV56/mMosxbxgIHvH9n8QvrARa2OK9WVa/x6S/Bp64RPMj4D
wv6tvNL5b9PlnywXzO1kJG7nFW9/gmwlsQ3hYKoYv6XynrSZjpNw/8XMucIAUiXtjNiPuq6wQQ9P
V6BqlcD8yQaDgBLcm8dsVLAU/MGAi6MmdkUP8NmDAS/c+lM9qmODEvA89rMSyh6ObuV4MQyAKdBX
OZp2scbKBQpajuBLBrQQYnEmbdvsHIN5m0ZUQIUIYSBT0YVonSTpJFOvABpYVIrwfKyyX58f4EzC
zNBPuc9F4Z6B0BJFFKA0PlgFFxn4qp+kRjXfCqC1t2Wn+TTajVjjpAhQBvRa4nzkj78gfWdQokcR
lS5v3kAMBot5/trbvAeDH8HlRhqa9dOrFICU49BHhrLpPHrx9S6QeJsW7iL+D3ZijsTDErYur+WS
63mjuJzF0sx8T+R4hcCTBWyxa31wqGa2lHNvuAdO5VhBXeYGjKKV+dKNxhdOPAiy/sIMWVUuXQVI
ifKCcGm3+TICjMui3/eUbM7JmmLEa1cAAhouDWhZOALcQaUjGXMVhJ/6ulwqgKLBx4plebyPjkxi
hNKsH4GjaCGT/nmGu5OhWWa061eF46G1r/QyRFLHHELfHSIUwMRAHojuGvnRCg8+Bs8Lu//s/aw3
jSUsatnKvbTXgNFqIRuFKBTJ29fzPt3O9wMXme8MmlYEmr4+VCypICHszOhb2I0ChV1SqoJahGYR
Zf/O/Xty4av7S/HJo1PpwH8R26bLfWHF95EbPiyx7x8tZiBfZL+oWpPYYdqgEgkIp+NU1PbHzrfH
PEjK/6pMG1xveHDdFwb/eMFaPS5boufe1v/IqIwZfhfNoUI9ANOM8v/aC2SaKDkA8hw8SRivArkE
PVTyunCWeB1bj4aT3XvRONhA6k/Z3Mg0zl3yLM2OQIRwWeQ1b8HeGKH8hMsCFbBwsG04NDJcQENZ
TdKc6krrE7T37uyCt6jrepkJOXBj4z+AKb6B5nAG8wzhf1gfYrXrdFZwZPP/ojRhEPbj2NNEfB7V
oiwlXHWr9FKn6I6XRa/54g2PtqN2KIH1brNScx+uyfhiBhRlEZb/LUkPixdMl9Mn9XujwEj1d4AU
7OYPS7e4qg4WbKinJQVCmhoFxJiWAMUiJsE0t9DPAikRZp2P0wxIEX+WWpVkY2M1Se4ODBEBeeKl
cAdpUoC/vufpKFqee3L2aH0TI384SRqSZZQLSKOLwUHz4YvBysQPTm0lwgk9JxfoHIZY83FpAM1Z
B1CJT6UJjjoQo7XCpFPRTzQcvJDs2MXvxH+i6W6eb5gxJoXzgQmKnavqSu75apvog8O9jbNCNUKI
Ff+3CGfZoJQjr9sYRHDPjK/q0fAYkVf2WhgH/C9nRbrVT4RWp68dfALFNhT08eJIkfh2+mDNkxAZ
zbIheE9OJhgiar6mKAKWo3a/vJ6QnSnZygmjLkcKXZl+ysd5fycWrPsoQiCj86ENlb5Cmqu6Gln7
xRIyvlznxkgcWsuIUOuUKj4HktbhS7ULEBrK0gck5GPDvtz+yCsLA8s0n3l7v4ZB1ggiVkX1Z7/P
BblzCE38ypq31xsB9W8VARpG1EblOsqcIW1CJpqg5sJuSVujnvGNSgRy/Yw70bGfMwJUmKa/ArH8
C1r+iPAzW9x/mFzYrbb6wSvLpwpeHTUZA7bLF2PzJoOmBpHxTF8CQovGQF5pBtc+af5LyBgLks2G
q2dS825NNucP5AIYDT9ck3D9NJX9hP3FvFw+V303JYGVaUj3tGxmBci3of1G9xz+pKn8bo4fqpNe
Eo/UoGe4gyG5v+996a3mDWviu2qKYhNL3Ie2j1xpaMQXGSag4fdQttb23iJ/4T+F2JBk4zgBF7Fg
Uf4blNNbu+k5t6ncfpnL4+8mVnMpLkxHnLDmgB2A9Kmom61ZmcGQJTdI8KVn0IVh2wKeYZxGDkob
FcZHq1XzzSFXIQo2qSF2iMB2xgJOY3nCoYmgWbLYD8canObTIFZE8+RawqEDuy/kyq+NIPfQXxsZ
NQUfneAbjED7/LRjVA0mo2GA51B252pp5ZM3V/ZvvsjrSi0WBDdVOTqY6dXXbPR7YqIkjuUKTEq+
440JnCeUWd9JSMC+braTKhgBxypw9uFqKfebxcQw7KdhPcxpwoOK9O5/Tjd4GdaGVw7dhxf34Bo9
oIRfx99cS9AveOWEu89p+zx6cXNu8+KVoL09WZsX8ntY/PB5ajhlzXj0pFh3RWKgTkvwCtZCack1
O9FSzmzG/zDNWAzOmKwekwb80JaKvdguIp9tVXAZPtJ5I415VKxBEE0zGof0El2nwkDWG4sQQLbb
kNkcwzfiJdCqxidRbKunjXjQwIXuKy5ojHjsKIDgTdsy5HsFpGEMJUBdtejip3QoOX6v9GJWnF/q
o6FxlRKNoSHwn4an7qsrvJ/+RnRi/MG+xnPddyxpiUYhyHAYDzHhROc7WMfFxt54gSXBAxwGbfY2
9bucw3qWAEVr4p/HkSjHAN75rn0QrOu7csA92n1H7Una71qePQk8NtCXYPt/zHIJEoy6WIYF68Ld
BU21codsexHSezH8p2pcPwRCIpWEml3COYMHaAnX3UWp4+Apeg1tovrRWoXATJw7z10k/8omx1EK
OiMC4J0bwUwbhlP8mlk+bBJligU+6wA4p+wxSKnQ9Kn7gPQt1y5SniGBWUa1dhQStMUq5Nu2RT8T
XiT0P1l/a2C7vWksMa4Eb1GbCnpb5f2HF/OnZW8HvypShd8pbX63fbgB5YQTi1NoSpU4DlRvelbd
VG6wY3OCGs0+vYsyqbB532Mv5nAb5gbo2OgLRLtOZdz7Z1z5hwu7CDkh/5ZnPfnCf45pjynKNWRG
p/bD3DNcilLkLhhdfpMkWn0Fnw1NrCI1D48Vanwk37Tw0FTNiq0NEyfF4UqmEDEvoPZn98LBC2UF
cbNVHv2N6LqFsaZ9S0m2ccj2maDAfVKp8+ReP6PKrwPOtKhlUA/xnGOZhaka/AtZ3djRW2aRMLxm
CHlvMgvZvxX1DuYwd96dBcgJ92tPVbN5l6T73Fr3/FyB4GIpYmCAEtt0BwmCN7tC8CxTmYQvlECM
iYmRlsKxU32pZjUp8O0A87wxnjY7pgGLILs58coiuTOSR7jQ2JT0WJk2tCrWliZ8suuU1R8F9M+V
fkl9cXtrX4v9i8Tr3GKZY69JzdYBY1GJ6ZunvVxhgiT6bhd4nC9xClXpqSwLoGEc73ESSxE/9uJI
7ZP1rHG9uwr/qIcUcr57aUceDMocm/XTrjsfi098oBGTEO9slKata9DlTx6g/nOlvHikSD7lEBlE
JEoKUQmkzIEIFou68kugqZOF4xhdk8lpl2LJ2ypCb8dLNJpyhZ7lFNkCg+vVM4TkaNPVvoFVO8fR
hIzRG6gy6uDct2sIA8lN8ar83VAYYA2S9iR1SywetJg4lKZ3SabwB83wmAoLOuuwcdvQMqPUnqMi
ZwDhww54FgQblsJD+iPlbwj+0ZNiS74pW/i4rBXmuLDkI3fBFvlHRd0XMWop59JNNA7r7c02BW/k
MjDpA3hvUJuREOXA7xvy2MgytjAx2jyKYITJ3mh4kR9zSp1wgDUJ1TF8XMABAmhm19P7Rze410Wd
4PvDwNtq/E8IHjpoengfJYIJNVj2bnsQy7V4OVTNe6fwqLxkF5NxAfYIOqBTKscWEvKW8ngk45vG
jFA0QB/GnBFbp3ybXqFNyTRUMO421G/JBQLyPNrWPqNl741HFF3dW4ZS8/UqSPZIIwhwTHY1BLYW
kT3L67eT3hMf+F3O/V+UKEhxNCCIvNdwKVTs45uZmt6cmOsiiV4wQgOEkIBCAMK1xPF6ISCcGp+5
dl5gbuTSCVWjmqrUVttn1XBWDWLu0kgTe9a4yvKktsritZt5DI8ZjYjTbMlqosLk1UeEzjSIgohc
Wm1jCgPClZY23egxIxVvx1zXYv4IAoyO2usdj73WSOVxCSYh5DPMuesvzLszY7FRTBZmnnkLOHDC
nDnifU+KPzIg6sJg/+ozUZVIIS42H2SzYKKY7sjJ0a4Pz5G8vqDlcxP7cEPUpDjJUk8ND8hTjQp2
vVKmE+mNV/VBJhu65OVOuPGPHzjrl+8GLy/oODY0SUmsp0nXaKCkFmrFIB5G58+me8tdx1pEDfHP
516voWB//SWe3eMyRzZQ9beUIhNSN/zXKitfu5KnRzh/thd0iHfLC8l2HpQ+79rOZbfW04QDL4tD
9HvzQgFQYa1AXOiCbQ8QGLlPIKHjjtzTPZpo/zdKafDa4HQT6PUJgH322k5b0cgiFJJpm7impTYd
M5QyAWojoEXVwKUPnpTO/p6wxdJbO9Hl12AYAav+T3gQ9qXlkfXeLxWC0iEGmrLH4/CxQYTCFry4
HmGUzNB7itDy8T+aiHLdlodrfR2Ezyl6OILHwMu78Tz5N3y3kBsFQKyN6Lrc/s/lcVQLEfUpEj1Y
QE/Wj8OAmwBeR8u34O80SPpMbTRBX4git/i/1MhXngPVXo1l0Uv4UFfBILtOUGW2MV7/brnbQeD1
c1ieRVEKEu3n7/271g2J69pdeAXcZV0I6Ij1dvdV0NrhfMTVHNox5tB8E0ZPSakyDwB8QJHJEMU4
jZ9uuwUGWdaowS2eColAC1cOdRp0OjuSBQHpcm6qNszCu8lC0CzEfXou2rUuZNRMGHtyyHBIh0UM
ZUYUtmvugNhnJxElEHDdBBGWI+sWM9yRtZCy25pjGuag6BMVLVynfrisHV1qA3HCLRSb76GXRqtm
NmSoJngyh+2jmgzMoVPIE8ciJSfa7dMDKr1uzdRnVglfKYDWQs1md5pJLFaySeVpgqDnkdIHFMVt
kAf22ZZdnOtp/1gVKrJuU+fHS0eSWNwaGbQHdAqanMApVXvu0jP+lahwHcC88OrTDZF3C3yJQtpm
U+PJDx3bsI9rQvqCRjPn9auGbZ6fpBlh98Rvobb3F06E1vhMcO3Oekbi5P3+aEZFBJTzwxHKAZj9
ETebLkqPgPHcea0czwKsR3CiwyDT+4XC8lyP1RZR9dqjehtcWb7siXlFC467wX+ug8D5isu3Siz6
pYO/MTtK5U8smfZhn8ySYaCuRPegMGAhAecTUFcPkXzi3scMHMwS3EhvsHDEc70Jtz8DFq44+mJP
XwvkhyhjNfmNSBMsiBW3zeNVlcyi8JU2vPZiKnUGw80l5nEnDGsdYpp7nlzIFiRp3RECY0R76TXk
TqpVjRLznPa9zxFBzEiZJE8IuTTKmhOr/ssAUzaCcGpLvaohOlex3rhTb5Pp3e+3Y/7ci7VAvoQL
IVD7OJuTorgzTybblgAXg5Kl5m6DsNepwMOE46vC12Q5A7BoC0CxL1PeDJixl/SuiujrHlMqCG+Y
RDgFtqEXkF52jIxGMmdE3vypZic+9mmNwV+iVgTbLS39xzzeVsgTAoKB5azHN6EMVGfb8FS6Kxa6
wZjUO26bq1ziQl78LiILmsQnXQSc8NSh4II3/5LyHMNqseZ31CE9S12gWtbndGrnKaJB3mBSMBw0
AKHTHld7fplWnB68J4GZH87zQG+xdqePJKHoVFtIUezx2x2F6Qzq/zYUBVbjopdmC6OpUNu1pWa+
m0MCjq4cQmtqhclGCMrhvAz8hzM/F2maP9DdOMbYnMAbp5Ezw/7Zd2aigxj0Bb2GFY5k/QLsmCki
khPkWYPP2BtUByjhV8XJUF/rOyuzA9iIEmyLdYV1+KS5uCOimxLap3kIywxqXvz3qTKCi7F/l5H+
4lPfWdG103ai8mTAaHcho8PaLNomnZdOYEj92tUQDvbGLyHQ4hlN5BMETF+H5wJ9cVJAycP4NcrL
9Q6NlxluwC3al40cujGApExtBs76cJRZ7DwKRe9v75NQaU3n6eNJn2UBldSILmVrNXPUM9Lgy/yQ
MMK9m+mwngery+mYxpKaaevsJgTCiSU41KD6BXi3ewieCtJCcLlAEmQrZUcOVQYXF7AEB6mB5XQx
txPraeR66MNOAVykZg7kCRn1lqcGYLYNpZObl2oTlOStOlxITFW+MoTs5BL6ulsA4UFF+4pqyxNY
fewtR3Obnab/sltbFNS3vQImDx7WR9a7okh2X/TeGUylSbns4WlfAY/YW8clYldO6vIF4pUCwzTK
zrFmlSGwWMu57YY3I6HEss9y/C0vw6Pizltsqhsy2JK/HUxx/vspoigLDvrW3jUYx/kmq6lw11z1
1b6BCQ56NbnJ4HngtqNJtyC1Pi29LGGhDDrwyMOGUbec0F+0L1TTunPYHRvcTBtFL0UxR4QuVJJG
f1SL4s3f73ZZbOfDxQ141V5twlAANNrasFIftJepOuxdC5sCc6sX8xooNAlAAiIKyf1FAQli09MI
DYiHtlvX//PADuuEFi5PZ3UHdw1zsoSP3TmzzkQU/G6DhpAdl2eatYkMcqBOXg75uwvFzDnpa3eJ
ecRRkNa0vvkBNyjrqvzC9SFevFsQVX0syabFMjBPt/MzVCDbofkQD8cvSH7IXvClfLJwrvnA6DHM
oxg8ey1xWrOOT75EXGNqxXTbGKJCpQEEghtFyMTU8/YUrg64FonkQcIX6JnYn/mxa+W9dpXYntnF
8N0K/CKRuiXn7niPfvrbwD6o/RtrJltu2t9VVq+OVfcNrlImAut7JE/a8Vt3it+k6i2evIAp9PoE
99vSmUcv81GgL8wL8LoOeDrKQZME1pHtjnQ9DnZbGqFYwrGDXW7OG1fw8kT4s7FZsnqXWDkAJWKn
cGW4oKlr42KpVCy+W/cA3EBydjuE9CIQLvxgkd/Mcf3qakcT0Y6EEvtTPiw4TXK5fky3uP1mLBXH
p/5cjgko15okKXYelgET6A3eocyY3I1pqlJUhM/GUBxgC8WXt7DcoMhMPiuwoyMuB0CiZ8gNDVLh
3Ei0c6hcnRq3M/GWVR5E/MvsPZxm//hd8IoYjY3wMXFbCNx+FAelr7Nt07UAoYQuXyYk4k5IfshX
btTcO6+bBhwLe3VSDVI8dMO4idT7Jx+YXAjzUHptz8vrCqdtORdzXeoHVZC03PQDJokZ3zH/aMEN
YwlqXqh1yDZ/qEeftp1EKfNLdErRI1qfUd3sXkfrgHOGX3Dv0SfFIvr9/4Y1JbsCD2Zfz477P+Om
j55UTCEhoVbjM0hULhS8V6TRefXnY7BG3Z6yTTaGA25qg9T1/zReIbVv7MGboGYe/wgBEtPnUkDZ
u5Ux02zTfGpl2crNwg7w6yRcL9DhrkDaa08wwayhTwY4Wr8b3akEDwX3lZtmJnHjRnelFS2ww49v
fwimD/7CZ4rrwiAn51BpdTI0heQWPj9tn4fuVROhrlyu9KW8AVzS0ZGqbzTBr/KK36JYX6WQcosy
4ZcjNMvK6YribcJQgEDHy9wBLH6LThsY0SM3FvWQk13jGeYpABRAaNIW0LrY1KjjB4IdjQK4N+CG
1z/MOxrNNGUmuyFJeJSDOtgdhnMrvdK3pJn9v3nPZ32s+HgZxq+gRSfT669kGFiRXgCgrT7v6NSt
T94w1M+XWr1AbNZQESEqFIB56CQ6m9N1VrlbX0QQb6llbfi1ZVllqE3SkUKJQ/0eN3/Oujid1Q/b
IF9vqlCQZiw/Ft2Y7SkOqdsDJg4vYO7aM8RnpNDawucAdcYNFt4Fi+3BCYi8uILvjBCX9pLvhF96
HPG0hgq8gs4u7KFJoynwUofUIdNJoP/VlBA484Blz7fjDmk170ymKhBFobjNz+9XsKNw4co/BNkH
Zbx7/LwG/VtcHVnEGjS4BeuuANWh2tNqq/HJFL5LAgpBrAa0rh3C07SjCXy5sGCie84X7lO7x0FF
nxgK1WHOkkn/VuCGx0IZzsFTZyE39U0dIJQ7ZfO5sOdS8PTkD7TIm5cPCujbYOMKXUbnAHh4OJ4O
6NB7V/RpAlvE/8SLYKD/obDPrGkOGf70e61AlOb8KpMvRztZH82Dx3zgqoHLAPhE8rySOi8WX8Nn
HtTS4+Rfbaiqose3FDjKbq7m9HBmSYE93RHFAiXChtDvKIoX0mDccCOu5P87oSLN7CBlfU4RJPr1
K23Tvytb2WfC2qGr1LgI7H+VbaA2/TWauYxUTueUuXuzab6zdzeH9eN3dN86Ftcn1HZRjl4hkJPv
FgkMi04IzaI/Tj1rezwGNsns4T045aBDFm/UuUPFlee98lpWG+bJ/FDwsqfgaNclNuyQoDNKhTf/
6jK55Yv29YB4a+1IRv5aper82SnR8cfuOYxkJRxcA/pu+F6ekukOLwPeiK7DGQ8YPdyzN/vM0SjK
T8hPfkx40jMJNvP+JAy3o/HhgsdGz1wLNA9zqpeafrX1OWSofCxIYrzgXxOnIfGXJNg6soniQ1T4
I9Cbpyj9N2LQvyimlPXcO7jwpyGJ95vduz4KEbG+eAbXr70o4wEhjgwk9C/TdhsSpxfHwmjhZ1Mq
XCI5ZU1HhI/lQRwDSx9ZMz7N+V7JnxT8TtV9323N/DkKKB2bMG6UFUdoTpmQpEVGwUb8C6ub3FE3
f9Qt1Qp/zUbDJIq/wD1KkB6EohG6e/T5Y5n7LsoUypwPF4ChNiImA/1sONS1VaDdeAHKn3BwCfie
9w12/2EdN2LDjus2RlBrRQsslaNx65VsATI2dBf4JiCKtGf323aZh0KZtOi1Kx3D8CSyZLKJbvx+
4208oY97CdrCJWYgw0eNFS7ZnQVZdwGmh6jtSIoD/efHr7ht0ox2IB2l5xKuKFYBR+EA/pp7Dv2z
T1hbG67/LRzppM9V+ASNuD/c8LQe4/d12RYat6ySCoJB98+bYv49sq3Re9F4ftqa3BfIywH0F6D4
71JpQRHeWGKuiOaZYnipbYWDM36IThmLv6lMrpQoPF3L/UG1HF7WUfqFwLtPQBClT7ynqFOe1VI3
nqZcxnXr/FndrJMyohgF6iHRBqmd6K811594CtyYMzTDSvxz5LGUPCJqrEPk4luUGqWlhg4oBnKv
x3/N80a4RQpWCL8KJbCxj/GOQU/vxU890NjRogUaFzRiMBd3Bo1NZoQe+lOtv2/fobAMZ7I06o9P
pjdRVcoIkElkPBGCkQhA22D+tDWqOyBoLg21in4uGu4nuYulqI0HxWsbfG4PLkagYtInhKU+ouAX
9Xu/RmX3Utz2wyCmQhsUtTvmbEd8z6E0rC6XyNwInHmRO1NOcPwIcJtgXoadg+w0Ffo0drjcyt9p
PldR1uUEhaf5jtZdLbAIyMxkSVez+9OKuDhIfL/oGX1x7+RyysY9WUQ7HTq9wVqv7tEr/DItzrri
0IkrGs9RhQLprngLxVfHp06InGi2/PZlJhGxFPqh4sCnqwekGLr9PBWKEQ4iHYtxooumZgw2aV4R
8xvfAwvrvNQIRNaYlKANr9IBNG3b2mcqlUpeGlxDmPhpAlEc2UcoVubULJyi1sUpxAAra1SIck3a
eI0w7AHlYI+Ol33ze6z2Jh7/qSDtBU/AOdRqDu37WnWVT+CUAfNxP/SFenpTSusegjNTc8BbGp3O
Yt+W7kuhhLNOKbuzzGXz0DS+gprMQKA4BD+9bN7yvIkwB0EIQrgly0USHT71QSr6mgo/vjx8nG5x
QruRk1cKgCDvtuE7fEYX3BOZnzdDc4dklskdDwpP5B3lHwVjglvoFSB/ZrEi23O/dPqecZ+pTiSE
B5xij+g7jlHekJzndr6AGKYY3nnIVunvtdCS8YX+h6i+DDD/hUaar0X/6WsSk8kHxyoDSHIzDeW8
3DjD5Ip7P/mpUOu9SghRYMbuUMw+w3wbdC1FpCnfkalys80pPFAMsHR9PTVYcLWrsxeS/CKIcFa+
/hrLoHc8mm6uaKyG3T8BPct7cIi/R2Rt3P9S9igwvB5xZtwtgxos3yOhgHPij7JGJ4Ps754j0vo1
mTTGNzQ0fF2LRSAO1OxShw+5/vlkNVNlk0+8sqPG7JH815bSBtYSLKTloixLkVZfoCYiTR1MwkH3
cJvfVqzsCuzvYsY5sJiFRPdlY9IbzcDsxC3pk8Ko9876uCVGScOkEghbJBc2CdC0pa3yu4hjVvPN
Qnk12YlV0yaNaJ1KwiIoJVqr9AGVExGm2yJQ0FbH7C66XYMc9usLRx7PVwdkHp0idl9SdH114c5r
gJeSo36CUV2RpaReOnwRYtNaB1MPjKmwGXn2QVGw9DUjdAFBPaEwpv6FqJlfelPFT1hGGNaTFcKJ
BkWjtiB5luGPTmohPdbCSNiljbJxHYkbbY1APpPJ8pz+i7DQmEgRL7xz9hHdQS7hQTmhC3zbieFK
Lx1qoZjvBZrOkws8x29e20NXUhEu/Ry3RmXgUBEbW93m8veKJFYqCG3FA/F1403jXc2/6MJcCOjb
sDSk8ptVxBTGz55Zd1LN5SX8hWG3Ds+hHm77W66jzTb58vPmzAUHxKkKzmi+JRrlDQBm6MHD9HKc
QOtMhQUuqx/Avq18ex+9zdw0U4HkGeYhKV47mS2m3Bmsrhdvk2Yyt8++pypTW8yfmN8aSyIghPXX
o194EP1WRo11QU3+/wDnMlFiu1d+iJs6DplaFdxQ5c340c9SwcgmJ0/m5+pH6mb0FR7HYb9Xpk2C
Tb7XWeZ/FoZHzwlyylUXxGjD1TpiAGHLTdOc4Me+RAbbmfRK8CjuVaBSEje0uRArzhfuL50iP+Lw
IDC34hlkQkNlLuR8lFuSH4uxBMbkSSCp1XcF2zJ2k4J/Tha4u/h8JnI2PuhAhNkwjR6NRxHmAYJg
cZfFUTtzXiJ7lRYWoE8FqYNrXndBYXPUjgzLlkYcWP1wTrwU8M8j2h7sDKKCuzypxsPtzZxZaWUT
ah3qa1wAk3HosbywZuCIqUnrs3fh1L8Fpt9ESb2kZfzs+5PiX4Alets8Zen1bJDsUzk1PD+RvZsv
e1KN9sG+jsXOjV7fBMclKoZ7hZMgDve7SX/PR86xmHLnDWXsoAhdRihs8rlZR8JI1kGxxCnmqy+F
xuavPtM7bx+S6Bnca1pQh9aC2iPAqgq6MlOmEwx0La4hoYAxUdvoSEXgYz/kZiaafA6NL3DLt7zv
tBc/dqrm4DJAZ4gmXQe8Dsvpc2DEfjboKuHOHO1bsxdxtXiIEsoF2rVyJH+x9qRZw5BwFrZZvGUU
CCWyyZDU+3bjxH0kNT2YhhqLrsZJvtzrrM3Wqc8mkKifyPptZcgpzfqB621wcQEwXaQJsQJuOy72
Vinh2/ABPhuwHI8aJUuuCLrmqy0PCSpgW3YXDkPPs2wVzvmDZTXaZngt1LtwL/AUZpMvp81LFtHp
TKo2O/KCOfSj47Xw5jfv+LyHqm2BL29JzoQAvw0XWmg6OOhj82fQdLHbxu6zSJTGbibwYFD/UPaL
ImccqvSfAxSlbC1jg3T5WfEe1RU1sXYpPK3I8gL1vIdvIZVoHs4Msi7cUxhIGZTZ2dOTRM6C9l3x
6RFjl+u/Wp152opLe2nnJ1QVrX0NvC02qaEQABqEtkOzWtmbPgS5llWsq5hfpxW9G/UxZYfyjoUL
+NRW1/GTeOWI4hS87yZ1gnuSMZiX4VE6r5FKdodGUGZ86/66NbbNkROaPKg+O4Z97xoGfn6Wa+dP
KDRW5uWDqgWvJANLpEyXfF3Y7DIvUXYzs5BT6K25lUf2CHn2yboTWodST96Lj50y35KDXeZ6y1RB
nZiStECXk4rOJlTum2FbRfMvARokcxteU831aIgwgPHtkIh/ui1Xt7jbbyUO1B2XtcWHG3he2JUj
g/GYuvbCO+JI5voN6lTnIo0b4BgqqvM4IxeCHlp8kJP6ZEmjZtp9rt9yCPe7cM3Gw7xMQRKX6p1L
Efqbtn128EqOF5zPyl73whRxH44hYTdQ3cQ5T0IP0KicBmX2m/C7rmsVPcXsjDeMerDiZw+XNFuh
Nsw9/TTItwmWJV0skD+k/hLlZ7pma4W6FSeOu8oLM2Em5HR6x6SWVIfe99P6wrEvgR5e4/aRBjnW
O1xzwxTxl8OGpnCCGosN0XoTeKy1rHPLlzsBZVt96/LcPg8/WoEqhnjUFuARzPZzk5T0yl0aylC6
SMmA6D4deIV9GRh9udKYlpqjyVEgIQKzM40s8aKGdpV9bdo8DDcZ4T6MvqTAHTESHAXQPw8Bhk2n
qDryt0rw0WPxw3lSsmtQG2SiX+OZaaCMNunSZKnypkdwuIxRZdKLk9vdH+vA+PSFt70QWzBkg5LX
SsAirPttVClHpp1zdAE9rW6cleztEEIvDpiH2H4Vc7919+/TITTinSc/LDgkUKanNmOW4af6jy93
Gw9JubUZQPx5d/7/oINDG9s9sUukV9PoHNNp0iIr+5j4VkUZ8Gc+NLJJwVudDDTEY8T7GBI9K+6J
4JAlyX+UL8JIpdn3XwqGlDVStNxgUjsiH0Tkw44OjF+yX8c97EBt9EX75JDPL1GKWLDo9tR5Qg2c
JD+8OjQGLNsA5VUUvdmOxFCPqD679iw+lFJNFSeWve52W+Y4LTVc9JodUf4pLr9LZhGSOu38i0HR
2zoI4RUxNe3KjHHxfGBsvd7l19cFY/82fcmFqVjphQIrP0dOthnFdo0c84WL2tuAcHVUL7Mn/MEb
xKzUbdkvV0oR6WJnUm1GwChsn5AzIa1l3Mxm6Kf2P1468URQlPG6rXuVD4vUPiW7oJRAAuNbE4l8
WmxG0VpsBOD3bQl/N4w7tm/DTO5+RZbzOQpBshhn2B5CUKKsxaiu8GaLr1KamGqHTA7ry6ewwkoz
s/FSsW9UzwoibDdoZAXJ8VDbfj1kO5LmyQ83BKuxZb8okydHYZd5daT9qVeBnoO4JbKaUGMsBxHv
XyAoXCPRZL3IbGDmeMjbi9SSO4PXCECLjJ1wIuBzXuzr3cYnNp4h6BFjA8zLjvjUL6lAE73YFgOt
XdGir/O/2kxUQlcRWHMIPDkWzYCRfWoe+UwQ6BzaUV2zUNLPpjTQRHPXAif+sxBp0Oix2nwtJrVg
ESdZzrs39i7JQbN0q8jF5x7f8xiSIgA9vaDdyqcMkIfmyXnVBZLqP8mYLwaxDSrSwg2H/4QLVXuT
buM2TFUmXjr3vMU164jDIkBJGZPRj3kHWUYbJLhLgiekLVmfMLvk6E2yDjjimz/1iCm5JP+7s6kb
wHTj0iOWjHLEZOxWeJxdKkTNRNmAEirFdMnGyw+Xf91Z3pN2zQ+BALxTVNSJTeRIjKnnaaBdcgQo
lJ8VbPccB6UsSqM84bowKBbwq9aB0XgMD1mZofKT6BCfjSxpx1GJ9ATvIlF4H07aVVMulqDOKgHl
F6LivDnTkdYkjZtgH4Lg+34K0mkH6X9mCd8FhrXRKk6PnCkO+wAJ5JX1LeVz2jyvNiM7HEz+UY9i
7TQZ9BNOx3f4qPbkjsFafznuEM1Aw3bwih0KX8aonWjZFUTyaYPQd5c+8npGqraVPZSbRuK2207d
ec7gc29XSpZor2rCqvLpYES3uGyAjDm33ZIeO5Pj4EXD0foPcTzthJqRXIaMGpt6FtxJUcV1ymkO
XNuj+gVSsUIAFUYwTlRSwRxISYVet3b0l+11zetJ4Ay1+ZLx6TK08jNxzIV/Zru3fNFmTtt+mt1M
OB0YMnLNscUnIQUL8S33ogL4ZeboV9SJNor7VeWKAbpUizzNqv2/x+gjjvtkohwvmae8aGdtaaXl
nBoIdlIVzorjdJS1d1JeTWXBw5qE9AL72IjfZH15M8D0j7BEkHaKDzN4BAiXRqNEh+l4KZZaKkSs
lRG/FlyoI/9ZIs+2zfHrvMcxnG0jtqLuBnaiiVqFLJlgqLSqMnzGvuV4BFJV80TRsmMshZmOLE/j
m52Ey+mSW7TCufiV+MCyMjqutJXSiDMO4otUP7Tf41KP+781byaAvXWdDLI1S5yZ8lycAYEudX+d
YNKgRqAYgeWf/Re4iaXgywdTeBhoDLmmN1ZWXkoxmEIy2w45Wwqn1pF0LzeWPQetf4k7pbw/6tDD
fGHCIyo3Z93HToIroku+2Lg/0zlk0fQDaJpHfLMvUMbCscR6bqDIoPG+YhLcseXEC1onQtHybYzy
XBYCStkGzP536p68F3cO6gM+8ziS/tXzAzVIIL2admPxTq/HQEc5tL9hZShZUneP2fRZPwZwh60B
x3YO0DVINfmXTDrXEyBDtkHySTB+mR7PDNB2cpW9t/TUlcYAQ+OEnFGz2MGSQiW+vJDQP3aFVwF7
uoxUuARaemcNsyOHWVaOrEla3DJQ+fsFyl9m90vuoLNs0w+QCjIPhdfLtScrBTxV1puBsFXvSNxu
ZpETkpYtb3ZacAWQKFfTbWNByM5sT5VN9ahCr74lXar/62Gaa9a9oakZ8qnGwIcuAzjb2EWAmfUa
K4ttHpgv5px+4XN2UiCE9vdZqyudFG5XKt0Xi7I1zXazWe6pXRrPLuaQAppSYYijUqxVQOVZr7z4
OgCx/BxGvNwhA+4xW43/nnyWEpvDu1U0gmKIRUOF1vP/HR8/x6KRfJjjb9KAl9ZjAi5rpP7tbR7+
D2+vzqEPJe4Q7zVx5BlwQk13qsPmQS80UByiR7kBZXRsrbacLX+Xdy2MKvrAh8272oP1PS/umYVC
wfrM3AQBahvGXWhWFum8DjiXoel7J6XOnsOG51ZmPCK6xX5hudRXfI8pUUT9anNL1DKB2FaSRHv7
PhWz6B1HnjK9DLURw8iG8QH5fkmtXxJWMEkrrPiiMKbBt6ti0mRKXOITleOB4l/IrfpxRXdSE7FS
BLbNWcJ+8aOxJjXANeBvUTuzUb74Y6h1B/UHiJR1Z8g/D2isM2K3o5o5Y883SimYFJvfnlM/NEDR
ESNfyIA72NPBZ83f5rXLcnOuliNVh7vJXvZ/xJ10hadF81/H6JOHckUzi9LqgP5BoxLdeZtciXTm
03JNyl6xjLP5V/iDRYXaVtDpEXPcigpQFT+3cBmBpbVBRyx2BB+Oc9gT/EHy3fVPUJIrG1F++Hve
RDe4yyjWtGopDQ9HOlicmgfFmbFdF+eWjqL5QYpASd54cBEWMz9OiB6GSzO+w3VvswJox8z+Id+P
5TkceWUBAvjPSrju1NpjJ8sI7aeUvyOEQgA8P8iIxBNZhWNuq9ZL6O6PRgPmjd6aRJklLkiTkFq2
ttDCdtlB8A2IqB5Vc6x9oecnW9DEFxKb/tMjqYknFLpFjTWzgpBZCC4CSZqa47a20QxvNi+qeflx
GiG8fTYnccDiihLRYBm03h6Nx6G9YUJRFbSwEFRAFCx1hM7vIT3tI/ma/Ce4CE99iVX+stL6w8ao
RhoyGfytAHMK2Y1wTgns3PnjU63lGD24C9SFA967TfKQUkGNwFFn54Zfp1WfG0EKga7O/jD8PMEC
2sSqf4/73Dw2DvzDe/dTZlo1jlG24Mh25rKniEVDPRyk1LtP8VjBA1neKnGnDk++ueVi5MF6rrTp
cbpy9n25xm8rAeEAgMFSAh07UXI38yELKEY9Oit/EH3aA2IhF6TOnmP5rxB8vFuIdc338ILIIHlK
sBTE7F2Dn18v3kJuSFdlr3fDqXwck4y8c+Sk9IDaergOsx8oqSyxQLSGZ2fD5jIqH6Q/lujAYVv7
52JuR0Qb5um4iLDFBtIUKWR3PeY1KpDyqzyIsbWQi+cSJn3pEL4RcdK0vwjzrbg53Gk+oECVCl8R
0w2eJTQD9xy3gLO1N2A5j9sZI9vD8kDH7x9VJfm3Gclvv5emm96GLl+P9pnhw4Gi/UKrOE+Lnofn
HXKm7cQy0xC8Zil0AbMY6Se/pe30hSCv7E0cjvO3XWZPjAYbbWKMKxceMn7cb5BkXahejh6kX+eP
rl76ub2WNnp0CQGd3vpGr/zTQQB8fhk2P4buINODBTxavs2DEk//S7aL8D4wFtA6jHwmpoZQMn2f
iiHwMKaMhVgDGYQ3FE12I87Ej1P2vRwnK3Ehmj7TwKr9Lqj69fpASy8PsojWQwuqW7Sd4H9DQFlC
iaUuD018l72RrrlGwmyzs6jiaX/1XLIciwSTOH1NC30q9So+L+9ay/1ImBvbNdBU5smcp4rm6XJI
I3fgKlseEIiSK8fFm/FX8Ilc2Q2NJMC/rkRGbFn0bGnU3DpA5L37oIH/i0aeCd7pxrk63x7RZYl/
NlNDUJPe8f4tJ2fzIW6PWpMDyVldfp5d0K6LtZfWS+GnF3UheWt2qcVTRQO8LM5Yxfzn+fKgkmhr
Qrn9LSxm92o/EpA871MnFWtnjheOhqWzCFzP1pZO+XZY4fWMhMKhsPeEB0bkKeaoMqJtOycom+fB
WAJ5BwJ2SCb9NCX6O3n/U7EFS16YB9Dgc5jhHWZqi8WGtBuWSP+ueTCEnvmQIFq9aDuRslcTGJFQ
n/+5DQG6+nKsq7hgJ7Dyk2jI5n5h7725txaEX+ehvYQaMI+CCXy+BIflyos2E2BDKXRKYlpyAspq
i6nB2zS508aWpyzB2WtmYyEXiI858DePDy1wt3MrMjzd0PvckRzbfmLLAkAszvNSE3IotWXwlRXQ
Qm9I+3xkNovxRk9/cICfSfpYFDRqXq2T1KUQveBXIQMu6cRYQQjgb5pEqswhBdfeYSay6fH9AXhf
dvtHoNJ18kYBL2MwJlExbGrjEcAimFigP47sYu2laHhYqX/7kE1Ks1TBWmkaJGOk0UQ5IHKvstK9
MpXAJIcGdd7BYurpTTYDIN7j41MTV48cwIifUkLhK1DsdDR+TTTkZ8yn6wThAxltxHihL8LqNd1E
NnBrj0Q4PLVUJqEoHS0DiL61X7OjcZR7IExdN/ujmVtQs9CMZ+ZVod8FyLMJPwNmQpScpvh39IEc
MHBkjy/M7XXglgYmwyk03Ux0j1zkj0hjOfwDG7Rt3Yk7gFdYa0Xi0GG0Tyg3OpH0onrjnFv9qH3M
mBLctUgbDhjbri+D11oeJWhCP63Trj18r5CRZ3XJujPdtzdOloZGhx2eun5sBScetZafDLs6jenT
gjnETg2V6EcANnzi3O/iY6Ooi/IwPDQSDZQFV8Pcmf5tflbQbrwXzbdzha4moQLbYElv2Zfll5UJ
VRJaGsNEBBRlKABbFbEwb78or0oXDuN6A+dYOWRIDjg4zs0Ak69qRc5xqBWaBYQ+Pj7dlXHlxEz2
Ny9KX7itJPyRZFHEP/148CxfARbhyG4XIaEilg4xvKa1bq49mZTuBMMVEt6bJPFVXeSRwImIq6qT
VcIjErfvy1pCJ6V5abyOTpXpgL8QTczjuiH3dbOEpVCHkEl5CAGxSRGHGPy8d0qC5cFIpwizJtVW
y10DKZbtVBYPdrY8vefgpykYX+OzPtO2jSFPDc68MlQoaEQleqQUPAZHx8qyd6qYNLyrrsIkykDX
O3cPr9JXIaVMDWkl0bpr/xDW8RqOWD6TcCs++zSkIWK6jeDPDePFycSoDhVtnZLfdIM7HzM9SrYF
iFKaNFxkS3MzfL8jRsl1rbA3FX7TFNZJYfmvolY86Xfrjg3rvbD8090gBsL3Y4P5LFsnv2azeEUh
goObOLS/m0BDLlQ/O0wCIBI7yS23SIIjo8cv6hO8JjP/JLGqE625deR01KPHug5ppJcD3Jc/3BPE
+s5smD0C+pQ4F0dpt3Ioya8TI3LgkSAXOjpNqp5NMlt9iMQn0z/GE4jQAdzQrsH6VSEKTbzUCMAV
RE8h6XQEE5kfC9yN6kT5uh8jqcuvRvrE/qsykLoZU2Bd9mG3yyxKDhRYe+EbpEeLgaftuc2iyutn
3Bbd1MiGz8XexziVX5UsWt+knyainptZNlZezfdayspv8GQk7EdLACWCBljn5GPDAHXIRVErSD9m
qfAgDEb9LGzrJzSzMlmWcJeFNAjyQ8tJnG4NU8oIe3zkvzg8EBiHt0LOm5SPHGtjUb+NJrwqGFXW
IcvoqFjt4cJ1qlC9pWTlKr7S/uK2N0qRMl3iueDKNuSsZbamP3QgCAdVk4x80BB/c+UD8756aB2C
o2baoxVTxWsOm/NOzq+4Avj0WC1vfrSuuaFhxjQ3xNfSbn5YhbrkCF9A11D+jLxnXa8njf04EcH2
/wYq2jw0pTExqI+o5F+DtQupeKet1eTWVB7d4VkTxiu5fpnzgPU3gxUaqnu2CkBqXwv3gylSsbc8
kAbK4RGIVP61C21EcmGXQMe43L6Zfs+UxrJ2sxZBWY8OIWy0QELiVsvWW2xXc9ZzB9GdZPtjS9oE
k37Q2RLX/0/YnC8i6EItM8lbZsk8AXdD8S2DMyr9HlQGDimpewT/ynQ0lHgHZwlyvnBon7pamaaw
LQBTGj9ZjEuOV8q9h5wgIfUH61Ff+IwxZY2e1yIBYTYQhczERo1QcTJl7LeFSyQpwlMV/xwq+jlx
uiwFCiXJRGYt7o5mb+WZ0xorn8eoiYRYQRrqIRtxJr1iYPg296ePZ8LGWOLZdJUdBtjVpBxJCK/o
x1NIxqucKh9FEccQkDXK2tPIvFLwMvrWQFZNYzS3QeWfqV7VZCijUpLqqyur+ZYljPfp6yHX074n
r7xYPc6pu3/zornaBQE+25ThBpEz8mkVLbqKfuixdHAlxWnAbhv+9hnHvrJ0wC2mRs/gPqzhXx3h
MEvrIydgXVa1wZ9o33UggsOPCQ3RH0YW8PPpZkH8/MTWo4EN0IhFhaN8bbuhY++c3Btmx4TZZWRj
/2I/+zpXQ50vJ7NJ9PLhN+tuXrL/caxFRh1D3x7p/g8+hdNgwsG9dqEnmIEIQgmeBSiyZu7SA8rO
RcgnuXSyJvJWoURjmWjRu77GiaeLOJfBvGGG3FRvAbsGBx78Y98hdn9C/vqSy9qpKYY0u2ewS9m9
k3RE2Zc8lAgjreYtPncQNOyFPbAsSiu5m4XqzmmS9BQd+sGoFmi0B6NX7bChoLjtzqz3oLgB3OVd
ixqaLQSWngU7pvq9iZiD0FOyzQtN2qPlB8KCix0q5TZw+MnzJo9eoUOGZVidHvDeLcZvV1SX/pB9
Mo1WkvlM0dau3jGDXwSFG0L3AX8Q2F42rVFwDsiUCUcghtlq44Bo5gJCh1C/F2ASHC+BwD8ymtL3
CgX6h3uszmMLWWgWUptmjafrnIzn5hceUwlneX73lEEr6JLzu0amzoVPqRJNvc135Nb5/9RnweY0
DEqRV6Yqr9ok72dcv+kYQfq0tF2f5VI9Nx7F1ol1KGtZKwYAer/YTC7LtZG6gdIKEHHKiPJgGF4M
PgyvZ6Wxds+uid13LJZ2fbVXSPDesVCkkcigyspRLAYDx/HnBZbr9S7LKZjaYSP3l7CtCCE1hKqZ
gTQWbV/T5Lcv0T19fKtigOMEnouwzeo2SP8wKLKWTqE5f55NaKqbTNMW83RUpQo7r59P5h6fWF3I
C48Yvug68xTTqI0B3sH84S5CUQkpN8NIoG82oGvjEHnB3ne3p0T1ecXHopQL27NyheUHMjcOP6yN
aGEJvQNRO+6/8reT8zyH9p/TYooAtMrJnh9xtF2yiktIGAr7ZBjj3UOTA3R61IzTKmXW+KweaV0Q
N4FvRTFJzQXSZ/CnO5+TonVBJ88FbXQhfk3AVs623s2z+NpuxlL6aToBiGD3mJ1qbcAqG14u3dzj
m0RuiLXcHlI5rKxFfhkI4cVyval1XK1+k8o8iwqda7vUR2AUA60zyQPAPp5Our22AQisMfIq7qvG
fcCLI9kPLMA4Qni9q4lJ0uzkCckHqbKuIejldEirpES9nRnIuu9qJcXq7ZSbuYFZ8z3vGPG9ps6N
sddd9vpgjnu9nV6DdSa0hB3al+yw8JxKHu9Ihe0++W5n8DwJS2Zu9kX4UURaZusSAeMZu+V3QRlY
D3mMeZAZTVudHH+1+UPyicibnpnSsv//dyxf3Lsu+ro+AIVz30s2+80/yU1ejkOCX0199Do8DAVq
r7Ypn1pDQ0Q6nLUmrSmAaXHdGU+ENbPU/KIThZBudK+aSQz68+DoJB++t8bVdve6psL2CBY5OUWA
06wWQgMByZbn0MKZ/QVjxa+RGfQESgjGGmZC9ygCpS2LKPEOO8AGHg3A81j0O4i0FlEH2LOmxSHJ
R24Wn+0AWxVVzEe2zyhpuScAB/2+f37ipVXLA9foS8gMS3B11z7K97nVmubVXPTSF0JkQJb8vGlQ
cBBuPpK7Ura9Q5WosJgMQ+AGBjAyFIZ04oUCOuImM7fBGfd8jSkp2XDdfRPA59mwc1YaosSw/dJw
0fM41qOZOQl6JGtAGo5Pe1Py9UOdIRvp9njVogNUyxt1xumHDKTjD9Xm2ZzGGpWkEE7gk8O0yOSf
u6r7/9cgpxwQXoYfusi8nNVwdrN7UicEu0oimMN6lUVIBu2VoHy/InZf5YXQNql4Uy69MFtQLCto
bP5z6PNKjaMz1n08r42K5B9+eANSoT8pLmnU7uxZvxrgfab6LSvRUQVSnSIQc/1CkW9U18aREiv6
TTOPm93SkhMfiZAIlbhRni8W5U4NZAKeP+NRW5hP8I90g0hBug3npBh+ivFzSJGXOmtm9GfELIWr
tWg6xbRJVgEYpzUriKwU6BfKQ32czKQVmWYzXRpNHlWV7yQnZ3b5Tcnhh1M/pJHK5khrzTQN8Eyc
L0aAZysSA/ILL5e+z7YrqxhCaHKUJvusAEgHNZaQTUF2iuRfwmZvb7IZ/4M8WEAXEhk/xLEVp9lQ
++O58/UVpEZVhBgMYjn0SUdYm4++1Jdrz2ZK9Vg/ZS3ckuAutynG/qqbV1Grnj0xb+vaF/OAkERp
LEjEekbVZ2e2oLu8kKSsS3V6Cptq8n3sGa4+4QUtyTk899PMqTHKaNXDymPaDGxug7OX7e1JhZPB
S7nXeOfNgOslEJVf1IOgD2PsJJ9GC/g41kZa8sLL/yztktWFbMJPwe7uxSy4pfFIzJ6GAtJqDP8W
Lhqk5pHsH8D8KWhiQ33zZUkfzpZZVe9ygtrBwHL0VqKwIUNtZiTRGxtY5KpuGmCMyiP+Kfv9Rl1M
tavyoBFSVbVd1Mi7W7Vum3kI+bjmcXNjqbubDfVJI84lDw6u5AX/qDUcfKhfitYUeTWX4PCM79dy
BlOU5EBdGsOQQFqQQ4f/abdyux8zspZl11xCNejX5t4QsSFl+4LdjwSUj89u6zQOfA6ZLuhN2rWu
0NcMuQ+BeIo7dffOwGUMiKEqXUr43yX7YrfzT+SGYrqb+8W6UGfB3qxB9wafswxdNTDCSNdfSZhE
xst21n36MxLGVhW1GnLXJECbuh07hNQA18ud2esEjnHBxAK83R8jcmFHmCrUeWTfugMDb9qN5yyZ
EPS8zZexVqtyayQWsyk6lCY1xjn6QGCqgK7Jx28n6hcn3QzDlJumTFkTkSdkqkRhbucfDj3dYo98
rvxb2XEjyBYjnYZMlL7izZaXZE7ONQAc+5Ymm/O6mvBShUapyaS4L4Ic5YZVTVwvDXW+QSPUaqDI
IHkpWbb7gndLmPsm7PNGVoznqOeYK7ALZ7NIbl0QobHV9p2XTQ35uhVDsC0PdHCfTVlNIaDGK69Z
hbOvSXpR7fO0RDIVMYCxOSD5Ie7TYL30Hg3dtvfDL+VOP0/q+5bG55nJo4O4T6x+91RjizOmqpds
s2+kc91jJWnvARsS4g1jjGis26CvMuu9RGFFSRU/yjxwntaP+pxoK5tuw0OOcGAfzup6gF+HwbpC
NrhMnYlDvKb7v7Zjua8moXeLD/KMYfWdFFnxndr2tH60SSC8WBhZaa2SYd63SZtVYnNoT0x3VeB1
6pFrg0+pIivQImMIhupwTM1Jj88+mr/IGoAdz0W+prvshDpAKJoY0kfjkAbTqVNpk/Oin9HhFP1d
aayaW01rzmH8jPGlGNhd2AHOX8Wcwq8DwU/aWhyfpkpURLBETzkHhbk+A/bRf7h9JQAERwLTq4KR
KOt+S53v8PmC8Vi4FR0vlWBRlgK9sENdWGrkwrGyuFUxi61GNJdEdqpre/0dJ+C3vYshqlghuwgX
EUjHpMWcSjdGuhs8LaWso2hjYT/HNfSPUERaZnrpV2kz2nk7HEQYvO9BFCt1SUfUK0JSaT6XzOdx
PbCcRWWHuB1kb348MJTnroGwWFFXUE22x+RrnH0WGD/VQqWzJK8/pXbC69NU932HGYr72ji/fMYk
WYFoxil16ROuSZfMRZzHXD/NIDkawcvpZeR/HXL4IQXSqOZn84jIW3ghl7Wv4rkGxID7gBK/ctz8
RHf0XB7K/RydODrm7OetGzFVXs9K/cjUn39OI74DBiHBuccMO5MDvJJLDixDjxaFbxUty5ZVCVLl
ll6ewjUHe+Ryv4RoiG/fK0hgeF6M3ejkTJNleKIrZQ4WC0cXHptF6FXtBrG+frySSShdAhG5F4c/
R3s5Mqy6t1X3kZl+KIm/EP069D/jO6Dm1/0J15qGgWPr0ZweDyPKsfi5mDzwnJjwR5at/ns6+Xj6
gH8UxXw42oT7YlNf+yyaw+lESqVZ8ag8t/pO6ezhz0zFAileIe/j13D1SrdA3CKYAoFS4IJnXpD6
dy+LCxXEcbrWLqNULiCyad18A/Bk6cl0ZBqsqc+FbojS9bYF41u2nR1L7a1JQc/IO4OHpM1KjKis
zpO0iYvj0szU6h2y/ZWH8Y6zG23Sf1bCBdloBkr0CJhY+Kh/fxIoQr24cr+AAkXEgBZDTGtEETRX
eHZv5VXuuRFo+gog7pFoC8jgRXM/3D60k7VbVxI3rcO+EIsvgzZnjj0itL8zwrhdvsn1rVEbXhGL
DEzbWh83uBHwzY0vn/A82CrUPTAkocBmWN3IDGkhwfo6Dkykh2q+ZC9o1fmmV6PONf0Q8FrFR4QH
1NLNQSOo9rq4nP1zIlykeWg6Swn/gsD//GpxkBSO7HoF7C6G0jMXsNBn8+Ok0Xy+zKOsBaJRl1uk
nIFTUAI9ymIoAUC2GIX8e+6X7mVJh54RfCIjbGNjfPPj5Ntz9PZT4uSRbi1/zqBIQVysSVyPa87f
gFcd54s9eo/3NYHfWqU+TyHdHtQmkLZxvioSBDgjT0QVb4Lkh7E+UWEmUKECnemj+nHesdnb6WdW
A9kCZdqPZkQhaBPaR1u0XCB9YDpi6oj2UwUZ1jgiMfD2R95YMU8nyByxCydgA597BFPlAo1+OnZX
aX2DgGihsLAswY6J3ezM5z/HEcHv9OS0oyXeW0NJ7zOwQk6rR/Kr7oIAXB4Mscd51rnaTXaTMEw8
WC1hfR/MmmhTmsjAfNFbIX7vbPkwx2NaavqWHzny6nIWR8Ouz2S7YNKpxpSJPVXPcK6xwU+/lyit
bdSeJIobOHaaSJbbT9fVkOCcAfbXVUIpKPepk6P4EOGlkCfDoiXoGqUz21bAlKVpb0YAEZ8JEPBR
14uJp21Y56HKQa0iFNG9J7VlkyevDOhKW73CtEZTTxcV0qLnWKLh7/BLEgvwFJw8VhZXiEJMkBrA
FJAAWaR7pqyu4R2Rs7UYbZAGepu9tEXnw82nqaOfT5gqZefCOpGEtfcjjcffEBq/CjLLuZnEzVzf
jTt209OFqEpWfaDHqpsrN53WQxIWv0CDz27Cr1Yyhb1edRRL0DRgCyChMDJSw030bAALoF0Chh9j
luHUn0OUvokgjSvxiiuIrxe9BMjHHoK3W7o14+34Bues9BZGciBLekQ9FemsV1tS5AdGAWdenf1R
AdsdAJ6SGQC1tBCHap5gkP6nOmzsRqtCiIfWmoNlDMB/KQZc5j9QN/FaFP5naC8kB9S6H+9QmbuQ
gWirD2AX8fut+TqLc/j0YnAS1EMrc1VfA+qUG3tVGTX7bfex5oxrZsjdDkZvqQ8qsxti8K6Wh+Di
V5Jf+WF9+2k4+RK5lhe4pa2o077O38T9jzP1wKVTNma65/YFG/ehDAHYe2sPhv0CSkIcz7X+DUqf
tEYi9udM4zyk7eVokfT5U+gXy8QD5SVGYrNIag5UuSuwtmYsO1XHvKkuqkX+h95WIA7Mg/wOw8XK
MwEb5xxYZooiYvpwQpLyHSFDSp/MaOkhRSqAuY7BlcqMLdC3KiA/+XBaj6SubRwJjGLaHLnHtpW3
jtMh53jlSCtDEBduJgulhGU/MwKKyovOYZF4q0Pk5GKCA4iLQZWihdaJlVJM6oarYsOXQAz0wCtU
7S1uqsXxVmUmYg64UXXVKuOB8z9xrX33X5DuYWxTLnr/D6g35JWa/CPIIsKM8Zl+zA9Fs+K56vMK
eqALu65LYOE4T6vKhIMCbWCrBI9ZXI1BC2+uOJYaRLZrNmnFMDdWIfu1vtGD63YcSFBUpn6JgP/P
futBhozjsfinkRR7SRdovaSw3ryOra9Gcv8LVqJU+TRTdXNNnwqd1NHboMeAiP7KUSFJSjwHZLW8
49rax+v1YRPDVWbBSOu+uI5ykZfe0WTQkHyaUXL9EBFZ16sUuT/DesKZPX4B9HTk/7+njDC2SgEs
opgDw3uvAk32SqC5jmLHtTlTRTs7O/5nK90rA5SZjaqfxNKJ5617txA0qLaM731CcRlpOb66Zs6C
3oobdB8TmWRRWg0kza1JkFIv5R1ftOJTlXZpd27GlVvBoiUTQ113G6WDN3UfjpSWXYYKcygT3IVA
OLJxTSgDOOZ+fgK/HD8ZXEjGkn37F5I1CD2g/kdealGfk51WjRxJdB6SwxGg3wx1fVwTRKjxzEvP
j2xLDh00khexSoN04iQvFxx7Lsat4BbvrARybTYP8egqdqalYfbqGOQ1hrGzVNjjTgC1oY+OEY5M
NjDgU59b6CTxH2XIWY1kUqfOPeyOuaK+XGKMNYt0/mfQZ5HLEwH7k30JoONJjWC3lrMgRnURdAad
Ngp0rfUvP1cU1oJ7k1z8VijF64p9QhgfLYsrMkeUqL71Zh6/mvp83DGv2Bft0xOE0/F2Nhq9FMfc
h7JV9ycYyhHXUtNtyd5K0jrlunWTkX0MtYdqV4O6ztFbWXkqsLqAQCCyDGSjkn14hj8S1FaRHSuS
PI5uGdVclBHlMdPYwOtcAL59m+dNEp+3wngTtYpBLggUJ4SeCq93aPIdZJwKs/lcZskFy/wmUFKI
oROMlEmxA+LL7ml7+A5Y5MLliTXQLB0L+6uwCErwGp8OWK5f7Yuei4qX8gIB3c1I57rKqgSoTD1q
P2ee12sn833hxY9qxSIowoAX4aqv1wteup/KmVHgylv3f5fT7Lvjnsf1Zh/0ubgEZ95H6yvNcB9P
U23JkTHhwLh0xOcPBJ6g1A6VO0NIrfv7ShmuwZ7FxDoouJpuUcIoYpraa8UgEwIXsPii3Npkq7dj
QIHlh7Uou2P9MIOJ7JM/TqrNwk4IK3LK06z9l5IZ7Or2edI7U9JLsHZ8Z0iFbEB2rlkp1VinWGlU
8+2Y2q+KEySdL+YyWN5PyLZdC96XYJ64EW3MIwsMglZzRSIRcaULYkTL7pRbN91Ceu/4VpX07gTY
GuQx6W+PKaVBMTllsTl6WPafz6jxYHnL3pf6TTQgbutsDSl36yPoBBp5eBxQxDyda6PP3BVNHBd0
GHkEJO6nnY/UD+zLzdhPCCo42foGjskfri7akCloDeHfks5/8gHGLSVH3/JZr91DLGIl9zV8tbCk
qhpqWCQG8/4c48Un5YVAHB57iLj5M4UXxu8eaGWIOLvdfOWw7z0EOFcNU9OCKX28DztlB7aPgyYV
osyv4jqDD3/UworY6Fxy/TYltDG0TtlGNPw+OMNwq8pXH+MEOzwixqXxKbWTtIJP6xb5WbXpZOft
WcAvUxK9FDPD1rSAwp/q7tTrRZssiSaCZrahFOJP3Zch9QvXlQDdO1HzSEqjTr72dasvjd73DZ4m
gDVSjnVD0tYoSPUEbWcpDouIDYdS9iioOhIEOcxbqDHhmNqz4N5sevBjXNS/0cw8iWxoc5BRPTL1
DaTI/JEAMgofW4nuTKK/iKN4gsbwsZMXWJbALE7Ky9fZdo4zE0jXujMg5CMpZ8IuqfMe+M2zqI0s
onKXElDkauquWWbpQAQ5iTz2oggdcsAglncIsnlhpvJkkUvYztXqC5j13qtDBTNlYtCpEA8XZCUP
4ZS5Ahk/gh3KQE9w+CimRz7CGWcqhn1f5dfVe7XEieAc6S7KTGJMuKCtOUgRX9R5uzDZs8rB9hIp
/hTsDLb8za1Bt4mmYrKYsS0zm9GSUWj3lTbb8Zrdy/KDNi21TIoK4BNFIxchWEIoutCvHVa7mrPg
f/AsKxxbb6MdKwmPwlsTP3u2NuJYSPUlYySJKZL7AF/f1mkHKQy4w2/tdy8rarweSv/7H4ILx5QC
FhORdb+C2kP9EnquRbLgkFQFHJ23Kul+UjhINEhrp8/qhxHGVidBph+5Z++Th0trHEnW+vcO/MxV
f+pPCH0zQl2KlU36TY/MwO4zdI8voeppJDgpXtNw6ZHQdkV9bhIiZAIz6EBuKP3ZRk1CjOPeeawj
T9tc50NRUbLDRZrou3skGYU+zxvF6BlCiWG2D1AFpriNtjHh1mE+4SWHrJqdXi9Gl6ISuIANZp8N
X7YxEjYGqod2W5OAafVxNfKsb3+gKywgUyMUourn5PH9ND1D9qoZwKiysvvh+2yjMtCpVfAPmFpQ
8Th+KQ7GXq6nV5bB1GDtUrjRAAdQp54eQCrNg3SbUX+lS+Nvw5fbEFdAbyGiawcQhTMp5y24TlBh
UW999YsN1jF3d64jrL6p2oJlR811gkUe0/13pj43DKMqqHI/EvgxfVHELOX3g7wFk1vdCLEVivyW
jKm1i26IAYT4jHhh7/R3Gne3VIL1JMQaNo5/8BE7tGh3BG6uJ7qVXQeMXkXh3m0LPjecihUJsAYx
Bz0OZiCuGw0375pXA+aR7zvln/MV96dYS+89sabpnFstZH9b9WI1zJ9IMZ3+r+k7zlfNo0b33eBG
GKeZnFzwRwbdnHkER7j8T5qUa/IiBaQkoDnxQkdSY0jiMUTnZAUGsmLpTO0Tbu3Zmv/nvIW5IKCg
I4EQlXXaIEFbeT7tT2OKH/FmYVxWcXAgAT6DyLQyZXk6sDzd2YPAKn7M8C20IhRsoOGW1HGWaOXZ
B2DmgCRmHqeT9nTqoPk9PkjKJjsi6uaWnkxcrw38uMFsX3SJMbVcdXBhgB74wQnUV/wn32sg+Rzh
HofXYthvIo40wwwmUkch+7yushm1YCh2evaluczQ8ZOh/tcAJGLvCaTjqmhVCMm8BVZm7ubQTnwU
X5oX/ex+B6+5wYJhMBSWW7xHQve48VIvadalVNT/ATBvifEygwYzqHCYolAcobhRJuZr352VRRu2
iqFvOB9pgpXyvhnc4sGw51OiFo7+VCZEuRAP0rx8XwjuEYxk6pw1RWGqQahW8DYPpnDHiL7oXTVc
oz6RhUiia9DXRQ9d9brnb4gwXvaYnguVEWSK5IujfO7JYDVG2cBKl656A7+XKGD4HSUz+TBSVVEQ
IGFXKWzzD4aFVpIRR56YREJb1OstjIGIztMkta0A0PT+TdOhfjvdmUDowaMNxzdq1rlNefoTW74g
dxMYMRUJTsOSlikvYUmtdBLfV2DZqsFicY72ljoceklCVE07t6V5Df7RJ8m3xRj+dCmBFbwHMS9V
IijUsNm/W/5tt77SvcMO7EiuH4ca/Q5aw6mgQy7GHZ9azO+VnYbhlTxDAXWg2+8bPVMuGu1YMj7b
PzYXVMWaWLo+lhUqvoZcCdjpp949Cnh+xVQC/BexA+CoAAF9sjvsMoG9E3mH6Gf0icziJDyWLxHr
plyivnXmXnR18HTVZJt8USi5zE1nq/HMFNW/Vw+03nFYSzC8qGWgq00XLXTc+PHazDwYzFhW75BU
8TDZSfrGAnOsoJMeG6bf96sW9qe4mNpu1yXtvZ3+vEWKhqgGDufHVcIEC59mTC4XFJ5yoPrn1sup
RqmcDgB4Jcsd78/v+1nvX1P0YK2pjHwiBJolusW/eX39vgcT71pbkdhZcEIZBdtXQz+Y1Oy9LkrT
t9KG2Y0sCgxnjQTwDaTRTqB/h0P3msZ4OPaHofY5VLUlR7pvZ80TtPPgQ90NfP3amY9xQ6ORO354
JXKso2MEoGmvs1o2AgWA2432J/+zcrQxvM/D7o0DvVJuaXU1a5D0Fvb79c8rb3pMYdeE1CzylhPJ
SMfFpLeEGBbDOGmjrWY9iTNEDFjnVUCZZ8NFc+hXkBVRVcQ8nFRxUl4OizKuI3mW28ADN05i2+R7
Nou+BIgMm+t8xeiPayila73yw+Ij4uRDHWL6GQr1wlt3lsE3jyqJrV2bHhG+m7G6nc2BdnfUeX2i
AHjDSws6sxcoZOmUthVlpz05Wsr/cC/0NqnZuQDgxJERgE/20qgU+tyjNqdH4/2bJzz6Xd1OgwOU
80AGrrKrzPvTR02kVbWS8+YM40Ehx6WdlBUG/MgWicbaC5at6/2iZhSKC9g9nlfQpCqQ9ETVx5Dw
eVVx9qnEqvrdsUPXuFm2OJCmrbRcVf8AAFLTQ9XtLTGeu67jzQVZYt2A5E3h5fghvVkuf1Q8I1KH
x7DnxHRtsIKrnj9ETLpB+uraNCxjPJSQw9NllsxuBwBpNRvmOeanlM20s1Mu02q3HQeR5FWwJ293
CDRXFuBxke+B9HQdHXGaRLm/OunuXaNtTj2pJQcxa/E5AtfN6tLVIYRzHT4sZ/3yRfzgEJjhIIMd
aCK8NVhvs/rmEpUC2QyMgtniHhlTA/2SwFRfruUyfLGDWTNDczWjrRFwu+hFz5Q/wG0+rlv9e3v7
6S0C8MnZCbXa/akeX4MUUbf7FDzdEK34oMMEPP4X8skqJDS/DmUmFT46ncq6YBVyoGt1DNSFQnNU
t1T+19piFdrN7dyrEwKDE8Io6A1VW8pAD6vmOzrTsX7f8AJKj80tF7G/ZBF021CG9pqc7DJh0yZt
NiFUhmykulLy9xkFjmJXMAKy739Y6tV0kdMeHVVnIZy490Dy6G+Q80dERxsxbTqf6tGZhClaDGwe
yhvygc7Uz26B+VWlv0/HOEsAsuWT/hJttKSQrszA1fc/7Y565p6kR4Vc+lpkuKW5gRJLmO2QjO45
fA7yooIcnzVHSeCpnFcWrkgxjbWJpIS/eXOfsI6Wr6aNC3d9OX05X4+OCH26M3rfwTuPfkFZr9Nq
ZrBCGyDeMAEke7doajKmtLv4cZzUlSksHgkSM58d5Jp8VPbqMZgVGeV7sZdJW1ewgigMNlN9H6X8
hbKN1S2q6y2wsDPqRSaWKQFmv2Vb2BG5vCuMAcB34sJWWcF/yoH7/Zr77k16RNKrPdRKNvvPseqG
F4ADN4N2v2v7quhWIRT9tz0WpouU1EOLIdDdDsKrL7XAgVS82Jz+TPFar1sO6SHfme8UAYwl9dJ5
VD9tHa0/n78OiXj4CYghvzfXpE5C8T5NARMEE2OnoXMqswI+Mqrzw6151nO2n7SfYdQDRi6ACpeR
D387DlOjNEoP24hbrLi77CkGrdBmBPYdVVUroUeZPNF3bCnkByWvyUrw+jzHEISF/sSUFHAOEP7a
j2FoeIdM8nJD9G+k/34v+NjzQKUFAsvFsrobu4RRlPk4/j/mW9p8mnvqhE90SmV/VK7mgzG7AkBj
3MnaeJHjs/175r5rWJJ56bJVWtBiAXmfzlPG1sx8ia/uEcwZRXivUPlCiesPhl8fu4DjeoZr0zwy
PrVnCHnBF6GzT+9Kis8F/wI94/ctw9esL8ho42BILo565A+9/ry054Y0l8iYWh+XHQEdUNijfFQJ
n7e+rmeDfMX4MpNe/wbOukyVJmyKA6G8trExxDchgSWpvyus2UuUOiiLAc6gtOC2xndDN+rbKpGR
AyyhW6nn9I4PHWQMlX4ezndbD3hyTKlw6T0urezsjhfMEPkZI926/xKCLqdXyHmSAuMcS6BGoaKW
z5A/z3+apWbXA7HuLtD4WAeKp4dalqb25mPlFtOB8kArERG8hngb+st0Eb64t3BhatJnhK9c7y7E
/bhpbZRDKKvRXCIngxyYdHk7NWhgSdUcQ8Rff00N8WVekmXrcf28iNmKUJQ7BVqj/f9Qm/3rxJQB
FU3NTUv1Hq0jtGXSfH/9Iu4XHZQttOxKRXoCyAi6F7vY6PvPgTiOdfxXkW9q9Rq3ISFGSZiP66DO
RTvteqA5QKVW48EODBxX+/+kaLWOxUmyYzIQG0f9KQHPxPv6nESYFRqOleCtbN40TkrtY1tLKN11
Lj/5AYaeOdo1ritPBUrm2U1A4sDinYO5LvXTTKMHRF/DBwytOVRYDgC6h92aZs4XwHulOpG0qEwr
dUFbIttsVjpjTwPngBbOxSkaE/GoBbbVzyMmBKAWPxKQ+CTupfSyg7LX1WVCA6FVryNkuvEaznEB
l+7ELPtTCLH+IniaNlioOCs+ZulX2EnpqSe0lluKrX11za+2/mLg56qSk09rfvRsJpVLZHkKZaln
VkOa1NGXvsWawTvEckFJBPyJcQb31MU7aOiLjI8D+fjItAatMK1XhoCCA7Y7fpSTWf1tV2wmp9i0
mTV1cscDQNtrAPYNrhhEH3ReCHI9LfyYvsuQ+bFJfX481MDWQz51gnTxrKPaPvxQ6SwuzwYq6yKo
gJQ2Rcze1h2I1hO4GeZzpgSsHBgOhxnFTgS3qCiZHoda6nEhd3XLH3U0tCntpBFhJpAs1P0dJMKg
VUNuOGjpV+UVakVMF3HxsAZT8KP5rpzPH1911G1F8NzE+k/WAQ2pqI/ecVmpPb2wmG9lesVIJrn7
XmAmhpN8bbxDzUaQOUgQEUOygd5i59Q5VhKDgPmTSBqBqVPiPrMNFfxjffmxrxw4x704/ZCFZmI/
PrOpGwA2IngZvnB7l+K/paBeKKBYk1Q8yyaPwbGQLJYOZe7rPfAwfaGcydvh83tIX7vaZGNPK4oX
nMQmOQfdJomltywzVIVwuJjB2IMkNICxYTqS7+68H3Z0dIDrmCML+eG0noGmRxfZJ2mXKdBrjslh
EQ+K7p8NbL3SAYf7nORiMhebd4gH7hHbv1t6Rudy6GpY6noaFhdB3WwUrojnRZsNv2g4BP36NzBq
vimFcEZPQqHJJX/QjfaxADBwfugz0t3sdRQClMSZ+wvynf4NOQarjEqrWvtpG2yHapgWTDcyFloG
PWcxohXPP4JG2AZY1RjSUnymiF6sI5iJAnQe7nwoxJtoRk40S67q7u1MsSrlJu3G4GpUQz/zDqML
wVzMGWT4cIDXJedkkhNQ6eIo8nbDTnAV+2QR09Ikb+xMbv7CFRWs6H7wOgnilC/aJGT6xpw/y0l0
yUnNwYjL+5sdZFI4Hfq6sX/7F1RGgBCxzh8Bp5ho1Sp9J5XOQ1yPhyyJt6IeeN/oP264TSbfuzaV
/2w33vaLIoLGFF6oT+EhGv+/t1yLQHozOTukrKsU6C0MjcWMMCg8aRX+JiKy2Cq/qko94oB+VJ0q
2GQeXj5SxPVP2d9EulN0jGqGOlx8lfQ4MTsSBIc55O8jimUH6WwIIass1BbLP3CLmCGYM+Q0QiTy
noHCOvp65TBoYrsk9xwge7O5LUlmrSXOFtg4g4nKE5Z1c66Bf5YI8i9msDuHMYjjlTSmLlzAW5Qr
kEYB/quEdmrT7xSMEFrRW8CcU+KbE2ieG1MhQxokVlMaau8PxTPK7fR3G0M57UueNCd9DBReGFut
OrjUDDjRec50prE0KBb0yl7Vjh8JyndLbq1RvcQjGPpheOzjud6byY7gfcuHDY8RZvE5ppLgZyUQ
zIuU2EpDir1B/2PNVWFgm/tFh2qB4qFHp0GYcVYG0zjsloMqzL5eqqo2FZ9SxJ/bARB7EYoD7HxC
6KqNG+/kHolJYeoSkEmZkBLWLo9yWIuf7Dfp+4dR2o2Yazd/cOkkor6uqoXBUFBj8PqWkxb7F5I2
0pjJL/B6PaY213a3j9uazJawp3uI4UNHsqHRmSWiNRnIHWVh2a742TLjZ+AaOxOE8XCbbKBVaiwg
TsZWtKeS07dAw2S8Tfo/LFJHoqGWyiqcuuOjSh4KoPCbZO882+xPsO3P8GcRCS8mpcD6+rAoScVs
kM/KloFv7QqZXx/TFFWgx5mPsd54DEuFYm/1M5i1bYxeEXs1VmSY8QQobPdfV9lq9x4pyBwtDNqV
2ApcRSA18Tm5OUf+cpNFKOxbzPlKoNl8WiiDPa/aCHQy8T0+8zRr+gpCle7cHoAKzzkXZDzfuPio
PigXv3ww9+1M6scbc0Z5WKf3KA33+BS33N9MGPtSPrwGtKIJy8AfiM0SAw9zN7tk4wOgfcBc7tCM
BqUqL56ChJW8M2hJiBKVp95kLqPcZqd6vCOTDOfYqS0z0UPjsjLyj7Klp8a87XU9B9t2hmn2oMDu
hysL4YQHQ7DBCZtwIRqbhI3+rW/7wM/oLetMOiYO7i6U8KUS0Cg8Y6UFdVTEi3SOyQVi7tOeoadt
e9Wy6MDyLJe252QxBkP1jyJYyTVq7pmWkmDTORXTzKeGCp0S3BwB09H2R7Zw+md3jQsrQt6PSmcT
ymKp03/yyXlUj8LTr4/xcTY+G4ZUJ+elqxNwnMi2CmlWRwKQ3PPVCuJjkDxpdQ/LwywYVdhh5452
IKnE3MDa/7fl17XdR0Z1RkX6/UCSB29lzrf/gJbIEPhMFOBMdU2OzUiJOWaxByUqZrqMNXD8UmWH
sT3cqWjB/SF+1vZvEvAqNOMtaonicG12T7rYIcfXdpFKQXPjjkouD8NgG7voIGESBAk6gfZ6tPfd
oWj4nVpnNiKjyvZqYnofIE/+fDPcPJ1plZoZFqPXDQnalv7CgXavunXnl/4NgMxH8XqqagrByfbp
ERTurZ1rvUuW0u1lBAJhpo0Z0XQNO1pCpRYtE7G/s+FBxs8AaZNIHa2R69mu9MwTL0kncI/63dOv
BNey/qbaOvEcPEYTp5Af1zqSYQuHKjpsG2B5oEtHt6pjBMtoWhJl/vJOWFX3Tj9T0pX4+pvdtytX
AhfdQaQnAQZLWLLL8gzzbiu04m54V8474JULhRlyvVE5f0DsB7n4+g2d2SOYnBGzGX2KkjoMcsKJ
iK8ymPgzFbO+9BdNgNiWignXOpdjxNRQbOqM/B94pKxC2dLKYyA4lo088AG+P7HL2EJDHqzlMtDj
DFviubQnC+sxgLvA5Q0qh/TGeM113rVQl7PuKFy21g7F+hyCIUWGTa/l8pFpgDte0YJFBJ21/Hd0
65m0SrG8HW2ys6L+TYcHXDXagRBx6thC98B6h7H+PCaPwuEKRn33d/iNJhyzM+njG+6z20pl7jaH
wK8Bbu1/4S7MSN7CI2OiaaXrKmAL3qZBH0wj/9c9WdNaief1AqElyeqCtYFQmjf6eRkeEO0zhe1y
HK8O0fZs+GXhL3JroN8o29CyRroMxX2Zk6Rw4zljlnNcyzuuHOPxdOS1fhBlXYbjlxlLfKMluTm1
1MQXbtxeXGAKEhbmj/F+kApS9BQEKMza/FcY4Vi2awoR5U/M9VLG//RtjRiTADr0GoGei36U6od+
I/9LwxfBT/d/TClK3CJbr4GJZfJA8zoBFzM+K0MQzbk0Ux0hqwTNGJKz3eLcXFnccr68HrnJE45J
Xf3r1Gd94tVefsj7/L0QoEB6/IPlHHWHq6XGu2DZNzaBEtd6xfeAIq4w1fKzdJ6856+QG0fXdudS
Vl8raJJFOD7JJ6d5/UdtPfEDl88vBdTP6zLR/HL+IaagqoyPYZhvLuTVrV8CxS7patKv9fz1M0kK
xBY/UxEDrNgem8it6PndNxDEnap4Q80vabrHQUFWpy/rkxoLC/Zaj9B81LD3kdlExYNub6ER3KJV
UrC+XZ9xv+fVg0SlZfVZc62O1joQXvt5CRVneHhQNkb4V2jB068kGeNENr5zYLHDvYF4lCspRtNA
WW1jpZnd8ThaWR2oLU8Ryzmn38BxIfYmhjTK1evN/+q1/4U2roK4lcQqJmaiqpTSbnBhSLId8ubu
rwVwxDjsUXegpjlv0SIx8GhluU5SjtPkpxOo/NTqSyloSdd64flf8UQ4rzVCKn6mxNp6Ye85n8bs
Mcw5gwFkIu0VnvDeMUrW437egmar3dvU636KRskXrwHnUD1sYlTF7+i5LWOC/AkYTpclF30qLEnZ
ZATndNjnfS657RL2yfQzetboah8cObUEX0zo/XpnAdG1ULPjnXo7+D564A9pkpwxcH21blQjuXTv
5DkXrJj/jxumL0OaxKOXOes6pC4x+LtV+WbSJQt6iagw798oygPpzUeF/cFSkQH6sFVsxrMg+2p2
tV9Ro0ASYC9FWtsrgAjqX0L3WWUoNCMyIblB41tZb09YpvXBPhSBZcNGrnLHmdi+YwcJK7XbQmrB
tVe/ksNYFxc43cjyNpaTtjIHyTFBt+ZKkSFA/LXUqJltbqPGPS0Lluhj7Wn4YY+iHKlPCwyfOOYF
0KERdso2lh3EtJ5EpJO7sWB/y7c6oyZvOsxH97r0xorafDmaVOpWf/+xQhbytjfURskflelleTLZ
LrQgYOacJFnF0QN7XfZfostdMmE6ZACi1CCBQVxTC71jko44aTwv1qEsp2Ep3AmpGKwiFIRJ6Zc2
/pRNCeO1pOsMEpxM7h4OpjxWi4wgUMuNHlIt7tw4AFU5BqfcTWVBPpd9wrd5nqym5+L4a/lsTPbw
XwrYWd/BFnTjXNOCLtOktccg5Az2D2+0Sy+WnlVNkXY09JP8qklHtZSoZBv+lWfn+SJTmVXyUnBP
a2F2UFWQU105HTgJiZ4vp246SksPqiQHNEGKYwY0Pt3z2N9yQ+FI2iE1ZBZ8q1zGEKzZnMrBfDl3
Floj2j/zGNZxzQHMqYG8QXYu0OhcUDSiKkdMT7jnJXVxivrkFaw/wPJmeCADxP63sVvC7nc9c5Bc
eoJJqkdjNcx6MHq6gN1ssJchg5cT0tngykm/fufPHCGlwnPVIDJmNTKR99owJwLGEoBt0UnP2MWP
A0szavZ6YX9iunNdxZP/WWMx8r4H65/7OES5aW0HQJjw2nFvB/FN5MvkUdsb7zF8Y5UY30TnB7VC
L+HO4dCxIBS0qaaCbQyBrgGaEoXqcCJmYburPc7YcxjhnpxSzn5cUlCGZe21i8oCPWmupEbmzZqO
MLkOxCzuZzLFhuGr187W8Z9fTvfOip/ZhvKxP7PQYpBzCBecB848BDY01JQsPhts8E3l/GOERNyu
t1MsVKnoBXcRnoCY9nzarAQSjpMHZdfNitNFtnY4KMhpJ4DOSIvLyBI13piY3PHdK7nlpaChT+EA
6CrOB9pSlRt96tdlsHbZeT7rd1wuSuXsa5txgKKjehQH4H05dME8Q6e+BnKMJL5+aa1cLhrh7IQC
ufdGydZmnAtw8NxAZzMxFJBDG8jXgOczF21W20+lCgMQUWSBwZDpiBd2KJBy71YtZS0gpJC52LSI
ZaOtROWbjy2+BZG0mRFw+lJpkCQVvi2iQdTtKTeuxu3m4bxp8QgZvHOd+o/IFFNSggfWXK4m/DEb
va2FRKl/f74+kM1bYxZvaVX5jIzpWwN8SB0skP6Ws24hfs4IP7MPFbno55Whn+r8JxrqaqMpN95F
zY1/Dch5jC2YcDO9gXPTjS7i4ilSmN2zBZ7JLQ7Nzky5nXSG95LH6H0xnPItAicEkAqOh6VR+iZ1
r9TNTTzLngZ/Oq/zrn1KrqUbg1kxUZK4FXWBbvyFlWnYNYH2fXhlN08yMQCtQnEXzhsolMZf9QCd
1BElJ8l51AcuvUGnRkORXfZQtjhNSB11H90L52ZW0OEHHCrYKrsr+dAwikAxA1fXDP2MdY1UVJsV
/Ef5ofEhn7Tl6N9FTOJzF8SraTqlepTUEKkI5iU52NaseEWj5DyWYnbemOlQw45WghYPTa6jdkQv
li7W1COQNPKVM2C421ZgYvMVz1ul8YcbwOdKbpwEaj2+omfCsHTwFP+R2Kf8mwwh/39KzN+81Q+i
YMaJXwJ+Yod4t5eNo/jekyV72QP5VBWYgLwr2g1VBO3jyz+GUfdUZJFFIvmQkO5q38M0EHFAFfBF
4X39JRfwKINfdx/VvBim8NH+bPtJlxYBF5zm1JfNUPwIPEII4bwPVoJKYIeHly9cIqzmL8aJx2w5
gxeHz569ccDL8rw0lIzyaGYrNakgTTld9P0wlPVwnUN5p5+W2S8x7nf7aM6H3qdiNETN3tuMebJ+
uLGO8EOdmqj0I4ZJZYIpENmM5IgTcOUMmxbhFd8wg+gOS8sLanCw+oUiKoaDdJ1gPN6EyCvM1Fyn
aSR95QIrfylA2f/GuEcfGTQka4HvyDvxf/pPGfhk8vVW/JlN6faW8LbLcyAX2sjsVg+tmzBt1ZXm
6Huk/T1Qza6XWJs976Snkb7qrx5N6NvELOd2GLH60Nb7l3qftLoS9T8I+Ayh1T/KJr0hCmeD/OaQ
n4kBuN+cUNHF//Gq5nw2TC4d4jXUT9lghmvvyhFxyWcBIM53BT5LCce57FfFRMF3yOCRuDkNDgPP
gFYUA6S5gO5019hZjTTP0H4nh0pjNY6nVnvk1qArSDSYCXQgv5/X5yFlAzUf+s2nQVb1uRoN2Z1B
QLahLCvsrnh+Vv37TsWh532t479gNvgwEgvmeeSbFssif2ZD1KuFkw8byrjdSo2QA0oK4LUQaRi/
UmDZC+T18UO6qeyR4bFuD+DqwlUKFfq8b8/nTZeMgd25BJhRRxh4Zs9vXFPhpRtfV7nNuO34SQlE
VpYDxnxzP/3QxwfzAGxBqM8gAKe57ex2dgllZ+VVf/GCUTCJGsOKOL/LHYZVAHNq/bn12CEDvNms
3j5hTMk9jN/RoUfSNk6rJaej/bhOBG6XVYsKf73Z3u0gEHSNj/EFBg1lZX4fHG/eDE51x3x3VAZ8
xclYIz4Q7RV25AkY2H9JWYK3bSaUJXc2hbuDvw4nzxhbzD4D5PdvoFZYe6nMRAo8+9HC00wdUuHM
+ChtELaKt8QETZ9l1zr3fUQxFhlA3bBNJWoz2laZ3cVcOLQfvsPz3RTSl9PQRDIQAuKsjhzSfIFJ
BDFqnAcEv5r/KJ15mE8C/mmDxsXOLL7MCc/LjcWsBfl0xJc/yybDSA58nd5s0y+qRW/ncLrNuZ2e
KKZ8RcTeTKQ63/TDaGtXKS2usuxcvx3L9gPTWoSGAF1c3WgAKb45uYXXF5Bbyj7wM9BJAkYLXnn2
0lUxhxsnAJ/5bvLhNBFz1XylkzvE1uoycGlsMiGpl2mHMIR+QrNDPN9nDFtv/PA6JWEmX+83OI+t
WJMPk9UvSBR6fBnw0GUXvDcc7QwSThtxwPKv0Wf/ZbYrwQGFSat+VonyyNzcMCfF/gMakbECxONV
F+wYJj3Z1s2h/fsmFRVG9P9OWfH3BshuXda5vP4EjsaEC9mmzkSDcukggGcN8NnfhZJojQ+IK0hP
9y6xB1AFb24J0hu7Rgi1w4yqmTRtAqYKIER99FZlcTo51xd/HcqGXwKFrQNIS5qSMgzAT6hheqxa
7iK5UljTHYrqtsOJa/CBtPlwAq3Cu6FLYCzz9DkDeLkjclTvPvmu8uMxMAVQcd8ihEzB4HoBl687
HlGrvCXXDBLtrvtOPFVJ7Dmyt1VrbTMKFE8IY3QHRaDDfVC6cO7nXaPpW6KbacvcyUotjNGdw0Bs
oAqQwTWUb5EmnmAQoUay2NnWOd4/vaFT910/oSmqIP7+GVwk5pw/BEW6Qbo3nJ8MrLuib2ubhooK
Vc1abjO3PDJIyMLymNkXouC3QDF+iRk/HHEeK6f8nEYSUuM+yEWUvfAqJ/ILw3U87VWbpBE3V9d1
OePVvwIoWhUGmJeoQLH9i6QWMWQ2mxXM+t1TqM8aMkpdAMRWh4CjcEfp2t5nUkGbTHPAog8jtLAx
8SSTVo6Do4aU+73wLGNvb4QtGON5MffXStAludT4/JbzkUpVkBz5CjdmIVO/nYzu3f1efYcj7V7Z
/hTX5je74xk/PcBSe7isf3/QcGXpLiA5ZSlndfzsj3QIqfYs0w8dSYku3L2w5jKZSnKsRJ/pcH5A
7/tlyrFIUf/KsyMb+zTCRzfEvH0KrzphqBCNv0uvAlkIUegYtl1NnYdEHwXB5hLMRhZqDfSq3Oh2
p8y6Bxit0f/EQuu0dcNNpyhpHKe+b6NcW2W5kkX16gedD0mSMrAsyZ2FMQDKQ9h1yO0V2FlMlwCR
FLfnNe32MDoGDyXExlQOc0rzRs+m0ouzPKGVN+nOrriBR8o5V4GBJTAp98RRIz3y8gyxfFtdsPYd
PEJi4A551px5rc3NIfXTynWZVWSaV5ZCQUjI3T75JXmBlwTKK9vZIFCor1WPuXrm6ANSVJLA5KVO
cCkWdqm8A3LBnWXXkRJpXealBjKI1kZvSFVA4X6oltH0hHD88SiUAmp5cr7NFP9UtZRPXlNg4gcL
3dKnbCG+I68gP0ZWGqDQN1dZC2ipOVeMc6OfqGZ0AsgEs2x2pPQLcVsC/+WS1cyfwV+Qc+1ZYy9m
F8gAeQysk2dGgCwioXOzIOHgLULotkka2JZU755Ink6cN3bEmgDmd6ShpLahCLIxArSV5WhzMGgs
4TxyBpBdzwd9aXzp5bvTVMw2QCybMxh8J5GlMpPiLGveOtXvZAotRz4OrK+E+PbziFprV7G8Qj6G
PzocYX66qcgF6wWt9RRHPmSQJEKD+POHatgmpBnFuIwO3vlzZCSdnjiRklfWF3csmxZ0VJGZ0kLc
7h7LausjSRdiiUbNPv7BQ08TFqWWkjh/D26AIAB3EeLWW44HAGjntou6aAI0HcS8kOOq+hj3L44f
Mi5GVh3ZuyNoZDfeEii4sOQJnBDrIzrOWDTAXB7JJnK98M8RDWlRt81Z5fP8lesH5TMCRar/mC4e
g14w7aZS+ctSQS6dk5LDn5HmYLZcr2ZOJGiUjOvFpc+CECbyTgnnTd/JfYPbgVXzzpV6EYjMxpul
K7ee1YDbWMY6X5z1sqF7DiYBHNSMUCExyTmYyVEeTHZf09g+g5uM2OylWoSSrJmWLRQjcOJlj9HP
4YrGR9u9NxRTBJRBqiZjdZj0n+QhfcWM8P81APWb68PmioKx6yy8E5AqFvxnqAdT+oFJxiTLB7SD
X59xxxDlrRzgoj2CNDprRrArVr3rAjkG5wLFIu5543t13bc7DzqNFpXYoa8jZdbjmbnrc1BHYT7Y
FlkbaGeSu2Jy7mMn3I4CCxKdolZifywFEv1hbwgZrxlpR1DXjypgczHCrDUnt0cUV5AMdEmx1z4v
2mg2Qw6Stcih3gxTpbeUkA3jD7O9+If/vlSGSqA9pfP9TXt9OG7OXG0dN0i0/xwdN7K71LdULfZT
AKemf4w0xH8HbWY7Hcwt9sOh35sLWrK2kmyXG8V15gaifA3yCTxLGB9+JkK27Z7KisH8V9px8IXU
018DquAA6vTUVh65IQzZm85gKIRV1TFZY9bewYLEv9FUOFHny+wpgoVUFa9O7YzQ/LpLK6djUeLX
ODzZS2/V28rb8q61gAsfo6SbDKXWOXTT0R42OdD3Q1JO3GqAzsoGbQwdHggx5JtJXPTNGzwAxfkq
Ie7Sjv0HTwA4PLb3uDOL7Yi6PJm6d2/XoWBoFh82rPrtCXG+Z341h6B4BiAmZ12k1hriszuqgKpF
XVYLKfPYcUR4F6YsYYiIcx2Gd/Cwmhfk6SAZ/oxh83c6vF93q/LOfa9Dz+3rP3GFA+JC0fyn5KVa
7n/Ie64hyQrrPDsyCJj0AH0a4LQIZEPJMhP0Osb+A7lVZ75gIv/FCwgKNLJGwd7ilAgSq1Ytxymb
ksYm8tHfEFe8BqogcG+2p7p05WFGKOHy6IbysUdrxj5iqo06sSnQi+njeac+IH2K89OriHgLeAhZ
foGAml82NSZk+QR1PQshTg7XnqoXNpvCd3yjvhaoR3DJVk4npkvxKp4HTMnIyt17Hp977wEtXiZO
Pzl/8BBAhPT/+wu5kTEeUqZhUEuzTBqBJu+6N2ix3sHZrG7Vp+5DfD554qs5ZB1b5iO8QoYFj8KA
JByLPlp8koilAlbzdyR8Y6++IXzT9ZPgA5ma047lK3aK3jHEaN5S8YKMgT+qQD24x3C7bLPoBQYQ
kjVAMBf51koMU8blaP5euT5x83lESqpQPdrESVriGsCWQQQE1BTddO/CynoqAA7IM++XxJGXAWxb
RIPZEJiPZIM4ZDGVn06WKkhkPuFXX23Yi303E6AuasoxFLe7rZcvfpARyxGP8pAZELhFe3mvkzWM
OgerWjA3Jd+GWmsG522sQNDHlR+pAAFESQmJNlws+0EZHnB8xwl/SqKCjuMexN99ZECN8qXfSuBy
/AJGn3rUpJac6IRNXXuIpzKmHESi8J+OoSbLuRtj7Dj6BtSZJXwBFySgmEQ3wyWiCS8LAAzLIIOd
niIfNtKH0JL/aiVB+7tbd6GhkjD1vM/jSAyHuzSPYXTcwA0+NCZUYn1E+fjibwvrPnGRjAuS+f/+
T3LXqIUILIe+HaDyhVcL6J4VhnMVZlHL/5LjU69mSVeZtux/dVrh/uHTLMquPDEbZM2J9sAKMxDT
CIkNlOgxdnxIkg/l1EUjG5vUxhoknPd+VaP10rReVuDQ9aabQDPbq/5+2G/KV5rQofiuZYQsCKqe
Ax0X8/FmgeDQ2zi1uSK4TS0eO51sWx6r7QQX8CJlL8oZttD5V/cKNvTQtr89KTxN/vTrRysa2Qr4
kGjOJdKFqShp3muK+gv9WHpjVUZVv5fW7YFLGXCX005nKJoIwfKKxiU2bBe9L/Att9g8Y3uSjAt2
bMp++Q0R1ktj5MoCvE/OtqGTyGFGzcQtLc47x/aBP/kFrTGDGZNKDHVR7LSjLZz+zlpbEBYYoZdh
CicWjKpLazy4awJHzGoHotjuxR2jVMDgE+ucjP5ZsI/UGd9D15EPK1ldxudcuOnfXEhU06dYVjHx
awe5TsNnDhOpk44wHrOhkWsQSJnBmSmsriRulrE/vdCIGE4vnquW5+wjwkcIqNYAxfxgv72rtigp
P0V8sMHbt1HSaKNkQs2puzs2WIAUtS0jEr8k1CB443MYHUz0h3Gow9g8L74cyl8oW41KSlIGFUYL
WSv6WEcuF/NbcaoBHzV+dgpKICk77CnuXAyuJJHqBDDkeoYouqJgko2Qv7NMi5KUSp3xjo9uUe5U
06AJNCRT7yn0NMdDbu32gEGoTL0CmXCV0CC0FtMD1p7zKBmkrwnPEQ3ONbp/9U8uw6V0WIMGiu77
W0OANBkKoJMHLmxjpJnL3jBy7wyyfcKcIe8ejBqaHUaym0tYw80KluLzMrRC8EHyoomu8LfWegIn
PB3aHTZseTdllijuibvRzJ126ZB7F8ZOeAbVPMjg4i1qxNolvpJ3oFLOwLehOlvfK4h8+NQVo5GM
kTt4y2FW3C8SZUybtMpDMESJszm18sywP5KQGt+uxMn0PIREip8Ct/ZaN35UAn7X9QS2dVvrhPCT
HtHDkkr4iLb4KRTTetxVfNFNQKF9KHZPBYcLk7+4zItvw3zmqfnUNUSpeTN3CBwjuMXfPjDWKfc3
jrr2jAkOI7dY+jZYBHLRTgTSQxZHmpwX33gVjJUWAPpmMBtoWzid2NZCjmDlyjCGBpx5z4B24ySa
LUPt0zZ8u/A83dxq1xNzRoI5tKUfJULY2W/N7rIaib9fpd1izDzNPromrwLPUnU9zrak6j0DQ6lk
nUghihV28oglQG/dQA791vXFG+tB5TqG4aNiRms+ReJFy7zy90Xx0Y8cAIVjf6s4dQ4saIpqqKhp
6haF32fBSdygjfOY43KSANKsSWFNv/5dbQbhaSWu8DLnmdkv2j2CrZe09Gi76Ubu9Auc+2CMqGN5
Va2UO+3sai65as3XBycB6mRrof485H7SN3fuax3mnlDtxGwaaiSQXl+m4BYDuW553x7INDQTVMdy
hmy4FHqADoRQayl56cm9HHpITBLCPLmd24/vFiosE/WuiXlGXM3ttiTqVOcG1eB+v7xDkQyOIVJM
0xCz/kB1PFSQiKvTogDVgWzxsPUINj8yc1iEr8A8ScykIPeAu1khB4bF3mGqP28M3DQfbLvweGzq
rMS3hXPah4KqJ/Yuxc+DTA1jo8/7uAeMnjNFPW2YakTNK5OhWaMsuc5HWVQRFF1CFR461Jrc4LKf
JVmtCxD7YU+Jhk1umzcYGU7hnlBBSiDVdcWhxd4ts/LhrqzUosxC1+nEH65YmNNuR9q6zVNNtm8w
SD0C98Dm+qX/SmFA8P9xEYSaLlI2YsssiKZy1lzwC0N+yaAJd934qkvDi6J3lXxKWTZlrtoS0RSP
pFveItMvG2f413UG+8M2OSwjNJuWosqeveWUb3OQOJSmlVqfA560O19py47pAtqkZfe5laYWfGaG
8HcPyswO+1yASZwEktdaDTRB1etdYu7lFSCTlrM4A5gEl2mMEfWSUv2yo/4yT0ulUGTHkQqmv7jw
2pvcwtUEtSazwSXMSZJtoz9O0F7OifBfUSIh4m2ifYXW5shKclUgEuaNm/am91TJjJucCkA83TNv
vb7HYFmM9BsCgVTt0JBLmlb+dY21vzypSNqlOLIuKh/+KOTxl/jUX9nHEWNGL+CUyY0mFMk3RZ4h
0g5GXRI7OeZf2W3Ee6N4R/BAlTKtuhVOqViL59/Kws8EypF7uvzrrY+zVdq5CVsZ3eoKdNnTtLMV
a/SYwnyU+5IYuqGoXqoYxN1JvIc29FyGLFppbukuyl4ocLPoUQ/R4eOFR950OuBXH3BkG7QOxUGq
LhPmhisyONSXawOeHQVJca5x24J2Q+ZrmJkHRkak3D/Ig6HffgwMLkD/hk/xobr9Xf8RH4Nw/thV
VAFEratLd2iuCwHjVbBHIMOLULPueSQM4MpUpB1ZCLJZcsYoyx1MgCgzSLl2lajD4o9hj4NKlQtP
ScxVKtiUUHZAu+uu+wHMSpJmC6I/WhZutxIF67FLmIvRVvQCwunNUNVRNuQ45KhYM4hDIg2HY/CB
1Ol4vn0gJKKOUkq/qrGE6YckTm0q6ZxGdF/Wt++++IWalHiY/yqAaIEpOgV0RJR/ol98dJfTs2+j
dVaBIrV9ixamCtwAIThwC0KE2jdmrrmvsVxdvE5uVI4BwRKJUfIYIdcBMMKrcn5UlUyOviozqePK
/sqcjpx3TzfzhZx7hnZMTKkBzJNLhMiwG0Dj2mXCchvYMmMDgIQikElUofqY2ilmZeHHOP2Wf3D3
uCotwPZJCSV4p+vsLFLZIPViBFiArmJ0OebwxmbpLyN4sQep3ETAVUyoI+RHvOJeKUrCnX42tZMe
ae72VQEaW2fHL+bJdT4yithKyaMkzOaFY4zP7htmIPmngij4bVfnnXXo42F7xrZJzGitjRGR3/UY
7GNnri16aTN398SWDdAFOeTu4nqjRrTyIE7ffG31F+/9K1Q9Vjl4Vj7Y8NiQ229LVLzWpZqVAeoJ
YdvpJuFEeVyJXOrfrKQdcN02Ar7j2KB4ARS84DMQb09BQL/4tKjZhOeeYK7gm3KnuscV1uyGQNjb
Puopw8WEWtgu71fvV1oOE+mfveJ/g3Svwxv0YCtPsCz+kAC0Ta8fbpfPU9yYRqlCjnpXlhnnNZ5c
mzhC2DyvV/K+BN+Tq6NpEiaYND3kuaOEYI7tPLbnoP/K1MgCKB5oW4ig2UeBE5O0Ba0bX29oaGsS
5qH33QrJHsgEvVgAGbbD2VN4/u9G/9vlRCIhtv5IWy/fkKf8MG20d2OOjqqQ1KPe+ge6HAgvliFZ
dy+0/kAVjelxoKk0esVzVFSm5kqK5kcCpA3PtvFo6eFifHgOzsOWL1ZToypAN0buoWuOiu8S+1WP
In8TYzZihnoUYBw2DFjdT6tiI1RAu0lGdUFxAIUgoiSkoV0ndRRryUhlbYzycbYIR/kaJ/bnpRHX
u2n3yDrK9c1iZXmNYL2g6+rQIMrHQsNppTtzz5o2xCJh/VxLfOTEIlxyKKklHx0TB5KdDQ8SVd0i
by4uxdnfXzCjxsxJDic10GAUJwQSMuhTs1kmUtI54P0dt9/aiYxVilhb1151ttPmQe5kYJjmnpgl
pTw6qnWBJO7Eg1Rqwgp8lXNmw9BAGNynJAuT7lJulJ1kdrGUt4OLqssYnmjVsZMdy2w+5qycrneD
P04LDp6fEqkl1T869HGB1ojcuqMV0MNvVNoBLaCbVD/ablHA3ch7gl+SP2qX0o13k704D+2d8SBB
Cqlubk19rs1JlcLK42WnL/RvPFzu4TPI3DVf4pn2hMB1fL/Qzy3bghJV186CPPe+BYqCZgZhbNzu
GAf5fb8dW1n5MktI3SRY2fqweqn3BusMfwJJ/HFeDKOaSLC3QyKJq6rMSGPxybbfrErApJxw6MFV
yM0P+DOwswJSGGEYdKmQCSnOmVgyjb69CHzzdRTBbTuU8dfjJPYhOR80C779baNjZtchShMkW3Ea
BhDiP4GkcSjzTSidsL0Vxt1W4xV9igOS3BJXBjXRfzKiLO7WLSwPUZddwCECAC6j0y06Z1pjLdT9
lzuPD50OaQstfBXwpvef+pgwLE8ipy8EOJPl97mIAa6L2elD7KgxXbqI4BbpeWY2WC01qlfvwgKZ
li2Ael1cOWfI4A7Vf2wj9ZeOdLkv4cFsXOvnx/lxNnWyR9VyBm5r0nBCvvvUA9C6wxtp/jXEGz7r
FITesmoO/mJPiPA576h3KZ/gRwwFfw5qwLp/m+KBEYiynTqObfJo9H46amdLGpaWOZYCcW+3A2zY
0A1EuTtkF/hBMcAPisnWLSLdyzoadbmnkGKfrqdiV/sBQuuxNNmeSMScFlUXah7FdstT5J/nZr3f
K2vOA2IuNLrLCpSIHw1t7BOM92K/sOu8D9F7ARbm56IiW9zYfFIKyERYkdRfKDCF7XBarZnvMTGB
ZnOAusEYRCpGXO8lsOWbIxJSkn+oxeDviObkVnmS0+uaxvNmDdM6aTNVJ+ufZwwcvoOy3lH7Rhta
i1G58pLZlszRq8CLaX7zkmF9SfbKtBd9N71mEXoCa1v2pkdPcCSsSxtCm7aaIxQ7Jfnnns03O8tR
Eut00g1gFwkkCRZNZK6GcEUG2KO+q5+BTtALfoPM+zwUKF/dawzTqbCK5jK66BldiuanPAE2KxKI
Qtizabjkes+NObIEevZ+rq0qIA0Tym7gpCNyLgzUPwmgZpHUvVlCZFsYL/+vqTeSgfEXIWfvPoFf
32KjZrgnX7qW7jzLMgPJKUHzgTRXIGJTdrr50VX31HAUjECVRG5a3RCYzDAFDF19aa6oI9keh/en
M+Qn4fjPp/BvmPGYPKQg9YaQlrVIqCucMOAtux2BBPV1djZhqF1shx/CksEucMQgdG2Y0t2ULoec
8odfE0Hf9aHkQhAV7lPz6HIRK6Emv+xsLac0hXVsQvs2zVLa6RQcV2CcIqWn7sPz7aZNazPGQtew
M9u5KqWpoFGZA1d0GI7NVUrLKI23mx7bS80pWKyMa5U2M9Obd2PgGAcKTLFrwdVswlX2/4l2inSq
9fdJ3RFP1tGvhVVm/h646glbRaYKPGlg1YiiK8R7bouX4nHdSuB7Z4BV/8a3H1ct/GZWm/2O9eKi
WgypeQgQuXjU3IDpxG1yWfujcHoFPCFx8md2aLG8gFmfgKT+Alujyh46cVDwOMV7LZl2JVLqoEpU
f+hvBgZ2DQ9XOhBnlW0NAew4BtOhxmo9zDr8bBWpKORBk7MY/hIiE+VSl3gn2USoGTqxVUvj2JR9
6sL4iubijDd1fGJY7otcQI9NuH7oCx0U28++qEmvjAFmjg81gKkdmZxucKnmV/w76+9BDL+9MDTT
n4i3L49a/nX3Rk086jEXrGmU/RK6WqWTYJSjI1aoZfRQnACJmlCOiNvrC4l836AQ7Cuz+mdu8kVb
YCgsJh3Gcx/nGmEd5mSNneLdJCH2S/rYugAgV8PzUyAP1Bix22+2AGwAgScdxrWCl7dOvtZ2K1df
ms4dBPE2z1IR5cGYJvYaDt3krl/WAljKhhhfrKiea0+b1Ipq4DpHBN0aMIxu94ic6tegmSZZY502
/SZIUrq3oe+MUV/ssY0uV3vrHAnR/awd895h1LAxUmG+gDXjNVnAe87lWcXmiscwRLwgs0AYC123
7OxSl07rRLW40eF2A/K2dav/HJvJ7uZ+7F+BbXzXeUhxNai03/05lmsTfKqxNm94WTG9qE+fAD88
k4ZqBotBB/j1ghgAHv7lr+wJ3N21Sb8XlSY9bTQRSvBIREklS+FOXr2Q6JmvcJNG9FgQr0B2fpb7
LMiW5Yj8FmiBPDxZh6VRxv8UAVv2dyfw8u14pM/0TWTawypHZNdf0SS16YU0+eLQQU/EdMf42i2B
6LUhoWofUMA9BwP2bM/4Tez5M7MfMqisB2vkqt3xhKgeXR3wzrC0wAC7S9hCyuJZ0ml1lDuvLsEh
qGyYCtZvzGy1DOMH63AWROqldjw7c4PXzIWJVL0jfBbWQSoX12NyJQF+FxAy5833wuLXPD+PY0VC
+vkuSRRZAE/23gOJ10vqC2Rzjvq+Cy8Zblhj5qGpts35vLwJeyg4yh+ZHYsYcIcFaqJ2HMjrLcmJ
fQFUq/ONu9sb92xYnnVFyherac7USOP1BmsSemqWhzytWQAqB64mZE6utbzvjC+FgNJYQeuiSs/I
ZNiRBseqdyN+7UANgwZPJy4vACqWlvxHJBvGbt1ZpcSzGrT6DwS5Ux9YXG+cYeO24rAlOudNHFe8
LapDqH9VMVFJsxE5+05pxDbR2LYb8+B2WikQzRR4TqDnsEY4cZwOPkYpNbbgWx1BgoYYJIYYl8fS
zLVJaBOqMgCIGPtir4rO7Bss994Jno4YJRvajApZnuAR4Hf2iJSUgGPZjugZGzLiLFBq2MGENlC8
OnK1PXH1dBgVy/1gPJ28Buf1Wj9QkXQps3xzacsvOXkLPIRCZRQ7BiySQl4tENQOy8fbSqC8C+3w
MsLqN2H7C2DRqHPLnzlw2dwD2EK3edZBfjz8EY2k31jkEPeKec95SPY9PVU9G1x6FXRg86FUZmPO
wQJgMEkw196NR2EkNiL2mnSnXndVKbvfjpkrrSowOM2q5h9BSn7ouRH9PdLXFluqCbyplPr4d88l
PYzgvXZgC/JGPrs70KWaswRmUFJIgK8ehXeTQjWubGOAkQQdFdAG2ntdAaaoak/YFzkCzaof3Ato
9xkap98GabVgZwHDqeTba7+Hy9NfSazqaslcVABlzA7qiODW6/56pMYW26bxbUdemerN+NpykMDZ
rvAk9Z3vtpIcpuZ/fHHBZUuNy/vKxp9aWkyrcoiEn6EfixRJyBABWL1Spdwaaw7AqeO26Wy+IEJP
lur8vSncjTULHqqIs+iGSc3xZkdx+tG+6TCo8uDfEqXu/uyatbT05txJ3mNTc6r6Y3tKvn1welUL
jwRm8bucfHKpAzueSan1mZNeFafqGhfdREez30hmgoQgodWdyk4gVUUSj36GBvtPD8oay9eP2G2Z
mcCJmB08SmF4mgDxRuAozfMhmlLFBrCLR1CoAg+FUYKYCNI6oCG076Qv73NxDvRjdMl01ibggmEG
6jSfOMCbs3TwkheJ8G5+uF2XbicBLR6xBsEhEYk07b3tfeZsANpJooQsyxZVMsGqA1hsmrz4agIT
vCe4Hoc0mCfJRDKqMT/uyxUKRiHWNwHNEwZFV9ol7kU/pKx7iHEOHK9DS4h3utiXiO0CvuugI6xG
zvZyEm7qtfpfO45BYn3Y21kQJU5U4RS+SqROL/pzeKmQcfNbSR95sB2Ipxw84hLnADdv02Ycvemh
C264ucP71ehH/EYGAuMeTUOnpIZ1XvPd3yQIdwmNUp/uzBOjQm3FmNSdm0/94At5Ba+z+vFfWJfS
EGzFtK1iXyhuTjm7+LuRHkLp2TCnXGyTTeMSo77wJapusvvJTDlOsWF+HeVEeTg8Y0MBqsZ7kDYI
INXvB6XD2J89P2iKMaWiaqjcNiQ/KDNfY6coRk9UZjheIJzr+2/BOnQlxOSq2P9FY+DfQntgg92B
afdkT+9p5JgZKh95UdRThElzN1VAEJ/AVJCYh0o+R4hOXpPTXVmbeQLhEPvdSFLac0Wnvl0LjOhG
PcgxxZrMdqajz74wqZzZH8VF7D8Pw5xIC2tW/ouy8o7ixQvC1AvsJuBglPeoGJ1iWYQbqMK72qrl
Z1gRzpqSvO8SIyTL3LS0qJrodPNyJnVU8/+tGnQyw2G9x0ZWikG9bEfbXhwKeUYMp2QeRRFRdFyC
CnxGBvVorcUB7sPLmDDUhMZMFycQ9xmQ88yAi+qpdfbw5wWA6VTBVznMzOOFXtfoeYZbjObJBXJk
eSM6MvbWXEPDwb1FGQjEivNxDUEjqbpPdVKSIYFUansREOesKiPYVWawHpgfiqbVE5FB4sWzFoEN
a4YqiMyLcT89LAUDia0BkChOI25kHYGmM+kJh2G1vWenMZpb1y73OVMVzqYA4m2rlewvP4KOw91w
V3SrRyHYOi5fOyd491EN9VRgvMLDCnOn+XNnsqfNCuduo2BwPTrTgT3kCd2i0FlPwsa0huX6zL6x
NXVmshZCE/OCdnydOLCbhmPSB+6Cj3W3eWlGALrOVzDTyagzauWuNMhB+yJAPCiuOKwZoTVkQ/re
JVExwsuLA1EP9XxK87tmXQk/t+x/B9gu+G94/U6qVpbgfiChahnmd8YYr0fSYHYHRMfP9noWHkFT
+278pSVjNXXq55k/wpoF3iaQZvvr/QKZqXVOVAZkPvfcC48F6pAHaUFQh3fD1fF8inkd/u7tAcW4
HERFvs7E7DUNJlfOsi5I01RbpcNgvYBiysAYnFKxtRa8nbpbkg+jSd2rvCuaqDUgBz+gSKR0b5hv
ZYNQm6XU2g59whzjjIFFJm1zO2CENl4e+C3U+5exepwGHEmQGgMqHZT8/YlCSIO3+lSVpFYtM+IV
S8oMEDAAj2jLqsGE83bB+1dOqbbVRYEveOVfFSrTpKP4E+puTSMmdEIeNp/lCopnn6mufOYNSdEr
WzpcxMOYsxGhkk2NqIyM8ChBs4FjJFNJ2svce3Zfg2R429lpqgF55C93A0h81jnri0csc1bhycsC
4ZqMNGsh7TGUzmSJrYkaDrvRzO9vtdz4mFVNVOu/rudi4WwuQUnhDHMc0P0qzkRGMCWrDldo0ujR
SZE4n4+ucPebPzNWcpXjyXp7JeI0sBEIoCR5RSek7BvcUgrHAdRjC1L9fJyaHCtKR4OgZ0AojdtS
HiJGI8gzrmVSkFWMJNxnYcIhdSI9MiiALKeoXWZnB0qeHddSS8Rft0+uPnt4n37vGOus7R1k6Zah
XFlNpGVb/+xcUntwuexrRp/e8yox5L0rnv2AEYwHNmM4b7vTUXrxrzYKh08+AUDXnRggHmv2IJ4L
rmla7b0EDsfG9on61rItJ11O3NqDE1zp2xGqZDs49CyMRjmz2Y9xDaQvKC1/XCB8DHvZ70ADbixf
OW7P0tb1ovwPoIGB6ioIXAhPVmfdrhgiv8jpxUMANtVbURnh/x8/fDva22bsSEDxVhXxStmPbgNm
pIUNTQgntR0jBFD23qdgHzAi0/nSV4ph8gyPy6aDpaDmwls+luiD1WCvqixF2rbBRgRvS2u0FVyI
PVyOFeL65MWERaMCSLOslcf5jLT8EHcVV1oQEINnnXpr25/2rQnP+4WnhVMtLnNq0aUSMFqLFf/L
PN3Ty/3+0ZPqT0qGAwIphpGvmdfyPOJGvHeHuYc9Oe3B7oiYCFicq0ebPNfPglIZGVuylec/l16t
6++GGf9Cn+VFNf/ExSuZYVUuIcENRRpoNrYgdGi4remrYtsX5mpFR8iCfzn/3PIqui6jug0FEW2x
z9nrBBSxZN78ouk35qG49ZL+J5CSehnco6qIgTlb+b45/Ve1mZYqNPy8Y6irCLFqfCd+q3BwNApR
iKjrlN7jKwfivneniO2hIYtUfoNNqypVqWzMLg+xYGdVo/LZ+Z2MbY3ByCIrxe4ctLHRLecIgq2K
qL2QguATOz0kFKUAggkBc34C5MQcJfQS0ByzNdFNuQLh8qBi8U1CRwBI6biOWd8aiJfIoMjQHthc
E6h+Q6vCeJpQ3bzBvPNeMutSI+I1u7rhcusEW2N/ZZSVfdHWNXCPCWU1orJePnC29QBbD8TJQW2M
Y7aAD0CQvSQnb06ihJIUIX9JjNzn/VOaSelJBsnTDuMo7rleTjiIbMV471zhcvXxoMG6oBxireI6
/8vKzKHk7hhLAaZKRP3QuJU75UWve+oizmf9ayxKHyj/lvTjEIbfC1iSjiU8dEaq/I9xY8yrPy2l
4UcD8GEuisRX6fEe2Nvl683N2OTMqzM/zcRldeamcDN2H2WK0SkMTdxmKxaC3FZ8YKjAHbK910wZ
zAZhZlYFXZXP6Ixxew4U1iiVd6LlfWJEvA2EViNRtNqbIY9FL2gxKUeWh5F2weCouk9q1QG74coB
kBWu4LV3rcEWwETVXlAu+KS8wrI3fLvYcTbKDE2LwWUr8MnJ4CqEufXwvZwYJflkaqse4olWnUce
mGA2pDD0yyVI2MyUqV4wlrC9CDvRFHxCGWSytDeL2Nc9iCx86wYhYKHilyZxwC7wfyTE5jk1jDtE
8FPpnA2XMtxUBGQIReuwzEIjJ+DQu0XAJK7eXpuORHNK/HbisQzGXGOb6WzGe20JPFE7DM1GizJZ
RhaqUYzVOJObOMg3bq1hGa5I2gWns2kBtr1J/fgosh+blAChNBd6XgBDqANy9kWjiNxkImpw5Ye0
x0mn/0tQwPqiw2f3JimPD7/0qtVLBVSqsi1X+bbefpD2msrc5JObnL1YQ38M7ttDnbYGtQIWtrQk
0SrD32kgq7PeCo8G83nGIQEhwO1HhxT6Cpqq8Y9oGbV3L0rJzoVWEyE72AxQw6BtjsREIhl+Hb3E
JVCa1OuGgYGHndE7WMzuoE6CIRBU+QEN88q4ui86p+LqiUcFPrqbAI0HvsjRurduMhCB5t+6ZDQv
1rr0Zit/0vtM3UJLBTvJie/0kTLr+ssqI3ZwtUinMnb2zYmbZrEUzTfgmQGOEU6DXtnFlHP6+DER
eSOQDPU+NJPiqKfwazj//yJt46iaiTWRgVt2KsAeB4OJNPwvOxfIgexLdBsRSyywNDTeN+yEQM2n
KPDd7hUni9htMlE7OAbspfgIkCtJDoHrrqH9ZS00MdrJ2m5+GVOrBKrXAgeTQx/SP4FF/7D9aZ/S
ozPuy1zVuVzAfmxGGSw/tsRfFTsEj9wiSxpXHCzUxlLWQYMHnyNOlL0mtJFX0m3/XSHfTyLVy5fB
gLxSQzBGcSN0lsyMM4JER7AY83ZNTl3gfr5dedoLIIx57dgKW24Kjj8CdEWvwXcn5u10IrPfdBxk
wSHFABT+qPo6/eLzNpBTRHOnx8IQefjsNXBPt1uDNtsLExgSLzKYKHNmosWNqXHiAQlBTScP72NX
GRiM36+hlGojbD4H5V7aPU0ZCCoZrRu6VZ3vQgUyvAvYlFqfgIIOLMNlFNssX9aUWfCz06CR1H02
mbnrt5STjrwznkLwtJMmSKps7S/+Z7NA0IFJ39HQtFsuRDIVTRjLm4jamjtkD/YmdRqc8b1xnZpb
QJpFLC6Y2WCQRfIhWPUBEaUBl4Ug+cNS61TWgTMI8r6+ZtkPdtZg0ZVn59obV/37Xte9Yti3eiJR
fwLJapouysCfKoly17IOHbbYmJ5SdrZBPbttmRZfXLKryK9/LBagmFnu8BlzLZUseoTVHRpckuqv
hLH67F/hgubAaKnP5VvERlZEjRpdqIvWc4PaxibrWhbvvdteVAWiY7ceOdLZIHFxw2LNiJjhv6av
pSoSLVaBvtJkw+9Ub95GJyG6yMvL+z0jpWRnY5HVh7vFYpgH1O8iQg61q0PlK6KQEHDJQ3ax1tv5
i0ITIk+/a4JtLUO/SrtRRCO6LIBAneyFtR5zo2bAASSyMN+IcS9ZnEphwmgVNzpOqZVC/siSkJf0
npqtgPtRvTTP49ggRoGLA2r5Qv2L8hf/v+bu24FiM1kOqa6b12DYsXxNfXRy9s9e41P0aDS9wgiu
uicFq5lRi+RxwHpC3OMjj4YzKpKET6dVqsxYA8YS6c/MBt9oEvzGfK7O3iuww87fzvSaHJMVbaFa
q3GdtU5zDlAXnbFlVS1Edp0bQ61znNsIhjGHS/mFdhHse/3livQttzwC1c22crkzN/Qo7UuY0/2N
/BMHJrJJAlRAsHUPn5i6aQ+jJCqaCZX3ycfaKrcCW3FaI2iN/vuUzU0/kBIjeW+dBTtb8n7M44Ok
O+pXmVtx13ZRRDJioK87x+XSUq/PuhelrW3hsT6soPsb4+XBmNnhTzuEzIvM/ohz0gK2dBmM4X+W
SGlnYVfSugZGvbrU8kEfuMw48NYqVWC05SMlMU2yJDETIpvTL7IE1/KB1wo2Tdf5gN6dFqsoEW13
JcMAQCySB3NOKKypBHold/1OkFru+sNTPNZLdBtcWlHjgk4hyW7TfKVKD8Dvxn7PHBEc5zNp27UG
KM58TdX7T0kuKWB3Uw9dSuiJ3Yj6SV+yfByoZ8/SvfdWJmAnRSbB2hvuQO58JU8fCReVCtqVjqvv
bKUwSglesmyFF+eTOramYQ3NZekqja39Ao1q44oVX4GdqcwuYQPt7bVg+bjdK9O+iajkYg6vsTa9
YE31s+e/dbnW86H5HSI3rfzdAF6nZ8xMhTw0jy8trvc3AClrR7p7eFpv/2IsTE7LxCw0tuKt2Vy9
pRimZAqhMOgMOT03lewr+TiUP7WWcQUlNd7dcQz9gqRZGJ7BbQ+DRpvHvf+aBJ7myzmD43xsTXue
a5dOg23YgxSqoGbWPpiIh4nfYANzIRHBc+Q0dX7tyIIcBj9LecTbBOxOjP3cgN96WvzTInxd63ih
uFfaWF6CY7J9o7nfMm69Zr+3piwRThrxjltHkSF7Hp4WwM9INVFcMBh1e6uimFp6M1lDYzOBp0AU
66vP8hCPQ4Ha7l5NBov/h7sTq6LQOuKnAZrEyilHoAeGRKGUjyOGWImyCNXlocbaEjEo7/nvUG2z
EoEiebVA+6nFm4Ce3vc5bBEmsLmDuiAdHsp95du17TauSG5qN6SqADr1+XNoPwrksTMzvxgzB2HP
HowQ66ACWvlL8iZjOjPBQVX3MjJs5kxVpf2lfbbsxS+Rrtxxwcjpfnr5RIm7o6ZBz4G9dtBhSqjZ
MwVLmfrA/Xm5QxrKHygfu7rD7CznStSawa1TDhYsz70DnUswhQp6ZbdMokYnuVOYtk36iIKbun0/
2x0zOBvMZE10Phf0QbT5/vyAclbsU4dyOkIrduJtJZsOZDY58HzaOeTfv+3NSU++B2NNnsEDOJWs
1qL87Pfv7NolE2Rb7QQSoNMRuSNRtwT/GXC2J/hLcd0UB2TV2bnJvd437+cmK+ieTTlrxAerhlg2
gu5NtgclYZevOA0RBMft8jEy8yLKrUKyJOoXYSw+vpFhPo/7ATIG7676stoUdhl0nP01erV9JM7l
/6Chn2ch5fWiI+MyyfVu7T8J18FubpIy5pLtfhTZIl7G4CnSe8fsjclExzHECjAG/fa+JVKCdpBx
2WDabt3giXyT3ZUxZDDtO7kTKGSOr3yyeUJ/8nXqAgsB2UYfbnc3WbGyP+ppahg+3odUO7xgPpp4
FzOxgH3/el+YESM7ggew/gtNsg/SBd16rTh/8YtCARyoZ6kAk0+DghpYHUAwkeZHqm+EcAa/yaUG
TkEHGvXA66k1zpvOpX21OuMurmCulqh0djWIqQ3qEZKA/Fj6V6RWQ5A/evqjhW4hBofH9pNnKjyg
XwSBUgAZTV3lYN3Ho8+bImrklznK9/QYsgoXjJ/s2F6miruX19l1F4k21MhK3HqqSHfr4GQThmxf
EKomMM+v0VtkfSEM7FVT0y0Myc47wJGwKWvAiSIHUrKh75vvGT+S8qstlPzH4OLQ+lnbaC72zQX6
WxP5Wojq3A6EQ8bGVZhGz5VVdpoBgLYT6VZvNcyAL1oLbzZjEnPnjRfmS69rbK9/0TsjfbbZGcvt
iGss1jy0p+lAH+DYmNc5asOZoWYxNpkOw97qw1PDY9YgYiNeI7JZH4Q0zafQCzfNePfNRfRVGjS1
sJ3cKUi77AduysxH09lbzOh54fB7ON8GmfrPdse5btutaErz2EXzVgXrI9dKe3wU9vXXm8o2zhmy
v0WIjnyk1808ZpC5GY1dvYugGw7ZWZ/aeUnPMCNh5NqObopUZXZH1s9LcgYG16guKOExPjZoD0FG
76FzQDwOi+YY2/86LHE1XF6eWfIlwyVbab7i3/lNINx1KjY5gBs8NACU8e20uD/tOdCZa//BH/ra
lleqzYwYcP+JxhW+1nX2PuI54OvZivgvDOOHNQGOmy6RIrmxTdahjVTCrAnYnO3hdxliNn7ZMa6L
3eLN9ImspQWeJj8EJ31GXbA213zdNSUGKNPuTFMC4Tr4WBOXfGhwoceBjbOJIsLrWDzy5EMxvyib
XZ9G8VeI7GeIdDS5gNa0Dk/9CiPhZ9SMMnCSxW9C8kaxipUPqe7j0xjLG/jgy9J+ZaGR3jtkRG6H
32uyKosiftzMFKxK1pSEJKw6s7UscYttQE+7yZurXj66v3kQHgafi+4KY8R/VrpLpulDMIkS0jo6
hQpeGA/YBhZ9WtytCPqpZBF41XYCVF40azRRtrcI66Pen3vw/wdnnqVLQ+CFx4yWZmpHDw3r+nfj
e8vbpN7AOgRT6sH8tnVNntbFMfZgXIcgqg0ITHxhi9CmME+UwrBg+fJLRHX2vfQ505cSN29j0mcG
FD1qLVEn4HY6lzrWQoCo/eQhojqFTA2rOJ6Ou9jZwzWm6Hy1C5QmHijyUWOk6hhA52/mQEfiETSW
h4Ur2PPoK26R/pVasP5wIrf33DHnhLceB19tUOls1d5lby1WltqRJNKN8pWaacEDf5y4c7/ZwWvc
TwDSVsVMm14LtrwmfLdjspD+/sXXQX+p2KkOMKYSkj+gq52pIDksa7Cxu4fDG6HzD+f1j2Ok0Mb3
lrrnv0+30SZO4/IDShkpqfpBoTE1gKoeU1LvZRr/7gX5hfGXCWKOLknf7ZlsUQs6KXB3Z0Tirw9Y
106tqUkqRWO0iIDk34o39rvD7fswrAtoyw0TJQGD06HCt5s+ACgxuocvJ4LyDicilnmONi+gLwuJ
DJCs5NA+LrPG/7J8uCT2ZAVvZ/YgX8bOWDtBD9QPeVb5QCsCQx/pDcmuFdY9LoaGN7YHBVpXCQdH
rwjegefiP+Av/pghXIdPLzWFaHICl9a4N1J9lcuq/SZBlumgNx0tcWpMcdlu8dLkQy6cocqoIi+T
l06dWp5nswcGvkFTpzsCm93dJ/uvlh/eujDm9B26DjqoRIMUMAuKMuDiaX1oKGisVTyrDmQhJ4YX
aZe3XhOxh6TwGOjxuyzbmseBgFBgKerHjPLi/XIx7uQWbFIgxVonlAqLbkzb6xIz8nmZwHEuRJur
QSQqrPmj4ONmn5ka9D4NNI/dllxxxMMaViTEF6M1O8tr2T4pUHuwZ/ZaW1ZiSuzDJ3ekiqsezsBS
zqurrtbsCToGryTx4cAQ9VAUnMS2VLQORjPs9jj5l/JldLn5GZ7mRg8RZyL7lGCNybSXQqHSvKPM
5kj83alKdxEbVzRtR1dKhY9Yjqtol0Evw+jUwHt0kYzxkbVfAs4y0jZeX7H6Wnte5YzBaDABE8MB
8tSVQIgCSOzGwjuIhEpWi4th6y8GexB0HWmtXLbq/9BFT/PkbQPLuP/rYMpufUHeGjLbiErKx+E1
pUadsKmMaHf8kxuMEhQBjXpt0o0Dud6ynnEv9sBtajwRrok9zZpi2e4aSydyXB6CAuJipo7U01jw
yPWzBpQEzFBSATxNcH5WR2nZHEjTPmywSDRl3ZO3G9zGLCWduMJnb6O2Uv9f5otShpi4JtjcaCST
5vYEHhBhJ8dt5JZDp0mbMJtbKDGxW9HJzih9jVgaJJQtlM2tywWmfXaULw+s8m0nm/yhY012Gn1u
mIep3FCfqakqkwCs10l0JcTRtGbNZU/MkafNPAiw0FkXAOABAJpwLNfw0Df6f49yT+9aVM5+joMI
QxHy0TJtoY5LeTMufqwsWJg9DLQHaCg7HFKYLqqhvuvdIoBeU/aIk9Wp+4c7VVNqLJwDCY/OZrpK
wKkTxvupSaQjVd9QVq4ZvUkNc4oVt0+lHOGsmPkrU4ACgrGhyKW4tF2JLm5RmSBFxA9MU2XxsYVT
gMNX7Zj8VAL4iPdZtd0Zh8h56MxiOyAzYEKhytw4sXIjflMi07rFAcjnjpRfNWDH1xmHF5xcXYIw
2aYskISC0skkV6GlTyZDINipgV7KwNawPZCD2tFQ4JSmeSJ+amXuPC9NvgqYKKFfxEgiHLRdw/EY
C5RJS8diUsJMjDhG3xEs8d7aUzl6AOp9WRmlUXlTMUMkpp3Az0XNlHIj56KLLs68Z+WJE8Fg86J3
To8FpvXoru8wKznku974u123xGeJ3+IN1RCfNNURV70ykjWeJyedqN+FpawOe7ZtzQu9zTekg+Lz
rmVCY4YQBJIpxDE+oR6oSNaeuaxFV+gTRu6RCDLvby6jobClf1HER1b0nKz3IhSscMsq6BfaC3ki
uwT+6vqGbnm2e9kICY7b2eLo0zWA7Um2PmRieGgFkwUIPBWuDYCPGUNl8L/tFvSTnZ/Xey5YTzmo
EsHi9AopMxBmTUqeXS2X7ouNFWqBfhNtAJNnBcGS2tBsXRf4nCvqtrQDokpYAPqbyJ2C02LpvpFU
PasNKSdsg4yHbss8pqgT8U3SiQY0d/Lf/n80bEg34za4rt3kX61k3Gl3hgy1isb2GN5NsFHddSex
F0Qmo09xegDJdrzUmyXjcsKggPtteyFjjqvhaKWrLV3hXD7kNqrwOWEw8nR/xEDWBoLtSA4PzVfK
63h1A1aqRSktTUbVdbwmtN6nsSWRxU0YHIkqaleyCaR4t8RFQIo2XWxypHUVtlnOq1ijsTOct948
IjFZqYPQZKgV82ZXYP94tcEY38sLcgIx5BrvSCw+yHOBpmUlY1jH5uehCd5QKPQtF9UqfnRFs9xm
5A9j2y8BAm/P5KltOvnDldU88ag7VnYTZmgJcqxqDiWv1OGTqZjstoITr7EYtClrO55KKp914IwB
hiwB4lfvJ461WCpD41YzFMMg65MhpOaiTJ5WOsl/VGSAjv9X3jjXvcjXSprWREmY2l3LVPp/qGTN
PbTzWY5sBUzxAcDV/gzqMU2P/GI+O5R5K8HJqMpnjB4HEM0sqY/6FIRjyQ/vk5nP0TjQoQTZAJ/T
PnuleVOnySsyeKcWZHNUE0f8spfNp3gTt7kwE65fAByFSpTz67HgL7jgCraeLe6TME7WarTsNStG
HjRwUm0CyPluvX+6Y3KgZYY3R2dJ4BNb9oQUt0IiJ1m2VaNNrSNqFud4sSh/1IbKW3bFKCqCultK
YD0BWAChXmNs1+8QtR7fIGXS38gH1KxTNizEOoxxhJfkjSsYdktqN3sQ75xKWVa1wNnTiVtEhPkT
18mW7Aa5USsISrMCb84IHw5Su5zf6qbp5BhlBzgCM/8coTyOoeMeIzY+JlaGtZyVqt9/NLOHxiC5
QcCYnV8Y9A+1qtm+mc8HVR1y33Dk8hr9ldvgQF/TE4HTtU25kcM1OJEwyBuEJh4hNgRrrrDEMQkO
Oatb+3VbvJmeh8++LlocAtwv3R1Ri1Mv6f5uxpZHTAp6gt5diGYBvaZkWhmsdoW+lUKuL5P1zfuf
oR8Zljbyl+uHA6zLFNqHrCpkeeCPau6v5+rETkfBgDR39rqkVKh1AvDrgqsshrcIO2FRnhm8Sxwh
YjY4QdHPHivdCnN7SnJB8Nsh6lx+LtNnLHpXX7iTRFCEiE2SIm8hhM96lUidH9EZ0oVyn1wbkf1a
QG+O5W59NLGCuroW0e+67SRNxsF1tZ01sfGGRF2AzuUkV+QB3xBz/UstkxNSNW2PHlVXEllRhH4T
9y6qwselQ3O0++w28buoDXe7ZzxXAiBs6OzTNmPSUGvirA2fiv7Auy5ath6VENUCkkV5CNLCSQMY
3h0ZAnGuYGjjLnl8Bhxq2CltqArOeEVBhyn0e8AnY+gT+B482wy3IbtTM9qBmAfdkvJuDTrE3Q0W
7KUC2ZFCXn0w1wP3InyZYIPgrCqsM4Pb+mDRmcYJXDYekgw+TD+DEa7sxzGqqTDkpZw6IYXtviDf
uxmPT57YxmeOtRhjT+FdCPLiRwW/HnX8Cch0I+/ZypVUZjQgvRs/wmoAKFncpmPtUIg7/7Uca/nY
TcBigeVWYsXkKCGTC+BY/yFvVHazavVf6VSiED/KunSw8PEe04px0MEhu2QSXbg5oaTcR7hsKyRu
kfqRlLcHFRsUXx1hE1u14qxhF9lRIqM8h6FrmN+BOv7PTawsEOCT4b6WVIc9PKH0/f6qSVNBaZva
N4O4kO8ToINQmOtqws9/j9NE9SIzqzvTIBnnOx7ai+IzyHGuuiyJJydBvQpT8+2iui14ek6ZS7TE
/3aKmS5+AEooV0mLop3+rdrHOqyHGMFbZp2BdECA3Fc39lA7u839PkrusxWuseWktAMTvPGN5ODi
7gOjgeePPyfcmwlV7d1iAMf0hP2WBcBAgbURMoA34eSRyF6P8XZPDdAtPh9q24tVJ7HktJkf0F7u
d3KeufCAOl/bB1z7zf+xuP+IXLffuf0BH1iHkGnRB39gLZQov5N4TKrQsVn/tkO6nAl8Gzeo6BGL
unODay7AnzoXN8ACatNXpNRBql0e7XRRblk81SH7gIg6oqej9o6AuL/NsynnHiElIPyipaoS8sdn
42yQlfp4a/mK1o974TANeffhHkm+dcD8XQ2dy626lqIrzkb8K3W7pycb9TAR6xXfrWOBJC97TBFI
1cfVAqWGPtPBPfn6yU9Ta8yYugZvilwbobzBBouLkWW4FwHc/Uolz7yjLf23+2fqpk+IDsZQ22xS
91Gqk0DIiNwWS5O55pzGpzudF+tjvVMc8LXBvyqx+8h5ylQIO2+wgdEV9j/rj7NWJbqctdIDxJ1S
n5b9b76pJSp7lAzv4JZCsAXmRfIzKgu3Y1dxan3IWpmFOVfsYBK7hNOojrrxU6h60fFepDGWBygm
Aoy86pARgedDiI8/jOUtYWFHi2HrCOSvNYfzPcGvpEe1AS4PJTEM3Blrw/rFniQqSEDx8CBoMGbk
26pH6gbQROZZ2CEOnboTCNdz6UWSTyXchMnBRFqqNeCotJ37N/MUz3aXL1p1ItOkYWamG9Rk02b1
iLQHT0pjCh+2KS8WkOtRWThYtyc0UqFmaKFyLnkTvHrpSd6SH0/K2Na5XuYbUWKvIZgdsy9jjaat
nE7Vw+3IsCrjA6GLZiQN4v9LuhzgSrnNyswOVSRrMtD3eAvWMB6F3zdtE7+mK+LIUUnpYyVEXvOM
BN5tRFPlKhRBWL4wy9VCApwKDU19ClS9a/MyzwxiXdCkkbGvdzFnnMlGXgJ1rJtTUQ1XD1M7eT9q
0NDVV4rObN8CHQoHgcAHJVDwcOCYcBqVRE8y/PUceBcopK+cY3H4sUCcTEzLmn1VNrCh1DrHxKNN
JQzsPVA+Sk6vVzilrQ+GnmbMyWBQF7qfIvald2gH1KHXPmpFo5+ArWZuKwQtGoZpvs4EdHXI4Bh6
SF4E2eWQ94qtDK/aPafhg35G6hBzMeapcgHf5D/ilJvWHbHh7kRJ00567YhSk0RqjiYYNTPLvgSc
HNFHR967OwGG7g1qFJjnwGVwvmVUZPolpdpQQv54JgnI9eWo2UxWu7x65/FUZXlytHhe3tYmgZun
iZwp1aY4wKjG7P9LP3LyPASZV+Pvh6PDNYESggb/PPML7VG7uDiDMKNFQs74w1CjLGI2a20KlKPi
3WTiYtFpQsU60etd0r7P/IGT3jN+Ray9qmac4QRCC25P9jOT613g8UWxx/DsUYcep04hizD1H0AV
YmETwrqmHkWzf5livPBMM3r3TUTGoStSjDWgCoNpE9q/iLdgk2nmwB6YYvzeSH3lTgQEsMYBN38a
q2byDuYcX0qHTdeV/YoFYgyUOXXuthKRIMNbIV+1qEDy5vhfWRzuHJEDS+DzB4K45Uuds6gEPlQI
jC7e0v5JnRolV7QZrcAVdGKAeEeO7cto6emeBeBeiayB6gqwP9PoWMFNNmNCA8YGwOR///MHtEUo
GCyTk3rDb1hugjvEUeIczOGpmduDaF57WsL/oqPdw5HPgjgUj+EqcWCh9sR2JJK7zv7QzZYnZPS3
OQnbbnC7SD/6dioFiSRAxEHrg9j66zNGaokjMPGw5D4rfGxgqfRU8knv75huPEmHI6BBnHuYZ7bU
9tzw4YigydcCfMN4+BPrmexGH7NjwV3/3llWGHT2R5Ey12MLAey3nEd9FRHtdfIBL+7lfdens/1R
drFVlrBwCDd3xp5FoldDYsphyMv+qufmQOcqrjxZuz6REw0ZVtXxexp5rLL4VO9jOzRoyiMLTf3d
yibQMd2Yc9t4cKwyvf1ju8yfGSjT+85Loz7E3twqlH8ALS18QGQVkOjxcrpiwMIsS5a1VJGAXMGc
eampHd8vy8m+CE9z2ukdczw3no1nKhuhlnbSRdT7FXx0cHgiBnb6XYTOGN1OU++t8xadEtHhn5B5
tA5Akg6wTXzVCOJxdZlRiHP2T8BYg8eybHWBS6jl6i1eitJX93ow3KHqfi+wf2CDxRnCqDdAdltE
M/BPs57JocGPdtJlsxRIBjmSKAOjD5T4e32dCZ2C/x2YJ0jdT18YGE/7vnnKP8rz6pssjateCEp0
/Rxyb9xxJ/d9kxgTknXjHh7AsaDATaTzcHiFNyv/YBocqjEZxJ6pS4DcuCKDz2Z05EtFq5GGuqS1
b01L+xWrYj6YzadjP7GLoj6ZW+UJ3C1jGiqbWGZMn90PiuVvWrtGAzZ0X2KgR5yayRROu0Y/QDeo
El14631yeAgkvd89mL6vNP9Fa5SIJX36P8x4gE57IK6zXfCmPk6qTGyA3j4GNs3jFQf7slL+TZC9
MSfq3fqe+6n/9YrIS8xn68FhnZDMbe/dMpUaMGKGkg9NBRsmoc5g9RlVObh8SM36to7QjxhOy0rh
FOAtRWAQhg4tmgQFAa0zcggwL171lFS3JdMFGJ4mfsIvrT9aTeuSzKBqnm9XEqq/zueRpWttmiD5
znkOhWdTk3PuWm6gl+q3KzCK35OuaxCDNFF7gPHv0ozMzrxq5xC1HOqRRfKV9FfSND8WtS9qoDcb
wyHO7selRE8/FVxCi+26e0qU45FjzuYTUWc1mu9gxvsWUY9YFzylZLxq/Pcyb2rVPFbQKyg6idH/
wY2b4UcITEC++kHwV9Qc+Va+mvEXhiAaAgAKkItycSPK/AQaIMDibWcYekyIQaPE11i8lW51+2zl
6zet8fzw5gRm+jrpVcP0lIkQqTJBUBqZyQvl8029io/IVl1CxDxN42VVCm+8QeiUFqWvwJ7BPPwX
J6VXxLSyFcvHycDmulo+xJJLGkG/F34ks9QnYjZW9qiUh0jp5X/wVX9WHN5cgcZSTBya+PKFuDxI
yfDg5RYOcqZAiYy+/AaQ08nQdFAJIZsmV1iiCIEgRDgEy7qqAJLbzOVAuQ6mSzCPqa+F3vs+qeDe
O07IYvFwo4b8Hk7YF45IbfJMj0Xg/vkT6gITf+bby4eZzgvxQtYDPrOabWWBC/qJaD0IAJvQYd//
c0qsn6xHNLTcJPWGhs5pBgVcruRZ9MHG7aV9fCjM1zOq/Yyvo9nMt1MJ45BEF74m7v8f6AGiykNS
csSQba4XGNetI3XW5nO82o+1g2/nMgdSAp4qcj5RCTsbMEd7kRny7Di6X4nw3eG5KyjkTuYgTqBu
NuilEis/VxZzR4JP16pT8x/8D3900TyfVfrRzliG6HdDZsRt9iG4ThluhcTMLvaSaVvBSJFo9GSW
lyZSiOAlj8oYv+/zfe78oo/rOaIpaFD/ldy5dPfwn0yZqUvD/mNMAAy18QP98K4rP87ho7NYrPrA
LO6of+fUofJ9BWDegjHYRlahWhldy/7jqhANm181x3+tCXst/EaenMylxJM139BTY/SyHc/YMBSt
QrH0v6dzLDDiNYHrbZGnldPK7QLKbkCs6Y+Fj7Y8vvVul7wOq91a/NUF2UMfFCks6JZnP5/kZkAd
jiZ9EMESzNkGAaGQM8aEmjvGMKb+RfqWjE/hzvazGW2HGWaZ2QrwwvTe7ll5HPYFqSD0ufjC8KDo
6poabq+2p6T88BYXMFh6u3zj7lnXl9a/99ihNxOfSAHBSLmuebhAYe+i5hrS8FoRjtvzFN483Sjr
WmKlLgk0pFA9pph3GwYEiBzv70KIwXavDO742EySJgff8bHE+vzTGdY8th53J7Rp+drubFdDwDBA
kzJ5+Go6jSN/02g3PVr7fNd1fKPOpYqF4dXRkSfTYAR+KILD6CqWPcEf58ejgEwSrqYF8sd/qWAG
WxBZmgY0ZwbXNBcbhO4sw8XHiYYD9xVQ6518MNuLYUwdQ1x5bKXy/GM6sQDsYXc5mBhs1GTOgjkP
q/4KzGOr19L27scpYfcy7+KJCt8Z9cchN5/obgCvcJTle4JzzJr1CeHxldWjRSCxQzFIN9vDDdsr
mEz7oWciRnn3NR2c22RZDsKWb0ODzO9ETryMrzN2nxBHLTjLdbXLmBYHCDFJgWXEp7TIgYGNFLyN
rC109AvkUB2aLBGFL/EI7W5mVbHGP5KYd+d1hgs+DbkEmf4V8IM8x5HMYR9Z5ppGataqrQDrBwx+
FiEGO5EATjJgfk3jwKh9mIN9EC2qzzk7A5p/9f7al9HMJsVkrLDgzxmNKa8IvsylY3SjwRqCERdU
OiatAAFngK0gdN5ibue0irJKPxfbW9yFKS3ED0TNKprZBQA8JmSOT5FZ6mRtIKpyZkths92ZHPBW
mgl0I8cxjowibbPg7niu4XD8VQOu7MHsst4V0VaoEgfih797xxRJuei2QlWRFri9DNg2WIT7+IOX
4/rXl1+Y2Ua0ucP69UQAV/YO6D1BM+cHWQXn5h28lvDSyXJcAMKHCjowvNb8iZq4mJ6AXqpeBbY/
3+A9yC9/amAyugA+DtlBr0MJg0EjevezWnktNnecw+5mATN7WRt2OUPwfdgRFRk9W8xwDuRQGpmA
2LX+7xJBH0A/XGXcm5FZkvP/NwUDNXd8idqtmeoElLtCDnj6YxyaWhyz2KZLvWywypRFsHEje8Qq
hJGa3PmQ/BLVdQYQICCoQM1nikhASYG+kMpS5vWSXHw7JHr3lFzRjM4CO5H8nrA6n60L3FuiSXUN
zHGb72+iRoXz2YLktkMQoRKLKVUkvGM+fMdwAlunIKIuEbRDuSiEdIop1ucQn0wYIovq2nAVv2O5
K9fzaWLL2pf39fsfQst5KGk+RbmjOsqweJ3vP4dynNV4Z7zIuyDcmhWy+2ISEz1onSM1CDtyVKU3
Cug/NBEqDOhL1cRsP5abtegW5vmYIFDzgy9ziu87faoyCdWJzD7OnIHtB/LzPVNu0su9ICW+h9nS
U+43yH5zLX4zLGz9uaWiORChlfPmYhubjP6QsVbco2Bm8S7qTWC7Ya4eVwcufzYlqi69vJ1W8bDh
e7PMWAuURys5Zo85RdXce8uqjdqMV8vk6oOcDDMijvvjYeRR2tqsu/ah4OqIC/MWcpNbNAMHWr1X
+OIf82PruK3dgzVr8BtQiNtLcowQbhQG2oaf0HUH3G0F8lHAjDZigdFmlIFByQWvPjcliMF9XdFP
/UT/iczQh85LdNGEpwL6A+qCAEO1HHuAQta0vHHeozS69nh+4qzqsI3VpDR+tQeUFzVgjw3o2q8C
XXFzw4OgQHyJHF0QlZwT4+2sof5EHnPDcDHs2htNiIiyyAX+2p5mNsR+GsoQ/1zOWCUzdMp1x0Xu
Y6X2hS4Wa9Ho7MlRFl0A51xBH+gfRPBT8dDhvujai9/6r8wg7+eyO8J8o5Aiy9lz7182Tboib9CI
r+Rh+FFRD9wnnMOXBFWqqYUZjwJJfF9TjVd6bvnBkfyBQjFdRoYO9LWpAFOVSbW7qmYTlSGRivys
6iScE9MfBI7yPcXlQ6SGMxjO12PKMamrtT/OoFKAgoHWpH3LDxXhZcvCazo71ek2QUTGiWjxBVwF
0QZAV55zRxVK2HSd1EbKV5HU907rWZKgV7byfSHY8f+QrwHgLaG1yqlgyK9k7olcb+bGRo/+Wd06
/PmnCgpLn4mA+KNAXWh/sttixR1gGtDJWFEdjBuG6iEGAMcHtv59NIL9/nPuojshPSEA6L+m+nMF
ZhXXOIyzC3DDphjSOczqzm5Od0A6YrjaGDJUylUH4bjoLzHPXe0D0GWlOm2NXQxJkIVe/4y2cLDw
QIApmjMsoQpGQT/ozcfBZEuaL9jHyPeUTTTAGREBnQCsX+JUHDBXsPwh1aIjdzX30fRUk6PCSKxp
Z/crk3tNnwZ0lOHcop9tLsum9e67tYWcFOx5VRYn4qAcUbPRys5HSBwhhHugQGybbeUZT8qc6T1t
yUdJkdXe5ddMQaAA6w9CfBJweksGAvCoYbEpZLVOI5fFYrRgM3QT/IP2ch7FIWRg4bRXQsQDmdOI
T2tY+D2i8IZWxlu+F0lm+D61KdBaSyurDX+QKtw5UOSsqadUj1p2S3IBWzU4SLnuZZUGY4paZHM1
nKzO8/fCzwT360QsMgQrFYW4LMPR8zh5ZeoY1JJpdCW9eRj5LzQC75TSkQwPelfo9E+qfzCmy6Ob
DQvD4HAelsfGpomMVsGGU7aHUaycpCqR/hEHK11hj3y+/1z9q1+AsAUFuxAuin3qMQEBQYDcT9uZ
p2dRPRQ/22t9bfOON8MW3JJ9HbZhGOi6r8shBpbfHID6u+cWe9KVyDbEYCF9/xr3cZWcAJNOmY7o
1aoSKB/7Aff/OPROA5DuM2nDQUPCKnq19bqncr2Uxwpj8JZvTI8+NVDrb3SATvUyt6E1BU/2ZkjL
BHui/dCHHICraSerl2MH/xALaVAVRMYeSfqrhCy3RN1w1DhYwuNKdu0I7kV0FVYeIoweYhKU9br1
seJaGcA1SODJD3IyMorRoIac+dwWLSfaLFuyGSCWHP4cGXIgoDmMmSKYVqwctH+1dNz1T0+/mj6+
KT50pDox96EHqo875WYZLwBurxoRIIGr9JmMn8zYWkCcSWZaGgbw5TGmUly/9CF6qn+yO8/q0H39
qxaG7k5M1vmA4KdwzsTkrdKDnTXhAFKZgAb8YG1UvXH8ghzPaZWzGQcS+qC1WaAXWuVdBJKMxLI4
mg4i4WkvvAPgpNtAYOt1WfmwGKM5kpFzFKXkim75aZeHV7pBJwHvH86/er7Vd7noTgzZ/9XG1Cqd
OJKzXfVno2NYohJADmyxi9LPrWXoP/90eOBNYnmkqJtWwPRBPEWNoxxikIDpj/neLtfxMRNbeDBt
WgK7OIUufV46dvV6U4+jisxVejQvzy5JM+N6YTapGfUW+NH1EZmh1YjfPzQVIuhLySNur0T24I7m
VMeHXdI6byjVpDmufrKIEXVqsKtJqZ1UjBYgJX7sFjOddr6mCvUq7nBqw5pcNFhY2acIDu1141kd
p3DPcSO3Kdr0+V/Ou0ytpE4zPIk+Nj5zQqM+w9kyxhktgeGJGgviOGRK35ja+HrxNlzMrER4R/wz
DkLBN9iZvbj6WhkQocdltIQAZ4Sic1nAm9dziYAOPbIDTNdSBon8SWII8nUlo9O2Scet9HnvrYvJ
l+z5yKk7SX7ASDN+YHPf0UJiJVjDlGuo7SSZhvABr7z4XcwY2QZYs8ZsEQxjPPAbMFQGWrMM6xhl
TL/DUbLOQGK4N+jtfQEsplmMVPsDSZKgDQ3P9SMqRC1dMpU8oZ+IOrFqOgSmqjO7N1bnRLJspj0u
lnLMEU/7Q5nX5Muxx0+yvjwKnuh0MnrTNv2kD5B2Du+/gUF9uXEYeR0iwa7npZEBvRswNPauOJ1B
wbCHgiy+9X7tFwuWraTjaVsOhAWDKiT4Ver3m4KhEu9S4KAb+sS4XPR+ukiQrpwnjbq1h6Yl/qD/
Hdjcmj7ecTD/MdqGORTq+h929K4L3Lu/HeWBeRJcIGZPxnU5FksZkr/1iPi3CMUyEk6q7RRqri0q
1TV0bOfAWcgzXyXu+hwm20LO+2ni++ueo/X92rsI5AJj/SFLxCYvCRiFKPbxi3YjVAOcQHKarBMj
Um0heKLUScXmDoovGnvi5qZxerNqxdNkxwQaTnS0tddimxNiD13sRz+/v0flxMX2SYxBAW4jBmBM
0b2l/iqJN9Ik7zb12KSYybPCTIhkbPgC2oE0NVHK0qe792zRgQScbvrorHx3MPlYQgPjKt3sJBg4
usZJ1nOR2zzrtKCXbJAaShHzZl9U7kVj5tJ7YOe2pYuY0cMAzCnL6ESzBmvo3BeOrWTP7/e5ULY2
NL9HBuYXtVgEnU3msYevS70c8bDLe1KL5nywvA1pUwmrWCr7EcfCl0Twkv9gnhpNIE6j89wHPm21
VGKRHrpig5BfEFuZAh5SLi/7YcGZ7VPnqQSPIpX1LaK8BAAOyjXBEbD8PHt9OWWlBbzDpOs4z9T6
8r11z8PepFu02IQiRYn0p2PL/bDejuTMhPvqxF9OcjL6ouTMzXRVCXgcl2nIY1jurI4ihNO9Nctz
/B3GBC1MwXCKI2RgFqxUvmBcglH5Cs18RQjaGqk1j+Ww3CbdMTPbPnQbOpR0/BoJnKKGZUr5Hq2B
G+fvT7VaCS+TIJPvBt7WvsRVtqO5qP+HwTR3EOMVzffuiA5DYmXSCVMTXbeLFBmISCIWEDn2W2Nv
JmEurmkylmAwK0YImrmHOjZcs16LW/A/gM+rsnZzZo7gl7gEwMOSTTVsu+mHB+kUKqBs9wsrG+SM
/h63Cf76DUm46SpaUsbE3Ua9obOROtXm7LA1F5dFxaFcdTFCgbu1ML2D8K9su0sEZZvCyjyRv7m5
+2OG09w7XY1p1RPIZq85LL52gEHLDtGPDMG0dFNdb1Gd8chwxxS6pac5jLGxR/sKWH31u5CTL4nv
c3DZj5V4rsTzA1m/mz9iflV4ZjGTSQSjtteWRabbAcISFl7HOhXx++JhdzRyW6BrClIwk1zKE5hU
czkKm4+8EelSrI9CM4O78/+IxHFae7Btwciu3fMUD8jMEvICZAty5p78s6SA86A/ZHWxFdD/Vbn0
qY+lP/4EDvKy8V2TDK/nemF/5HY2BTzMfiRhB3TmYxtFtx4z/mGQ9KgWrXzLuKYZ0u8k1OmSO4fI
Seae60H8ew3xiLV8CCIOoguMLkeFEnLcCUsYXgUi0fIKIpVcNsl3Ur5DlWVe1SqZbbfI/PrkUfTq
mer/zJbkF02BgmUt/lMaGYk1zKQweZLKMYbVG4u4DjlN7El+zKOzZqdhqI0zJ0/nD4l8gnXx5o0K
goiob/B6c3cWjAtXQJ8CMRI9YnwtFRu/rK5vJrXhBpiYeLvot7tjs6GSGwV78+445QB6zlsuLKke
uMd/E/z+IQjjVt4gwDdjlB9cEwQc4nZ2FBRDwmXNzuf4hZMW9g0TUvJ15/gWx/ieWedYoMslkc2X
27qiOgAWg4ZGGDxPLWG5fA0yAT5XT8bDJ8KMAWaQniebXFiwvfw2iCQZKg2PVMtLvCoqeI3m5U9K
49KRPlNxXRlwJP1RciErxAOIat1Y0nzzrEAoiL4RZIRTH60Y06/LJ3IpXlucdVsR8shBJp3S1rsw
B6hokEWjJXrUjQiztjtaoQ60H2PGWWh8m+QdRuTG+4DryxwtpptxkQ9xAxCETwUZeJxi9r6E7QgV
1J92+gJDV4Z9aDXVlbTTWIWx9x/A7S8FocQdjx4AcKuWgr3r0OA389dSFaHtVrTMFHtv7G6zg0gT
8XlLGtrWUCV58pit3jtPDUHvrQ0eAS4cUe0F4QBIYZMuKrGbE+TXlqv4NEyXu21kOAGnoGyYdP+u
9sOUS9ufvZy1cPGC0SUnk5CGu0XhsB9A1/W1SguPvLOaTa7k/Jo/Uy3PdRHWr4kDvYrvfyL6fJtA
2N4Bgp9MYjSjdqHvd6rWqHZzajBFYyGRRlSMI1hOmVeb1itReUKnuYmiVzyzLZ2SnEVBb8ZByzE5
ab7KyF5saCYhM+NLnXG0dZXyaLcEiX1M1pdy8hKn0EIz3w7+hfhf18AIniEmJ6oxtFXgJLk1uuo2
GGIkg9uFUzN4uhRaO/oYyUzjJ8JOwhLcf8Q9f81J3v8iO0JQemTI0flaNM4T33KeniqXSliWCDKK
OIC5KVDYHSR9uFcTCYtxF/soXztZm2NKPVPwUZWByDvKdUkIlmROO7ZBWBcVFQ3HRFKADXjj1K0l
lHrthIW/v4NEdRa4bK/+ttui6LOUXOleq+6R6nVWyFkwR/8QnBeB2Cy6BQwBRxvd647OuYoIC+Nm
yi1APw0MXimgat1USlOed6Lx7Mmiqn4Goz/mrduLQG2kVHIprLMuru1Hu67OHi7v03GjqTFuogi/
Oc+rrrRNKxdC92bdgKw5HEnHrDLthrGdVjBK5G7X6xZNdihmttaUw4GcREEjiSWbz+3Ou1F7ZfkQ
epaEIpq5n1y+IrA78fhzck3uo+b0wq7Yworu/1y8iUOXzNmsu+MRSeLsxqYkwXXQOtu6TkpOubH9
VTKMcA5ln94QYCr650o59FtvriqPBhi+aUpUiQFGp4Vd276efJyy6mH5tG5QF+XeJJ7b7bUn6pig
f9RichkU5E+l883oR3n0x3yvZVuCNGin8UEM4juw0eMP78YZNNriEJ5Ouf1SlC4CP3tcFg9lcF71
f67Q7Q3jySZV0U1l0F1LMaWa3t7ae8tFyklcteU+/r++nYE+mPuGDZEAnUsX3i7wQ+QtRwCcNcA0
Qrgl47JDjkn58mKpfKDYMJwHnkpkcTF37EH/ZfmIwPyA1uqL4SJ8rpVzDjRlA+GeR4+B4rqzstWu
z0/cKLJRNq7IsnId75i2zKuyfRcnciGkJkZtDNDMoYnbayRpgXgGb56GkUzAtW2PvovXPW5HUNg4
W+bmTHhNRR9P8rVQrE6cFgLDSiTy7KHujbdL0d1h1/2BBCNAm7lrxngOB1eZp8GW5EV2pbhp514P
YjvxZT+wZRzPRU24mw3JDj+McDmWO6zHcWUKXJDBB+T3f5TXzNckHsXo7E7ZbgMzZqSOsJG7qclw
jTZKmvclRfia5HEMCmOVsHyKTvfggoYBMtPXtVyRy/Fbw88H+qJCQAtSzLk9LnhU5Ar/bVDSFDPD
+M3vqpwnXwwPGrhwTCzGDuj4pcTkgS6u5DJAn//bLK4zl8oJNbHcoJ0lVVCqt3jLjCv61uOFSeN4
icTEVMDLgAIxKgxoORPpjjDETDC0RMLr5xt8P5srHxzo160lhaIqfVCRyz44gMQrnhxuOL6m+bp5
GEFbQxIdSG2voqDXLwxNojOCLLqH26ZBkrhMhi0nfZlYFxqhfhCe+vnk+uQFZjRlxFnbgV5doE2Y
Ba03KlcnA4ex4GU8l0o5XnCf/WDVcuJfWAEcy2HrjLjdrvJQWm7mCr4CKPXmviq6yAteqzfvD1E3
POuvLOTrtlLUPHHwrJGbzOd0f6UU9MuNnJyL19fP5lwSf+AfcMukgn3xzf79tt/rDaDm2sY8aVFk
WG+4bCU/bxpuAVKzu6rFMj3sXNwFwbkhrWmkHUtp/yMJ6Oy4QVkbMIb4GCty2OrKTE9H6K2dkhcr
XF6A8EaBZsaCHIQSsmjGDssMCFnBw9mSM7mCB1M7DASqdgSJlVYmvpQYU18vk1+Q9raoWw/zhL9a
xXs7kfvjLl1xCTxFJGkeMd8GVQ4UytObeY5Y78o5oU0lRIk/NHaFjvpOonSHd/JS2YWK8iAfKSX9
VbsPeKFBWmNXafHtwwYKhB67znz6Qyyf3JwaAG4aPQHo6FXZElPiznH+MI6+84Bdr10zO3K8DplD
j34XA6ZlW70XC/8I0asH/gmN+cvaRctd+ND0uD5muTJE7oHMcdUHstv5jq1c929rdUQ7xTOXr7BS
uXn5uzaAGoYer4N0atqyM8+85mNW5y2OcYe3HduYLofZz+oN50b7dlHdLptNIIEspTtquQlBOnOU
aVo4PaYleW0uUUPzwBBmjGMDcW5fLKu1XIZQZ6Oy9lLGUzUMR9CeXMVGMD3nhytaTbn/ZsvGrw6N
oi6/0TdGDytvIOzY3/dg0qVaKVVlW38JS3y7WOTISn4wF4vIdISap/362sjIVRqcFQEZZC86IrY9
lNSugQE/dhLx+anJ2i8UPQT1Os1P6+PJocaYCtg2vgENEBo5NFP4SDtoYnQQCRHHvPBWg7crjtFF
XSMgRsuN6VIXZkl3Js1d6cYqPif5eE5YWXPzwLJxZ0jAAkTK8UdyzH1s+gO34gwPyU7Up8l8Lms0
c0glVtYhuKxEniQk3iGup/PizwEsPUjePRjtRBDmdbSNW58eaKDMvuMruC/UR7apN9jBG8kaADvI
jxD2NTP5+RR4iPztlVgv+WqLjAl3aWCpMMebmlkEIJuztwAKdCE/RKJ1RpC79Pjdfuno3mGJxrAF
tbAIKPzYgL3M19FheJIzYWPUkUwaFQIwV3tT8OMEdfkf+ywQCvQpoH8zNPSy+fLDqzw94iRJ5ErO
3HtKsrWQO2dMeO5tFODTY5NuvqU+5jTX2P3Fj276c6WYUkY4w+RUFZOQ5PkstnxLYaAwyIIWc3ZK
LLb7m9SRIWwKwHJWqsrEV4i7GWutT/q8A+bpo2yETgjOmDz+UY/IhNA1t1hVhfgPZofxdKbdoghX
lcFpT4wMQsyCuHQ6tm9mWbNwiDjPWx18Xj9k4+LrYJBKVkI0MxSRABnLfOPDvRRl+gLVrJqSIcaG
bKD8ppHPy9W3c8KZ/UtCCKM/PADKWIea8zDhs2rcbTYDUZhpRp3eGce02C2dYYG/zlhMbVqkgiyG
NIXL/rZANM3XClZ4JAEZpZt/57ufnHMv+3kNL6f/5q4Pt8ILCuZhvHb6U4d2scqqRS658LbNNjj/
mUxOBO07gz7ZCpBDWi47d9egWxudaWzcCf4zHxSRKLsN+ULXVQDeXHRzqmnGojlfB4Dz2XV6GboH
7qXJkxpN5fVQ0AnN+PfhrcR98pbZaMGJC2iHHu1bCf6JahAXGFgo1xRYmAwNYIO6JM41yjZQfsEd
tpEqx4I1wHl0ddEjYsmznjgkVBOBndy+qjr7hgMGzDMrT+RkLz0CPDh19cGwdS/qZONAHh8UXEY+
8rP9HTDHt5I3bLnFXFkhGIJ64rnVMp0ncgz5kG1tp9VVVbuzsA4okPCLizHxPFOG7cbcSXOKEBZT
FpUD5IzjTcNjzHE+yOIew4G0jzAkUAl28ZJ0Z/zzOFC5uMiFAbMh/8aVi9KyvkFnXDNObFpe+Wz/
8dewnF2qa2uD7S3sjyRZ/0SxhWbHuR4HYX6iac9DM94WgJ1cSofN67iaWsygWsDVhFCIsZJ5VA/N
XohQXmI6fmGeOTozihAoWFAyy1D8eEoquUWf4mWZ2LQm7Y4uUcs9DyDKCjbhxAfs8b7MV++9T59g
KPsdXCdHNG1b4EHZw7rxnnTsjoqhSkNo7yAAWWHc81xgzBKSDSIzReJw3SdkpGe/Jad3smgALVZl
nkkP5Pe1aAWPBsjIIeEdDZ3rO5hnSGUWgQL1MSiJjwjRqxJXWEhu93QWnilV3a4oplSPELMBL/F0
Yqdfxh05K9CcDe8f6yQQlTCLzlboxEETettUI6wGZYk5eZ08afvqiiULllO/+brGu2+x2C+eYkn5
HQOf8fxDiRgmJlQZ+pN8EfQJmsV7l+escISF8krqF0GaednSZIFv9eX6U4oW8xccxmOVPjj5cSWF
WbHgrngKx7UNMGn4hZJD80r1huSVHYvuybwlMTKwNpWh8XoreBPnjggAbkg/A52kUEOXRCwWnXYG
0G3TgFYe5HrdyphRz2LfJmqA5PM+XkCbmwEUKT7WeEZrKa62Mr2mmVTTRZjQ91FM7GTDC5EYtRp2
5wozckU1TtZ3ffhmouEDfApjk/sph/+rm/Tsnu/WMEW0hi8GELx1qejxIPqYuNiq1ZfGMLug7/xQ
FEbZ5yI2jbDZlWeLiHIdLOsl/g2vYkoFq8T3m7U+qkJkb0GrJa3o1HAr8l6v6+Xv1Iy371wx+AVA
7FYJb0CUkqtz+t3IOGojx3/6751gRWg3eOHMXApiI9pHCiVrzlI4pNumda1XvmSeN//nAdKW3FVA
Pc7tvMEzHcx0gk+kIX1FKVWztClDcwz52VYWo7TwbVq8arh2ovlbAr3wGuOUw1ZKDB46sh5rkoFe
/7XMFgHLyx7EHC5Aac9fP/OgzHG5Z4B7DDBLazvV2JRC4moyCfR6Z77CnnQ9PJMhQH7FvleP5WqA
hlC6zuSgqoZHdRYNXGIkFq6NcSUnNUoyCthbtbYrxajojvFntNGtPtMI/iEQc3a/zR+G0FqKXH92
3nb4GZMD1aP5966m/ZddARvLOgp9CGdEHc8oKJFuZmv32689Jn9L0P0ydHIXlqGYoZTFRBaxx16c
SsEu+jxUWF3SKPqSk201jyvcWEPeeQmtkS9AKP2uJY+JtCR1J/JVKQtLmj5Ky1XFM77jPctDdexH
t+tlk5h83Sf8RKcoQUlHl1fY69EKikpeeBFwqIhUctPGmzKuXM2ahomVEOq+Qdal0/n+JBhgXiwL
cSOgPQgWxGQR+dw2bDNZs99ndhp8RW2oPcLbncCT8zFTTu6X8+SXGgeOxeMJ4TvT0mta5lrifsUl
6/YOGMfjsrQUCWqHArYcxMHTdg45Ns7ef1jDMAHxCMgKQ3Ihox2FCKsYZpf5oErLcAifJ5ajM8Cn
sNQwGPZmJgbXv04rW3IsJQ8a3RvElURwtJ5YY6aRHL24tE1Il3cEmtP0sAKjNE5WyMKsYsk7c7to
WxSpCojb0IbSROJyGyzL+c4QJWwx2b6orIqdRDk0GWpssPOs0Lyldk21MCas6Fidm2h6jrLvWpzO
rsDxZywz8aLVD0CX5W2ErheZLVzaYjYShQS2XlCIUoMZxEMEAu2/6LM+ikMBIxNX1oUfRbO1qQZ8
jvDNk+rYrFFKG5B0FDx/eubuByBI8vDF53Up7guDncCrrEsSVr4QCxCz588t4h2jATMvVRwnumSo
ZDz0CBXUsC/IRNWG622RUAkFjuEy9Su6rZNhbXFjNsYiYTpEDd1xjV2wX5cMYWK6B4JAl2Jo1VZ8
trlC2LhZHCiW/v/7M28FIoakE9WcVp60YXWIMCrBe42Hv/Zdg9gZ5zHLk51rkqd6rNOEE0UnB3Nr
AIQzp+lk06FARgKkGWA4Y/gw0Io0Mt3ROaU6vWhcK+PM7lGmLrRM4n89Vr7AwhTWJX/GERc1w6Z6
JGL8Vby3FSWinr2KF5ealeklu2cubqbzO3/5Q0WRzoXRsq3IaLwBuolt9OGwe1uEGLLl1LiinHW8
yQ8B0FOJ7gnYyJy8emsuiuU8Yt8CEsvuYK0CFVwkOttX2/+7wGAUrFOcCy9SBVewaRFA89R4s1UW
dUeAvupTU8mQjXyLq+T4zBEXZ0mEMlQI+LkXo+yJ2hSxlMsqhgUkADmQgLnQoYRB0CKWcob6LP8K
EUAoEN8mkN7JvmaCSW+3adO/6W6TZmskZ1BUMjh18ojmvGrmr4yl0fJirFg5Xy6m1PF0gQBIkkap
nfIcNWdBevXG8Bgi1PpjjX2wEwNv2D6KJzJr/XWLJ0YfGddeIOiFnPMX89lJXfxTb9Zxyab7m4gv
os2vCLLbBJ3AGgUkYHzrMNAH7jekINbOG4J+nXCc95h5zekBQPChScurnzrVvZ+p4t8ebQe2rmLD
nhtfQp2sxxrE7UI2F96D4QUzWYXrmaZ8GYW1pXp6zYRzESPQX353ImfULWZkVE3mEoy8NEIT4p0P
cDhhUoD3Xik8wOPKfDDUA0iGVuhhd/AU64TACWLKv6ADi5bKvDGVYJIAU8xxDfN2cTmsMIuKjjzw
WhzcBKRjoUeXF8ODwMyT9JJ162hXoe3e/nE/BeLLXKOafjoqL1woqoJRSAbeXpaKGcpWbKIviU2k
4sgKoAyWN9EmBflm8C2S+6rU6k+WGShR/gjw8MmZ1F2xP2R7arBbp++4/c7y2BimXty2JsDPe1aC
qfTEtImt5bie2bqJXSoOVwraj7dX4TDD7G7LAH4o1D6NS80TML0sW7R11jB4zHaXUUWbk+gW17QY
na4yXjgrus2dCDZ5y6uh3eFwiH6JCz0ai+rQsyjxNZV4unln+nbwDaUSc8z0jqxXm6HHgsGKT3DU
WrkUj8vQk3ssrMFzpb25whLzFG8CHLeaXjJiOppMfo2o5Fn0tVgg4nr8TsONBjn2qVFrSauuHenD
pbXUkWrxkrb/N3qnK9/5xKrfKJ9D3+3/2ZRWMZ7xk+5YTMGYZvED2SQ1piqD7q+HNrwkoYNsxxhk
rQ8j7KjCp4eFDluYMz9sEkw75tgDtCoCUuOcjyx9XJ0qCwCdnYL+wTJ5H+YH1pQUGmXt2WHscKD1
+C+NhikfCn7pJb5oYpUKAgMWArG7DWNKI426H14akbeAit3v9V8b0czEAb9jZ19Odp6crDTycgw/
ApPkf7axCILXpjBc7WZu8NLeZgpV2cvQG4TF6zrSwSVMUhU9wHDr3kwHquaoGNiI+ICbsEVLGsn+
oSShaB/fgjCAvyl9ISnTr5FaMQOGiYwsdLT8lxNiWf+sNggftMZK9f5tKYTreyCfcBtkVxTQ5i1Z
oXt0jDy8cB0Jxao3vqknXA9ut2KFF6vbVkcp8RsENeKGpbHhMrTGSNA84G+eiBiWufI+jar5Ubtg
ErUTrAYeNAGPQNxNfph/koxwp2uK5mktPhdKBmAPbXZmEmEaA9vu+rMqYPXXLIVfLXHyUuW+z8Ul
4T6xEyVYXYhuvqI8fMbMbQ85EGev8m243OwjiCdYkmPeTlnV5pljllxU5ZA8kN3mX6bsqaJszYqo
KjMDn3MQN2nTaiRGQEcGbpz4YPGpSt0BUaXoDlA3VQbM+2i4xjn7oE3y5hruUhTF3iKXk8mJZv+l
MtDdCcNHO5e03AqY/B5ibmXMhm0hK6N+6aG3XC/Yzl8Ti+kufi6sZU/m9AvuLNZuGb4oYaXZ6KB0
9NBkhNYuT+h2cIHqrvEMc55evU9ZpKTyqeD91QVmy8c7B1nqEGUp+YC18BzdEXkmWwIIiSsakeVP
8lJXId0VIGMSFq3258gKi8C2nX8ZZ/BxosLtHCxngtl3/NYwwtZrxZGqPIULS3PEUTH1spBxfnkc
RVghHgBDToZMVTUBHpdWwow+A0B4MhEVpkDU6hUvIMHgE2gsFR+/5hMkLDxXDCKAHkF5g2muEQiz
UnW/wna5EtxrfNTsHeVH4dOfvwUomAfBCjt0jyTBr77Baj2G0wlPM/JOKfpT373OL5xK9GJ4UuzX
bf1QJCThvTxrJ0zpYV4TlNKYBR1DPLqgBnbwxiaPmrZAcLBrwu/0UpxTr5KQ3iOSxbQJmDVbCa5E
lqD3hv2UEnIx0Vs/afaPamm6tpgKbnLYWsvxKUKfY9qLwGGyocDUjV1gn07WjMUE6Tt8RczOuMRm
R4BUP1+drGFqbSwwdNuTiL5GKfU6igvI3zyf1IrDcsx1MI29KkCmOcem6My5xiazUCn1n/3DIRxa
qgC4VrYwCUyfnp5oacPPWAtpYE0Y42XxABlIWp9g2g5D7DC6NBI7YcNC59XPEwCzEafcWXIbAG6O
LWbn6fseKOfKN/h0goZySPEPJ7vWsMtCiS8jUQXPA1u6IWakaMx7g8f+2f4pj73xrHYuyj8wTNNi
X9OV7oiMD+No2PlKxjlt1mpoxlF3YOaqV9UF7iURTFbv09iLWV82huZTO7NvO4Eh/7+zCflvsWsO
BSwyjGtlRlv3Laf1YNz6+UqKgz0hoSNo1POlLcWX6VzqUsponKEQNtaaPDszXcEg/DoN6nlJP4PF
gb8DVtobNfUn6HNP2+lX8a7Fdq/nT2gKoa6GnJJXYcEIeCmEtbSTeX8trfFerhsW/TrmaNRnAbwa
OyZmgK05cVOKOFj5dJOLW6AO1W7OHInAjRFxBSKJwDZgh1iitK1QJTqDhTbL4LxUzsT1h5779v8G
hMYev0GDPjhSphWlJFp+5sePCMCZ55g/xjC60UxEL+V98x8xveA7E5fH8VcEPtoofcVqjTQXnlfO
NtEYdXJuCK7LkwVd6qfZIZb/+py4QpTLjSLsmqUv3awkuUpn0dXILAS3hTkAA3kbEHa75H9XLP6R
YGKFifWlq77VrQm08WxkfbVfY5Y0L88nfKoVn0HX+q7UdHowfO7daWS7a+3ZUmqK98PrXd1pJzst
TZq0iaLHDn85z9CDFF55Dqe7rNyxdhPoYfzCEJ/GyrVwsDcRkzP19w5F+hpEw/bDInBcr4nopjrn
xzXJAGwypYZs/x5KltbAkiAwyhwIKddWufMCzMRaL1WFpQJ5/RRp+8S/c968YoBrBqZVwYM4qqPd
NzRLA/nVNFc/aiybL7K6nH0dmZ8+GEhUWPXrw4m3vj0aB3655zLS4VktS+BYZ9eQPuiVm8t0L9Rw
sHowibzzhCNX4K1o66yk8H21lsSsvR5L3l2lo4xaow9MfCKG0SnZdZ6qBy2T9JnmjakHkYQ+jNHx
XXsfMpA/Gxxq9ytS/u1TAeqRMKDdYgRZhqxljm82dFf4NW4htI7ddnUAU5ZUzFwdDn4lzXqkyuYd
rbTZsDOjXEA92Gd5SYoSIWxp/jzZIEr7FHWp4OSA5X7QjscUYSog9hJlRwiP3fB/zpgocNfoG4LU
hpzm3GCaIsEcdYq815LPtcKPUqIdYEcBoBh1/WzRxLZV/KU5y4Q+dJSmbP6cEJhBiI5kEJvVv9Ne
y0XrUG4rPN5sY9pjzY30FVt73QVB9aqNFSQrcD9t7+kjRcObFk2g7UiyLRPz27Db+bYwYFN75Xeq
bVc1fC12XnuWRevrmGfrFKZZYKSCfXTDx0rxaB+xUplsRFHLeguqjA7yyH0WyZaqREaZUtA7ufFJ
8pL9AoM2zJ1NTniL/Y686hxsQy02MseLgttXbV7zvqcTziHJehFJ+msi0tzs+vyve1fVyuobdw9Z
ZCSsz6MyWG1sjcHd4FNaqVrvx9Bm8WDmPMrk2Q+hsBWSzKoQS1NNf3VaRhUYkbLaKZH7G/u32+2L
1GYwYw7mC407/QgBUQlyfNhxMZV+dRyLc6kTLOikc2Rbk0jzvZOKE/MvRsIHlLFr0G25/8JygS7f
EsOka6SBwbOJCdbz111e1ybEluDo7dSXSk1U2wiiQeX6Frg2vLH9p9MdVdDy3c0CPIwzKWSxfOiu
7STBN/0v1of/OhmR4mvaztFPWryscljUt96yEQpweL1VDZ3hMbiaQudmhbh8Ngh0mEBVjCjRF6zc
2OWvKgsE1wTSaODVxY92m3fAHNUxcIiKrBQLntftkBh/eM1F124NFZb/D7B3DovmERMR2f2bRY84
gP11JoN8Fl8n4AUdxQXBZsUND6zphrje5fPNgvbeUhWLaG5RL/Geg0XLNXZ/Q1qAPLwYjBeG5Osu
qd3XEYehHCtrY66rdGQa+50lrbz/m7NvoX10dFnlbTKdW7w54r6gWgLUQGYauuVx1Wf9OQOjiOx3
geryNded/G7OZUGwN+n4IfluFwK/Lv5YYOVwFZyxSBpXb4JI/grYzg2IKgSVNF29aWeok4COppM2
fDyvtANjGW24E2nR7gugVT6NhdrsJdVA76KA32EHb/6DS50pDWg2YKlD7yKc8FKMPnTjPHLUyIOQ
uBwHu2hXHGYMaL3gwyqKSmTSmmraH9FKoJ4wN52+4xcd/CPXSDCkUFz/jS6uJydyW1EWt5HuixCx
0vJY/Uhljv++Tro5wNEfE9VmkgB+c3P4xIgOUSFXuGyKVokiuaC/bErjR1XHYo5lk1TQZqrEXjwk
YqfNw8y5cePl69MNijVBExtw5fO9gNibYK9DGdGI14vfVzup4VQ7Q0gBNuaEapwb/LQ0vQU1OaRs
M2F7jLZkVJq5iPWGMKk4SEImG6Bh1H7tkUwn18s58jQ+3IUBTQIvY8OTjeaWtgYpC+7f9eO/9E3c
JWHALT5SqQ4ZjIJbFvH4ELuyxms7XtDVcNt90Gwv6ctUfQ90mq3gukJH699qA4K0lZovn6GId+VR
cp87YOcvEtvm+c+6Cj1lvaHCTYeiRpwwPVZ/NnnvvbUNMX4fqaUnWe8r+HTacqqHDeS/Gkbj8YaY
nmtNVRUWFBdMqYn6yFrvAJjJyGuN7dz0o0vr+8CW3j20FATeMe7KC4hKGu3xbw4jZ38HrYywBFf9
I2KCYw991qQ/mcaATSM7bDEcPM+G+AoPMfWkTfJeU7EK9pVqUdPtCAc1gKokHH2VV4nQ892d+NcA
150LIBcGo9HQTZZLt0uV70q1ta1EyiM/CQiuK5xrNUkVBODHtbXYBlRonM+bOsWaFywrH5pbRGP3
510IYdn6A0gKPJ2286SNX/YVCHmFvw+zkn5KLO41ArjAXYnXPkmsEyQZqN7P402lB9m3PglOKmsH
w/xGz929Wz7ZHHQ8CVaqrFFG02f9t7sywDlyBi6aA+3/ggBit8qamJBJ6zVkIf4MfxmVKkKTRH8P
XKg4EQ0t/Jsuu9HUjJUrb6gBPPb8iTMZkaHWuOY9Rifx2hl6SK1gScMJu8PW/meBuInNNdHD6z1P
2O2HFZKuUmSswYqKNToP/TEZttkyVev+gW/nCzT49RDTk8TO4eNezIL72OkDppVlmEOK9i+sAMPi
aeu1qlzSnJivr82JMlsujItQ44TESirow0ax1XmZSySD2VCksdlA66gdK8XZabmiKVEkvKKvf/r7
JayRDaXXRzj/pjhspKNskz5GOUc/F7Rl3DtOrT5hKG5pOpgzT69H06xAqnEoYkTjPjs+fvBHLWfg
rDaSpgn2JGPyIKT6FHGnF3/4EN4LlxLysxczUhGykzxc6gLEpBZozB0Mp25F3Bfgrd41JX4al48U
XZG6vLnW/9/uMKiyncQcNw0wg/kO6obBwTE3NTmo0YGd1krGQISk6wAhBJRDoaUUY9tZHacDWqpx
+FpTUw0ndK8/hBskRpsETd5/ZCk6YNfZ9x2qhfl15gA97cn2kNc1P6okHEhM7JrdB48ObauRNseY
kUnR8QnwzZQR3on2StDOc8SHBkkxUTRc+hHvFvbkQWd7eJRUNtn6mtRVhZgAHP5UfAed/3W5/SIB
KwkJ/l3rirS//UygUGdbY0IZC1YFOz0Rw14ji8Cm8Q2sJ7vGGD3LpuCg2OXXBFP11mH3dzDirlbK
BO0jh493Iu6FUm4cV0OD3fB+LvpIa94gS5k8rCouRqNs8XOdVVauF0tFhKEsg+SnMP0ByGTVSzLy
9imXqOkITNUlf1u7I3YqgnPHhMuaSFrUeGVmQo3Bdasy0c1Sgu90PGu+Um7mwfyi1QJgil0/W7OR
XmIXu7AFvYbTdVvEV1m2UE6FWkaj4MYQ/UKjqujW0oBk3It/JEN4pXTwtv7Xjz8THsW+a6Nf9As/
pEGLEdJ7Jp4Pgqg3+B1xhE4YnZR/rsVr9yiaoTAH27yRuJuOvII4rLPSlBfeD4OcIwRMYIp2kxk9
xv4r3FNROio3HSo+igfz5LvHNgexQd9ug76uu4onNSCSwKogIPbZOHkdNXwlHlRjz8iLS9dJLp7f
pACEZxazx2SDZ2EzKeazaa1CQxOslhGyMljWPG+8ZfypSUyCHsdaKNg2oM1yR9lPiDH94aJbSHlE
jxj8aoXOIYTdce1vf9aNWqW/WvKqharppvasUtSd25yOI4uMbiaRP7nAtQz7fXqc9Xi1f4X4ZlVm
TAWrIc3bRrSdCBR/NkCoqVjLErmJo7nKSQM4QZR1eWvjbaKLgehIuLS5GIT3jhjRGebFiPBD40do
AiVMZTOxrAOVCsuEOuPK3jNGmqE80nGHV7jmPwG51lSpld47aYTHwl5bhX1OwDbKhqv8CjI+sOzK
6kKrFlnzsaYh8cMJw4mFQUwf01AIq/C/TB7gkW5kPJCbAE4bID2Hsau/Z0FTk+Wub3L8EdzjTogO
WtOTMb0TUTx+yvCf6r2x/36rgY/jHI1CgeGvgvSzyyKKNoW20PNT+xWB2ZEOoBnbyV7XfYI/ruLH
mw2CTdM+6iJXdE0weWUPdXgfAKYZJC79mqndbAcx4UFbfbQgcAiRREZ3qCCV1c4NA8ziwaFeBeUE
XF6uAqLSFx6ZhFA/poGXSpLarlht7UQxufgwlhngrJJMPFfl35HqU+UTFQ60LLwSVExG4xuRMA/q
uZWf2SRgW3dzOX+TzwGhWj2CgYHE5eoEgvcpOxynVzlOLsoX6ks7a/imvy4OScmtsGuxOrNvHW8t
MiXak51VU3cbsZJTU7C35w88HwsGuTXBsaNsDcNYsJxnAjzrGl5E1y2gUzL7ies6rE04cx66DcX4
EoLewyfK5jwfKzocmkBEiYjZVQeUUNRDmShukCiHmP//2EUKxO5tIJqxrvSvnP4s5kPy1MjsrqCr
BZugZT47CVcvQ8/m4yShXYghmZsnFtuq60mz4aaZgvD3PYn1cRMip7+g1vq81JvNdAjYRnRUJZU5
VxvIx1R9FvJpG9la2F4pFgI/h1RuTjXw9M11BgB3t0PSBMcZvi3CHjN2aY82Y/ORg/wQsUomLyBb
GuPyekLuhE2xLlBDn2iyN/2KcVzA9d+OPwpjs4xbVaBlr4V0bY6lihGacBY7PrhLkwbO6BZovULx
z1wxDUb8tSQ1qyV0sVaK7LkYPd8l0knfq7+oE7nGCOagNkbaVSlDAxngYbgG0yOhWNLOxoKV2s7n
n9xZxB83e6nWOO5c0GIaCwvAKX5ReoMTQlb+/C39k/EMPxc756NX7DkymuiwimnXRHip2g7ZHbsJ
2sygRdNWXnACaeFn/ov0ebRI2sioFolbBmRZMD55olEGpnlRxe2Ow+0VcusMwhCwNQ2ETIp59aKI
3mUe3pjvj19T3fVoRSerYyZNxdq4LRaxgtbJQU3J5ve1grRhWhf3gJoc3NNVl6X6wf0VgycCFv3N
fHn666KQC7BAhJfqU0oW55gOjVzd0PG5bh35DVoSiaBOK55y3WvbUYqGJBgAeF4tlL5MXe9KZfZo
H13Ty74/Artgx8kbMlregNlxtrncauYJOtgoQVey5NO3vBjCi6KHSvy/gdKx1Nhs5CAdUGF0qxX/
caLnMuT6LwVrwObBSz8XGbyvVsdO3tlRKoirC+u3gN3Ln1dqYk13K8IPklPrth91x0vw+MsfEV59
45zptT7YhRJtjiX3MecTM7waWdNzDGcDSM4L58zjXpeKdWNyHOqUMCmocOmnzcgHf/ZVubvXCQrW
3qgZohaQ9/6iO06tQnAK3e/hwehqHzz0KkP2hjOFStOrEil/BzLi6kWbMgRfuJSXr8mVuT8oR3Xv
V0uDrs8rmnm0AyzjVFXo7kTlW0dqToq+73tDbGaTUGN2BtzKYVUCOFd3R7UGbQCbM5R8SkXtdnlj
waof1AI0vZxhNIM6hKVG3HgkCnnSTNdjaasUX9cQ4QQ6NBPWvJosd3/lzqM1ekt/Re4PMzj04USq
xYzzaJEOj9FywX6K7CZeknVTGg0TiNadECBPDL6UCBjXcGgAig+o7K91ksL5aJi6mHFlltmwjgBo
NJuysz8mPWBRD6ZEmxkrKw6KSA3kU2rug3c5k6Z8sIouw/rIdXELpEWs4tamm+XUttb8y1UJzy3g
85jM9zMiCiWQCi9Rrly5rdmz6XlGAoRiLt55/PepcQYsO74pJR36Tz29lJ9IEls22KK60vu5xTcn
5w4a+gNntwZPatC+LL41/iICcgxNi0mbimsWFN1AMhTJpOHnh7xDCtpAx0MaJxFlv7GDfMOknx0r
2S3qwRx2HyWXCCfJTmuEaKQLME5wCQj7KDaoAsbohSG5zGcQQkIhupV0FEqvqcQaYhek1HIhlsaO
l6OxFhSxcIpv1qNdKICA35z7yRHzgCR5ndZYrpwxZ6oBdar8R91a9X5uR85kBvfHqHEAiVgHDRYB
tB6AbmSozP+aui473L+lZEdg7+9CZSYnFtAc/PLoZsVd5sqjliNpbN+ciRYVoyAlAsFeUY67jw/5
a/Cz173P2YhkB4WJCAd+ZTXyMfNLh4pTrO9SclE7PkFXjIuqJgyIY/ue9Pa4rMGCuE9Td5pGe/z7
1mZ0QrwqzhoL35gWTdENg/OdzQTiwTvRye/wfiK3iYvv/ao4NcX+JafnxxGleo5gOHJF1kTpzbbo
TCzp0ncYNjhtHXDIywSJEBPf2AJCowtSFdDzKvvX7FXJ8lpjp8pd8hj69sEJMuqcXHN6998PiQM5
3yultG/FuThlb1R6BZZkt8L8E45u4VIq7a124SR+dSUwgziGezD5bM2bsLO4A6ZhWSFZ+VRO1jkc
zefp0IX55jviQkYoKE5jEmT17h600s/cGMBJcQZHbK2cAoWkhzxIJCecsJWO5a9FjPvmg+ZfqdXW
F4A8jXE7peodAj1pJ1glZ7pCDQ61U3Y/AZdSMID1BgzlhUwZNgDhSgYnrbPuTkkKeigyugxapYgH
Gnlee7RBsYJdBwqAP7ZtlM28dL8md+addYIdSoqmCGnTCnyka1O3wHDkHGhBimOkGmc7JrleT07B
I4bA3We3oKJxGnM8rkne/XsdvX1LsR9mj3ca4qtp09BovilWTDAmuGcLNcX1WCwAF6qBBhXkl7O/
bamwgh2vCsMkHvGx1p01LS2oFkhuXj+V++MfYXZpF7mOz7RIcA8oWEBHhaqjunQa+bpNbA5H4dje
47mvDnG1U8JJlJLOrFN2TSDpU3gbXppB1vYB++N57+AvnMz/ntsteq1aFdL2mwsUTdjT4HUXnwLL
AcTGu9/X0ddceewvVjHbEJ9ZyFPOhKK2jKMAlY9A0B/zefl1EBszP10T8WnrtHqcrMWACP7kGvdI
s1d4pQXT904TsRHrGktCza0DOSEIiRkr7ZhLXo+09WMyE0xl2yk2eLQgiYXRN5G1ObiGIyuDB1Z2
G7m2QHoVj4vd3OLyWOkFhusY7Y46If8OrYDQausOQjVZ8mIOOIEdkjBifPjIHvYV6fZY1XertgPr
lKCzswB0ukyxnfsAR1ceQX/3TLl+on17Tkvc31XJ3fTA4xjSt05yM2DDF+3Lb9o7Y6HsQjT85gEg
TEAD+g4d3Ss1rSDbnJRxryto5OQGMFOh2S3vzAR8K8PrgPjUIIu23tJNtZbYbhfzIp5D1HqYpx+b
seb2t+GeI94PDrOxjbv7+D5ICtJ32MzTJPMu85Oi9WIEHiqYckc2B6ASBYwJmlzaExLFPLY7eBOh
vh22gNDV657YAfOk7tSUQaz/bQehMQag35iauO3H3VC+ingP75Jiek3ytSZ96Ry1yz6JzATpVBhy
9PvVn2hTshmuCFisRYK25ibNBsagajVSdkO9Okd2oqfxLIQV7clG79XhWWmcAW+dI1oayoX2dHsW
cLKUoPDTwUbNPKMBFv4t8moQZqu7cmL4+xSJ8Kz5zIsNjBtx8EtESMojIK3po2TeEvawlrToobvn
5BXJ3oEBwZ2yUNZdCPFDXJ0hAbpeoKed6SAAdzIFEGEKnk3A+PRrvmC3afxEjtKbl/FIrEjdTtlJ
dBCedTMJuRLkoRBZVhCTv2a9M+gjZLqMiWra68Zo1yQosbnEX3bEVoEyPXsd6XLGR0UZut+esNLt
Jh/7NyJzP+nlcPAVk6H0E26l+qvf+j16grinM62nBAQbRpHMAsvGjE2OB5xSlKHBi/n+RrLw+/1a
h+3kfhFiaOiRgT91HE6/24OZoq8ibeBQLlQ88fK6VmupsTApeYiBDEJyTw0reOQogrrjwsaijpku
2FIskdhr8P/IUYKtbmfn7NeTIkIy6Fc8otkU6SNmZfWhmKkwhJOyCY+SfwmwdB9Q4AsURkA5Jl4I
nQgoj2SQwkOZ8lAENOqz3+A+f1ndgRuneImid4cVMNb36ay1IUJAQIWEdj7Ah3r4L5vZmM3nCTMJ
Tumk5eDMnVfJZUZa+rHB1MLLnl6xqcfTfzUfRIY3ffCS2nBA0YfLb51DOYYsNdK9RQ5/CNLtt8sA
6z4rb0s5Hz8Ph/T1X1nlJid+x1znk1ezhdZPg7YYUMoKtYtI6q0f/ytbQyfGHup9N7xBsoiSbvRH
SLnuVhs1Ex1+CXGog8WdnF4yPeXR3wmk17ryPh69pI6TaDva6+utK9IF3XnehVJD7i4mzOQn3TQk
aCt0CKru4XMIgBzN5L0lUAb3nPODJrgiV/wzZTo1DQ4I14Kls1tbLY1LW30vWk4iiWqIALhhSn2N
KqXVL7wCivxaPxYWwHc0zaRsVQedomS2BImjqNeJzkdFfkXX7xKTEX7CcDSJ0lYczzO2JTcI3rN3
5DTL9uM6wOg0v+/Olr83grBDwM4tQ8W1wyEzeXewhOv/QE8BRd2oeF5Q3+4EwOqgTsNgdCXfkFHc
hIdG6b3QaaYFvu7iw2OI9BaMSfb1a0Kg729+7/sg08OcL9pyrUVU+J0q5lX4grfvFPrURRuCznQG
Ip2bRwh+8Xu6Ey86qf0w8ptMLjqBvlG9NAEFQmIVqNfsMX/jUc4WEDU99uoqy19bQ8KXIv+qDlHM
cT7vPVEu4LiYnm1nVrXGc4hgPW3pjwgWIUQlxnvgWzF9n3FjXtu0Nh0vHmVMFH3zKbvbEOdizQLx
HzyEzmA+WzFLnduIJiyBKKvMn23gduhkobj6ixtoDDR0ga+U7DbBZVE4WUGqSkaLSgYHjfAtjSUo
x+3xq335d0qeE1lHT3ifAQ9UvAd6fr14OSAxnz5lS19XxSg07CP6iaD1e6f8jd0FCy80TtHeqvwA
7yriJVPGtOE+ctaUsbEpaYFYRV44Fl5UizbAEyIr3eSAMKJNpE/rccsqWpmAJq3DzAPxwwt7FP80
DfsmU/091xbyPYIa7puTMhY8BXfMZTEkDE5dT3j27CHlmQw5T6lQfWNVqbjioAzMySKz8rS2p6tr
Adh+yyIdb600edhyqcHAbA2KFidHaD5jLb+FIDHILPgRET49scSgmtZNyXOUX8u/cjAs8WhMC3An
FB/6vWgjYlnvm//89t5d+Fj3mRCSTJzH6OlEbLTUfPxCjL9A5Ai8pyAcGbBPRIdh2DVrdEajIrn9
fwwvTPJWZg8KsabpuukzPJai6tpht27zdu2X2QIhcYEN8AYO/jYhPHj9aSImDhdf3wqfXZ7tOagb
Cnsw/G/hivuB3YVdXdlrKbsrLCA7Ftz1N+n/VOSoGH3PVygOSU817b/4E+qVzikTn1p25EyTBh8h
3+mtzxhLxbx7zowkRGkzehvZW8VkPyCMqe+iNEqYs6X9L71zbgH6bcUds2pTov8alI11CpPyACZv
wAeSIsyQCQfogBwmGCb8taxEJ01NsNHylNovINCjOOdlx4pWpkDx9wWntbzHm/emDjZUtGA84BEl
P/GvXsO38GdjA+cNMeUsxl8shtVqNUyvoX1lZLP/e1N8Rn7y2pzQhDhvI68JlBmMqz/aWNXplE8Y
23VDpcA1FHiHOWS0YSKqyVWnq8kCqGMQIEez9Z0M4dtzh7StnRztYz25eKu9mXGmUgg0Y6Z7b87N
zWeDwbKMKM6qtARvUxcXzRS+7WdjpfjmtE0P3xtrSTLq0vdy8JP6ofT0wcdL04eI4swltYTmGdo3
ekv7Jf/wqq+t9+sP3UKDRj3bxmmkVqacjtfN1eUp/dWxZPgFpVee/2t/XXFMOqZOjk2cCsdxixV+
HaSIraA3s8mlKkYH5iGKYD9mxCtlaFesUjoXcHoITsD1zGhC0LDfEOfYFcG3LmSc8pk1Og971ccm
xFqpa4Vt34ryc4E2dsfzOQDH3MetSueqe4MShUUUt0IP3jobeYCJ8bZ5EHh/qDKytR5VHXVqDums
pYIEaiEHT2yQaMT9a5hF6YJP12qqWnsD28zejaKykplOKM9zu0sMozId46ngE2aWKmXjNNY58vFr
sV4hArzxGwNCQ4C9d4dM6323/Jh3jQ8ZIt/zVO7R0/kn4tgObT4WwfyDV9LBWf9IrQIb34S6LyMl
ALY4Mu5WlXNMBzcNpVhBktPAMYCLFQbC2PF4hM0T5hWST0Reh8YXL1YBRApmdfVvh3V5iKCL85NK
fP0Yyx7TV5tzlPsfJEyZfO/Z5s2dBmxJgot9h7P2XX04CF8Ze/Tim2Q58y3aep7+OCMtaq32MraH
GWawYcPc6/VfQ1kdnYUpXWk5qXwRnzpmpEL21MKZYkedkjT9I5ok2FdSEvmY2Bywecpaipmgefof
J8vlMMgF2l7qoZkoab8iaQOG3feknU5+8KjZP76d26C6gxX6jWs8HKcf/FcVp5tfw6Po0HKm7KIH
uNKiiTAtz4T1MI8RDqrH3db6SoJeDLM3SO1d3Wrz1XGqrWbKoa7NqUi1aftUDu3nIf9uqzArOYx9
varkk2JCniNQsRJJoZCStFU0/HvApR/E68FBblTO8zumflv5LtkCroEUqBSyL+vRyelVc9qaO1Bf
Bh4/MhzI6QlN/2rrDdAc8kARyh/Re44H62cJ755buu/TSYot6BMrglV0GpPCVLeGu0e5eU2cT4tC
G9OZMbIk4clXBzWnDe20VQfXWpccegUw56/JRMpfRe/KU6Q4oU1u3uCFGaIrQAIOXORe6y6JeRRq
YulLZk8ZmJ+udp6z5Ue6qO77Ij1YGxQk+8216Qgnu1ameLZa3eL8kq8F2FTSGDiNZlWa92kocNK6
m/xmLSRryoFsjKOY1WkE1LNNWGnwMNaiawdksiLS0rm6rLoa8UQlgZ9WtIrhox0CX3mKj7YUKdXu
2RXBLngC3vCo1bBRYfVj/9Xf4zAysriihLFuQ+EyyIUOvvbEKJARGGNZ38xcm9vCJ/naP2X4kMT9
wMHc/psrsT+CIfYneI7Ik9byrUcdPqAzy0md1zQgHgzO+b+ek4tgKYQhKtinhkemrggu5zJbNV2F
1ibQwVzel2j22v6Et+7MDt4htSwAdt34ClwGSg11NYvKHCx2iRGwuwzraB5bnvpLV4tqpQwmJiPc
cl/fmUlG8DOeH7OHiRenjPicz/S4aRs4nz40ce3a8O+TNAlWzHM1ootW+HfUcVk8H5zW3tOrsfVg
F+uogcd2E5FQTuQHG9ARWFD3pmlsVLEVbBqvKHFvW7xW82I69yymOF7+sBMYNumX3fncr48B4jgG
Y1eATAYsa14zNEqExeE+MwzrTyjq0dMLLJ7Gch9gz06my0qzipOEfcRkrt6uF69FADqsxOxi0j1c
4lcWt6urbmigZQZP9u9A9dcs/qmJfxNJbThJBETJQ/l1N8Ozq00u7Ysr1Z6ty7hzdVKntAXFTy6l
q2wS2PhPkXEDirmLFBZe5waiHQfUdWdTtgMjdr9qxHAYkT7sU9ZTbuIjwTiYj2E90m+p8VifNOFp
S/wz2ZaivMDXafqqL9wVuShOzgzuwGrI+oLokYfwEacp6/5nZ3rQdZI8fbDdh3Bk9gVbS5RLLF+t
wztUQ5Hb8yvKOeoK9ySpWWlA0zj/rYCFZRTzr7zjrPAqta1+7tQxiG5a7FDwj+DJ1YiSHSMvu/Kz
xp7ZX1o/gyGrKy/tee1zdsloVG1yC2vP8gSG6kUfn9OPKdbIsT6rpKUEK6IVX8W/mtzkINjbG2Ul
BKwiy8/lzcyNf3AhRujxD0SXfisW9xj0z441uxe9LeyEBlDcDtdSSA5+AkztReFMNTfoY0uvp0bg
SZ/1VYOtVCkzar/6stLWVFoOPcFLO566Vb6S2V4H7Ag+zxVlBVeKKQkh5uoAYZTjh4W9vw/eBMlg
IdAM0hIv1SSr16rlj4HB74MQwf8AFbg/YL4SYwoid5G+eUyDs/aCdLfuvxzWfZvqaFA9wW5qQ7Ap
5am4GX/piGSfS0VLVDcx16AjcAF3bu1gls22Y3ALXUWtxai6WxfI28pYMjqxlcLPpyS6hEYbX9ti
mB4g3BjwTdd9MwP1gldT7tGgLe7f6PjKNy8wGrhF/aQjsuEiD7wCKifLFvQU7Eb0VKOWfiMtiHWg
c9UCxMz5mH10xiLEY/urxhdsTOiCx1o+CL0e9eSd6ueBPBii6eE1wPzI14BjCbk8a4rcMBCXPHla
iyZ1ybQYJziCP1KKQKM2M44HUD0CSjV7s3rCcge5rHMoiH5bLZXZETe8BWtOmA3SnLRBgWcTtYJz
+mXz/tqZwgLgFC8KqJ2blzqAe/XJyGQbH1SK5P7B4fHTzBVmGyE4A58KSfdNL0hsWvzq7qyk9J58
2QHItMXrhwbSpRL2cn0E1fEgwCYMUISyXK4jXMCQi+ibniGM6i8mS8amDLMO2kjp2a6wLf4TJbW2
Md8fes8V1z/6r4OyOkzOCm18XJzbzcRsQSL5R1Pkp1ckvvB87WFRy1z3KJNSeLfrTjydXlW0GGRf
OY0mHcTa/vTm5j0Ll1BI6Xt9PM1Lx+IqBCoMHyieC44fiOdZNvlcauh//fbPAdDcPGdJKbS1PN5L
cIBAeOcAghiyD+2ngeUyTBmkuSzesJJmzvL9Nd1oE/EE6BCkSyDlcOyZR3JtXk6QqZBmayAYw3ip
nc9t+0pKIfGUQ6lnyaW2XUlWtsYi5GM8ZiRKwM5s4rrdDhuIzrzCTXc5oCbVVqkuNHjwcUz4Pql2
Wh7QQTXZ7znTI++A5BR9cqyNvs5Lw7x/RWd7wHYp2UhYJZXtBQKK+ZD7Txsjsgw4Da5Dqw4yKqd1
wvozmXMmwTBkz090CD6FDe6IUkNt+sB4OLac2O/shqBVYMzbr40h7w9z6u0WPPdiqeJrE/QdwFNv
+be+Ads10fRrq3nQyr/i9K6voslQVGvSQeJMXwgdlqiKkt0v2FpB7FmmyQ9ghOZYdAspfowzcF1B
ekW+IRSPC6or4YyMYjhb/uLb5T4XfgcIPVYYPlIn0uNn8P1qqcYcy1sCHxYGOu50OJbhlPax1KPp
xGQSDER9VX0i5D9lprc2mApjNN4crc90Q3g2mOR2yimV/y52lsKhncu3x5PPuBuP2Gm7RVEzo0dn
LlL0jlhUQjJ4J55GAAbOgzbFhoCEKFGHa82XoAJJ5ByT+y4+nqhwgp+9yJJ88wNgDPqFuqIezgmJ
nTmbP2i4Sm4fy/v5JuL3njAveif+o8yhFJZ2/6Xpq5Z0Fl5GUifYO+z+YVofOPxs6nDU3GHRgrkG
NuNpkT0OKQ76zCLLkCy8EiYdwj8oRLR7O5JWJNjPRp1VrnQbw3rGUiOEA0vP56yfn+2pxVxx2z/v
t4r49dIbokK5wau1uwKuzOfaEBptBR/bUmW/cWB1t1Q6kdiSDFTW27hdLNjQWyliAt3BV55IeSEz
xwZJNn+62yuPSvE/4P+JY8atJ3fyCgN6VRe7nzCvwBW4FQ3+fRd4q9UeLyKBq3e/lw9vTH33dlkC
gv8a3SBMLq1xqceGJp/6vpIGwP4nbbPq45mangowSocHGHIPH+z0Yamt1NOsA9Rpq065dxdNM0AL
5gKg3wDXEX/UYH509JPf9g5uk2o5XwcRMRnt8BwCcwQsevb7L/G/oXhezqIyusB4vKXHlP/uJk71
/Wh8ALotW8BazXRlrm6gw+0Ifq4OcTzWOzUvQ54aRFn/6K2ok7Kxnuz5oDjlVpfJCiFFo4FF2Pzn
BdNhgSrXdGi2lN2CekDLc9D3qWGdf7rognW+1SYcWejWx8pXFZK4tQSEx793HuGvM+hKtESnqiLW
abQjSGKFdPiWzjas7y1cK91LRxZcxI7LSbKhUGjh1EQM/DjAd4Dw3WAPCKyxVsmvTFzvZcJ+BSnX
IrYABqEGFe2WItH3Dm7rsg5LKbjrHbrebxvHsKuiD5SafGHWYBb+d0SETDBbeph0OQxHdzrQDVuU
fj6x6XcyPGqIg30Bp8viR22pl4pMTnfF/kUedbaQVkFFgNRVTWv3AwTs6qTXNV452dExtDJWdG32
aSD891df5FEjt/IkrTJmTgl+HBFkl6Rq3q11LtatQeJ5eTRsjD1DOco+kpXEXfjEOSeyJBecrtdC
QFom55KHqKpfaiwH+wTFxnM6q4hyHwWDS7aqpKrCL74iXgeI33FHWySIiBqJcgk0KLwJR2YfchcX
Cp1aPyb5dbWLIxNmWtw9lpliceYzqSRe2wdKGT/IZtXBv8v+6yIz2vu9Ziazt0TED3EZ1kQfe5Ps
AOiMzemlP92CNUmA96AjqGXQYjbhurKPuof3vKLYQh97j13LUyFdQVzpN+SpULTEVSX9cMLcr7f3
RCVfhpaGQYspu2xny11RvZC4rm61q2YMFII/NRQFN9Mi4cnxycPlBHZnHYTs3rJc+vIIORPSqgF5
fazscVqECkyPTZ8LcMUCOVo6XFTlntX5U8+VFLSWTbnWbCJJHCZytEjJIC1oW1K15gFP8P1QcoZQ
ww9Zrv5wAGqT7wgVA94J8tVlq97gnqPrwBrn49Ea5JjnDbniHtMOXCYvsA06EOWaxRV0vKUCbz2y
2YufJWK7St73pgOTKAtOmI00mD95ILuJILPavka4FjeOpenR+Z8AI3eMDj+aEdY7tDUdAuPWeE2Q
LJrX6ma2cJ4ziEW8H7U4Y8hcmnloKrDhuReM/9usPkRMlyrCQ2Y4Rveavi8vriyZ8CJDmgxDHg8X
eoY5VW/mz24ItdKFlV5Rfkm1G8z1x1a7HFDj0ZCBBXr5Q5uww/y0bJIqcuHYG/gCM971VVhnZIJl
Tjmt7iOQnff7fwYtLSC9DQNc8vh6KDzpC0vXnsexFBbcd2vukoOUVmFUfJOxtIfhj3RdrAWeje3K
tarhJWCCGx+R38GzTyxpqNdsynm4adgAw0uSr7B9ALb6V7j+XAvgRg0Q1P6bzhWNJfiCzMPLM67g
z3ZAiwgWWuFYJ7SbY6OY27vsJUgOCoXZeYnUKsZmKJ0zF+o3LE7vQlpOGwUaH03OL1z5Ah4SqqzT
U4usLF0mOtkigrxBFQTkLXKjVCte5L/8b+Bvw5WTiARumvFlbCmZ/pADF5Wk7AQ8ta/oN9JfePHb
guTK1QfKcS69ulb9uCEt7BNCFE0VBPaFI3kxdZuVErJUk0+NVtf0m0Q/X2BXb5mshIu2cweYzGsB
553ahQXNTgSFH0fKtzE2ef/k+G4x8Vjq70SzWuSwN7pJeT9ICNGTQrI3DVn1ZgSYbYDSCw5YbLJu
adIKB1kxvhuPaK/Bi+xUZVNqFCMwbAKO/dvJNUvXZITHfEWPmBN2ytd8McEgK1ZSzGXtZKNX/qz9
l9B6h4p4aQXDsqa15tnT4CfSLHvlMviDbJ6Noej2LpCs2xQfz3/meaEcFKnoXwHPQ7uM1Orc71I5
i0E4qO9ItoLT/1fDkwGuzC9uUzV5a8lH0oxjrpnwiDxR+uygUqBdeCbj088/U3R3t2l4Jf7IesJt
tnHhPmvguPAwHaBZeeWHhciRMD5FQm7LnzIpziP/HGUDVB4NBAK9JoT+eccsP13PZkWLg6lV67AF
rxPSlLq6UvXA8ghmfTTe0HJQH0GvfEhIINQ+5Vrsw04DRFQUiNcZXkyBavJH/LW4/SqW1GoZZfrY
WbqE9+k4565zhU6JBWi0RagsePXfz7vm55oC1Zz4iJ1of7ivva2s7T+UYXDLgxB8Mvmx9XARNYpc
YBF2v0MozVT5MTSF9Xi5tDgMlxmLnjGIsBVwfifaGYLaocg3JnES0weRO/Gwap5Bwk8YTjB4c3nt
MJ5ymzY2/y9Hs6mFKVbJIPja59rr/hJ9ZHopcfrdwmevCWfA4hGxH1e0F4kIehvLGcRejEs7adqd
G+ih+yVZB0yqHkOG9QTdvSJbmcT7dAbKwauCKGD4mhuj2UdYLYZdskRrSiMVqLTeAox1Z+AZ9aSE
8lxVqezDoEvoQ8zdds8OrJ74FpBZRxmq88xWeFig20fpOnh7NVZtCvrf5ut2dBaCUF1ww3bjJD1+
MY6meDALxlDC+gZ7M2IIjbe+CuMMmkFVuA3VKRgvwL8fTYLIoXWQRIRSS8w3irpyCtxvf/RDg0FR
Hs+JtXoEE3/Wivr4vBWqVhtJpuvhDHTbAbznjLrTNyMSJhQqgF3E1FmofU7xw34uqkFbPAzAbJ0w
I6vH2L0wxVdf9goeS8FqJ4TrfDmhrPb6gz9NR+0gr9bLTDVuLIFkVzUDlSUUJQ5qLTAwTs+jW4H8
2pTY5VuSUR0qwkvVky9NdQ8XGygLsz0CNmc7eYxJwHtFWxd8qpvplivJjug3PqpDIZW8KqDGPWYP
BAVLeKNR6qBUnVHZvmkcWIx0yKDhYtpUr4eztPjqR4HI/UdjjsxXIAuNZuMtTA0Gr/tp0NczCpgv
btfKOvCGHzrsPRq7nQSjMZpSQiQXGU0J/8fMeg0Y7purSjh3m3084UNlK3YNdS63T4xwVE+4IRZe
TTQf/5qhm3bfgWcQ0pMmJ65dKEP2Bt/nhZC2Uo+byQVZvzNuPhSMWkdfHB4b7+7WrOmoWhsx381Z
XVG28QDfWrRHBnFg+HZX5WwZNtqPH5/RSqCMUEOCv6IwBKEg9bTsQGH+O+Q+MqjuTWIO3y9ngRVh
UGk1dJZkeXRBcg/Nl+m8a6MUZEOvKhNhO7qq1x1nvi7/MH5b3kqDZiIml/7sW1CRC6s352Ws9tkI
Rm5z2Auu+S4pko1/1g3QGGkAzIa/rPg8Ib0hn9tMyMH7IlYlmqmMOdnwwJvThfqQzDihjoJTUNo3
RroF+zXF83wMw18t5bKzQXnRfGyhB2wnwqrGFQ4XfOoB45qhL79QwC8DwgaodoamefGSzpcrMfus
GUGaYkguGQC+CwNLZIBhz1RMIX94fmv4xcFW6watYxXDgOhsxEozKw5103EpHcaJKQHA3RBFDTuQ
WCpjB6eTSHVf2Jbzbfnfjg+RQv6rJgtbhqlCpHoulkFXOz+94v3wHFPTKlZn4E7L7NZMOCNbxgdn
CUT5f97kkY02rYh+xQ3q9Ar0mPYqlL5ud9eCVRZzMADGXkxQMw4DrqOhUdB1a2sQ+NAbgtptmULx
XyAhEydbizfNBA77kKQlFD7lFfXl68pfFuZJThVvgm8ybD2Gb04PHDJcstzcraDOHp5cppoPPoEH
JBJLOklfvyxupKTdsGJn0WqslfNNiIm0QSXer4V5Bk6nW53NSXWbLe6yb7evBJnhMwNrLpoCAoRM
sF7Arhhzqv7mUhG52YDgm+VEExlSbQnPVGs4upMfPbX3UDejI26zFzP3POsRMu0WX5jMQcQT4ArF
eUbCKp+SlH9p9lKqwyqZzJepL62BJJOOA5PSN2vUsInwuyefk84zNwHKUar/bz6e1p/QvFGKl2EK
fnG+b0klvEm5OIhCP4gZgo8CO4MnE/QKJfvzg18T8N0ycNdNiXae+af4nfaxpvc+/Ym5ri5K9erN
7N8Gao8+8LchBYQG1T+U36SfymXNILMBfqFYfNOOYscuZ/BdaID6UXgItw+3ycKgsmED3oo+JJEr
omdpvjlvAIhOr0+/hq1tRDz6+yGVplPtuENK6DyH0HEOAuddr5ONwNkU1re540naGMCmdO+UHQr4
FolUVv8ohsMp5z6DStr5xMexuGlwW76u2TIj/sQO9Cowin5UpVFab4Iblk3vn9pBM3zhPHwd5EJK
cPHhMim+29JwXYeYzdIFMCDuQ+AfzrKRqTYsfUkSOyCpQAP6xXL4oU4NitAGcHCS/j8jkwowjzjt
VuGcWZ/M+y2b2RwYi10FdC9y4kYoEp/yyn0we5yjLsNeUXqrkS2VRzM3zH5oawfZfEMZx0TWsTQB
jNSTtXp17AfgbfupCgkz+PJ1pR+kU1Whg+pOiWfwNtKFBaahg+W24IIj5T/v7JYsVBLA5LuRcRB1
oaKyRF35sr4dGFd/B7bnOe/RgtgpuOOVqf6WoaDX3gbezor4pwalj/lUcNvmBJjw5gNlSj21VYuK
Wtmcw7nRZzYwxAvhqhRPXfa65J06Sr5b5pRlbjxdcFRTz6OlOBYpt+09a09rlffsEEZTkVgouaR7
rY1mocoZuvHMOje1RMLBiFjLN+zRPriVet51CXtOEOSXjNRkEOdcKwMmAMUtcAEj285u2kD0SnPB
PmZ7kYA41TLucqZwbZfxMLzQY4MN/AUA0W8fnqVZxlhNlaSYcKZiYmvYi8CFQZ6cVMS6ihmc7icZ
RaGLuLysOfk8BaDErLU4Ve6AAegN3hDjKu8K/SsCwnpROSkTT26Cc2J5JNmHb7DQOv52Ua94NDzm
DgiKpQCV3Jv9Jl90+usBGzD7QWZ6/KgWdNxQ/XY+p0MhmnpnI60pmzrvE6nsmmqlRY9+ircEukeR
IOPG+WJHw3LB4UzG+/wLRcmcYEB2d9VxOX76HeJRLr4iBqvsyRk72NhIAfIRehKWeQRw0a2vsumw
xnQXcEsN1ryRU6YMhXPACELaW6rRBbavnmlu8svpLoAInKqj/TASPkrvtX3R2f45Q3ADOGmtZX5k
GbNwDf4hx/Rx9a4LzXukwCD/6/0e7ZS7raFvme6IzTQT+E7NJiS1RFLDS8+o9MUvKKBMROsjeOnX
P0n5AZnnjuN7QWMik3rr7MQx7xBk0FY7d1wgPgt4r+UCpP1eDNlSxTPM9epuGZ15Q5Ksh/ViaGbS
GaxbWNgbUo4HWr9mWAK/73MzMSknEJqxpGkhOmJKY0LdZgM7pWQOMTA5rjdh6EAt9RioALG90MKh
4eTJBHYNyZyBTJ6OBYTa73UEkaG5ADynfIOS0fUkln3sjAYMtpbpwd05y9EjVc9kLgoB1o5XICG3
VHtCgeDRboIg3COxIIL2p0yuqmas1l91DC2PM963ya9BfmaiP//SFe7K75Y453rXo3sj73cWo4Rc
HHRH3Xp4J7k01d6TOneWQTYMB6UsmbW9wHVoIpsvvtpizEUtTo12YakowXxB8ZANNiLFlfgWMopV
T0kj8YRJ5gWdzeJfA/NYgTPxxqI66Ce2LiYqz1TzCS75s+l3BH0o34Wjo3CfiArOM0TXIpTJIj+I
Op2Jqpfw9EGyeRtxFlznIgXg/oIBZh7bgKFu5A2UgCv0GJmAgk5zRnc+HNr13b4GHSrHkxYYrIKp
lWIJ52vgA+mITC+gsxtANzQN3tojGfzygxeOMOzLzOOHiGBIGIetTp/J9t5fDXuBThviJKDbxV0u
tytop+hRkIQXEcls7ZZG7FPg2QSItipwxJATQbk4n2WD0N9Twi3MHBbVAMkYNSTYUmyTiBZ1Xpzs
r6wruL+eN2i+v2SiqY5zrWJ8i2k0nvhJ9KqCoyzuBvM6kBzUeCqhqS/qmvrPGja76n+lcTspVqW2
tmCze2WXUvOKTw4k3BLRrwEx170k/D0XlIcYfmuMrRysD3jB+49LXUGaNY7/q13tcoH04Czlk0tM
Ecq9Cz48aaDNnPGjv6xzsHCwBZGpiz3rY7n0yX4s/FWANen0Bf0kM9j6lQ37oadWHphPilutUt9A
AjYnF7d6MHBc/qLp+yA2G+/kgefoFYrksBOUefs4KfQdgtDWIcOtAhJb9t4S5DEOCV8iZTVPUXRd
UjlpkLd3gY5p+X1NQlVtbByOtVI6/qx03vl0tMVevKb4YhnLZPDjPhoudbSsWaHxdhOVJgspCzmL
4Sm5P32ir8Z4FZHE89bnHFir9vT39rk4FAmWLKna+WKJu1FCg01/qP1hWdp2t+U5LWHgHh220/sL
xVoV+WEK9St2b68XqvLh5Uwn6TIrGKRdfpicxt83xyIEH2Tk/JBUemMmMkgyWzdkOTi1ctvvHtii
EcLTD7SYYTUITVY56Yw8SirToNddsMahiXN6Oc0F0NRjJhpkb25csF30QbOEVVvn1LOom6JyN1V2
Egi0zny1ewoQiujVwe0Dvm/uEL/XSUdJcreB62igCWYn2x45HT0x1oXwvAdWUVAzqK0Ui/qX3KkH
sgzn0axfez5wbAX9alpH9p5rohgMH4HUkLMYyoKymEcOxzcdPeqam5723Md8igqXeNvytOJGH2OW
dhLg55W6R2X3ymO0fKpF1HAHLB4SJ4KKdi7tA+LOxsN/gblJxV32gQa2SoPcFAJ0/mJEwrE90JUc
g+A44pICfSTD5WNRjGzbYdicHZb8k7zxoCAIA36dXa/mjB+7cHU89S5Ky0sQ5UCCR1ewWpavBZuP
hIJf9xILhat23K4o3pLx1tkkNZY9D72cbIfD97DTadsDEfRES5XmQ+q2064wsM3RmbCJN5Hm4M/U
qexszg+vpduWs1A51UT5naOstGDyqQh08Jq7phcW2lM0NnaF+D+VPaZVv0gMajxPu1YTxb7ZjQFW
w+cJgC8VIbQzsM0J976noe07xmeTXNMI/INPnpvAIiat2N/HxQhiZx3EyQj7WW9F6vtu0O+3SuBb
LfyIEelaaogWLyyv2bPGOLGmBnAlZfLUkyrTeiKnI4jw+saxo0qYg0kdmh0kkfspBaOEB4dFQhza
l+IRFZnwoVgF4Wj8CK2AVF+3QW8qDxaAH0LqS1xjWniniZC47I9mGfPuNoOj9JKZt58AMZ0iVlzD
cPUmK70+6lRG9zkagB3ufMpNckgLWZDCI5acjy9NJDa1aStt2YuEUQLBkVjjZ71iDSr0mCAQEGJl
3UxbWGZoG+Y1xDzgGwGAmW4S7yxcMgXb0OTWvC7NgKHOCiiMyDO8LWQ2aBfrNhAXwbpprtupEhry
AqqspMCK9Z2UbHDvQpM+QL6uUThwkm/k/fz8efZewtNjm9n8iFU9+u8DgoCLcfocZMm9IOAL8TgR
mLQvRcevM4/tkktV1guNzBeIUjUt3jTFpAYF3M6BsWAadQy2hfBCgT69lzkWUiVDJUtr43s4KhYV
uaoSl7XIyVgNMIG8lZGy/VaU6AmCoYpC2wJiFNVABpnfdWwc08hxN3QWLMgrafHm8MsS8PGpFffe
QsaImY1HaQHqwtflOsDswG6/jf6vxpLq7wL9JD+6AqIbBFjHMv+4dmSVHWDYYwN3XzaQ8IH3lVDc
U8q3xQPEbvvubNZL1Mkt6NMj9eMw0rx8iFuDKkwywQL2edo6seze7LfNXoj2XCYOIIORyd4N5ZE3
i3BX1v7TSlhxiePB+EJ82rhswN6KrtuYvf6TFAG0L2VK6drBfM93vtNlcnIFPS4Z0LcK4ycUdzBT
TsIAM3ssRVWK7N5pUclBTz6Q+vVR6GYrWPEiriQzigHPjFrwZwEWbFKgAx2OK6fn/d71z+2GxpNC
9UK2COCxQwo17X3PRTowOffkSJemoky0RPkejSzeqkAO0nleZOYduLnDJOk1Nu+rNOkc+MdI6Rqt
gfyt++dMm8J0R0br33QVTNGuPxtHUCOIWrKMKktNRTlsaW4GhtJw9qQVqkau0BUIw0DbLocKz6TC
dO1G+ULgv43guvipSxEDrSokwynQ1AqYPG45GOg9X7WzwXVTWd5wGUfkle0AIA9Knhu13av671CD
U+iI+PDgfPaANoi7fu/eZkPXL/J4S6Y1ZuH0zVmsAWCW42XWwHyq7hRUUy0iexAW1GCf6+RnYkzX
0w4/4uEwAjjj08y62bZ27kXL8gCga9N2hS4tglkhD9aZ4xNoHjovpgIqMytvG7VNwl2YBGl5ChX2
s7LpWpiXN7UWCjbws6WxdG5oujGeJxeBl6dvUhnQj8Wbd7QJNovI9/YNYcZZ2x8re1c8KKl/0LIB
+5gk3KOG86VXYRQA3EdvhvDQvNGKV/Jb1bQQoyFcRThI96Tu9eEVJpXL9nkOxKWLmcLncfwJUJ+l
eUvYZ0g880p/5l0k4fOtnQFenWAgonXHsm89SANUre0R/g5fOZN3KAsvqv/wZhyMLgandKohesiS
kNTwLTc9jWtcVPJSH9QkDz3XmChv8YTWX8OCFKwUKhqV2s40xqXLmQX3uy5ascnZVnDnqizxdUfU
FZEJbCwpkdAJleuN6HgJR2JsHUsuhVfteXWrQwY41ImhMUKP/9wRDMsmy+PvrAV0akZIFYSvBwC/
iR0Vybt3ptd8lItVv0ofOs78lY5K3Vd8z3o0IBHcrVTCU4kcUN0Q+kz67ipHrb53kZ5hwfquE7oZ
wwm68RNOnbgMtG1Jy+jwa51xUBdBxQ1cOGXmAIByaweL9pX2j+Lu3PLm6FYDn3Dtq9r/cetwlikr
xGg7viJxJ1lskz2YIVwyYJa4+mqueq5BtNaF8sayxctkJyEgRb1SiFNoajLyAqxEdx6BvWhp3q5h
7CsGClqJRyBZtkQ+YOHeWC05pG3WqOxjYtdACMB/wLh+fUYwCWQQl3Y8nRLkf4tauBfHgtvJ3DGT
ogIYc0Df7G/u5T1W5LACbpe4UT3OJyFoLSRD1BIfcLeyhyGOZc/h/RuTKCjsGLUxcSBF/LEr8uWh
2VRni39xLB1Tny23z/7wIRPayZL+aG6HJ8ei0QKtBmp5MlJ4O4CbtwV7zlPU6Y0btSkBulOP3QIS
zJIAubKdaKkjmmAcmySLqFYCJaIIDgIVRnS57dMq+HIPDHU5jsZ7xaal2SXEPWCkjhOyyxWmr8oj
E0kQO7gtBvK/YsEcp2f1hxt0s7O2a5GN9wp2jlsPmC+boZryIkX99RnHNd9TbmxhaJWjna5NOiPE
0JzV0xO7auEy+KOYZB4cMqoZ8o9SXPYlHBdSQJVezZZuTP3XRblAlqU257XUM6ps4ZjZymFUOrGu
NoKdDJlMjOE4ohIgZLF+KsF3zlt1KmakkZJTJ078Kp7cx2bmQkhkU5Ty5WkiUldgtGG5MZ29EYsE
F7CBwskKIFM+QkbssrtinQwAKPfqPRkJ3HOnz7h+wENxhiC526uiK2V9LOt1WhrWekKzdvVYa92z
LIJmb23D2RW1MlmHe92iYf9uO5Sv9ESMkjR9tzLONbiQaRkiiC5vW2j5BzBq9Turr+b9UJmPIEME
x3Im3BdpgA6/uF8NloEzeIVL5VVwVcYLHJyAsaZ8yyyV6G98hAATMEtRnJv4qMdFU5WL//KkZg/N
KNtAcxwHzXMHrpIa8Xa3ZekJ7oTFv2Q6LOXmbriRCn9/ZRaep/HvXS9/6Qb5C1sxyzd8teEP4QiT
v/M0vlpdJAeoWbEfkepvjhiCGIPLmH2N6IaeErqc+hNnb/RLeK/Cz1G0Cpi4Fe42Pnzd/oMRlgWy
632nyT4Dyjl3QpvU3kGTIfmk0nDdS+/nrjzacxo5yoK0V/eqhOWm1/rzgCBVemaQztsnvyK+3Z+S
LSGPwr6wfShkpuG/MqoW74CEjMZaKlXl4Sc5+3I4xkrAP0nnsGVgwlmMk3F6DNqmjjf8AJmsEqFK
zjyXKa2qM2S+Ju5lkcdEzTIhemk4JovY9Q8t0Vz3u/1e3V0sIOFtQ4Gx+6o5Ouiyj7ZvvVuskhmz
/GjRT105fHTliZDirfcaHsJtU2pgZLcgPlylQ+tPhknRoHDcm4oBmXpt6szaVv7WqwnJZIcJOqEp
gOMd7jNuTDjIlRc8kgpguQQuWh5XanwHFTpe6cLLXlnibnqRw6sacb9XH5saSk4bOZtprbDa5Uku
4uOK5qSaGqXRcr9dlYe8PPSqkSFfQUG9YfY5+bsXlU7kuUCL+S0Yk42rqOkJizOFH0Y1qTjftU1F
uGhrQi6Ed0s8cue6u/1Ouj0P3eVbiFAsvBnm0gq48VoXR3iA5TiziVgu+qlTITp47p9eFzRenUoo
npcfZ6fkzoQyGBVNTSNGlZeBqkR5rDhI8s5OTwrz8AzT6I5Y3RIi5vOmLEv0VrxmhvdR9zgMcLvo
dpyjHzMq9+yqzAYdNKXsxcYTRGromJJwBvkPQvODP6ScoMrrv/CGyr2HYymlYwXEMEDIt4ClSpj9
1wERXeV5gS9UBSpgQSUR7MgnDXqVllmBjSiCzgQ9PhwCtHEM+rVPhGXc7caUZzsHRiospBXDwRmc
U0+C/qIZ2xq8oyxwgRr3tX4yelBm3+qiiyYsx23WsWI2GUl7aFnOxwPKCkse+Zi6WYK3zLcbDNkf
p4u5Oznvsaik/kMlPIfaaQ8EykeA27bUdyrATLp5JLJ65IPUiRgmOWXKzMKN3I2yL86w3nQi4Qyv
Uo0VYtbzEK6+Hc+DexcvLUQATiokCQ1wZVWJ/s5inhUwDkj57ALLqXy9cyCFVVcwBjhbm7ERC59x
cu5Ph6OTxqAo9kq4uXezrcMBIQQ93KZj8DGPJjtjvg26e7xVbnXxTUgESwGUjIKT6WEWhCoFRDFq
VFMWup3V3h7e0NY/FzdAc0u5JJvmbW0fDf8bz2w3VxaMHOPqFrKyjBt2Om4xwXodTXZFJg4vNcOZ
l8yHw5IxdX+5FtMFbUIuuaqTy+e/ms5NgCDuj8X5+8hWoT0AshJXTRNuuc5JHfOx0XMAmeS+RHxr
IzE1S17jcIPgMhL0GxmAiiixZp2TO+zuO5Eh8TKJ+sAlFmUiKG9QKsz7VVbOPnu+wgg5QrR38w+F
n7Qu2NNykeyckGyHpc3KbTWaro5mUaELQCqnSKHz2YV6m6ZtAPZI9AMM4F+P404wk2hq55uHmwDk
A7t/RuCVL8FIHeMu52nAAAwKPfkM5X+EOd+RTjWkHsswvasft+KkqSly1W3HxH2YMc/DiWk+Xv3G
mJqf3GqB42x4SERqLjg/nlq2KF5v6DoXxDfDJzNUusPThZKWagI2H+WTVNVYVAEa1LRB5fCCh+6l
UGyEwdICJG+pC+8TnmxwFy7waMon0y2pHZxeTUoDJA5R8Yzio0/ohIpv7/wwZBVuDk2duAOiqlpC
xJfDzZYN5bbh1pes3HAlTv2+tnsfor9aYTAMUDqvchvuFYZNdPs7G3aEmKdjoGftTD1P6Iv/8Uuj
twVW2AsveRKqmfC52WtSe3FVICfZQElbmYwRFeasiA2aYmrGQiJE250DAOMxIGYK7Wd83z1SPUKy
5n394s69PxAO0M8f2lXn4uKV/MtQBSDkUKkOYMqh6ZoNVY1r649A+ksfCoBVL5bYnRvAYNcTVOl8
Q7CusJ/xPX3s4tbIIS5AnVKdnogWUk75GaMSLHSdPnpeDIh647V1NMaU5Ds1dOa+TO20HXkewyux
0F/gSsgYrffnPDUHtvE9tHMkxEuY0iTN/OKbuyVKUhltF+b7ZPPpiROc9Zgta9Ozj1p4Zp1fHKSi
R8qOT1PKC3lvpDWV7A9BqNFvwhItvV187d+ZpdIIyF01SvYOEotsbSgn7vVq9ISs5PYbqADP2i0w
FFi0837j4YQxxVgCnDoFxbP7i693BKuC3EyHBD67z6ijtsyVJHnN94H7TM8ef1kVXCRc4GxVX8PS
PcBs7fwfVjIqlrjGkGLbvU5bFLtksBSeTr0TisyPJGOER4/p4EtDGPUtYtvK3U618/Hi7g0Kwpa/
MHYu41yc6cdlvUIFhWfVjm0lpXQtsIicH0oiweB5CP2Trcau7XZ7sMG00KNh/XV+RgIMyCYxjlyb
rsAeZYqqGS9HZc9GnKmREXLGrB9CWoMBKrEy+5OAYjK4/zAjUB+PPLQGqVgs4sUvtTT7J7Y7v8YE
Aq98Uf4MXVxQFUQ5ddXStD8UO3mTli/DCIjTCEc+gtfm84pvzeLZBg0qWaxZnMRcvaLSQJNvPyOY
3FYHX2nIPRkRvEl62vYEDLZyQ0lQcCp4RIUzQ7Gul30FNH+ITVtdPq9mVeAKSotUqdDeZM93/++5
AC03pJip9dxAHKc3aUInLBvxu1iuD0/DWinURW4f7rKYMur7jNS42RJGE1M5XAA3yCm0nD2Ci5y/
1AiuONSahbNCWkg+BzUfefHPLvyMOPv23P2ixnIoondYOhwkyJRWw5CEF2WrZwlZyD2P93bxs3AM
9lRk1tGrybomlVHZTYe0GBvP+o8je2ycvc9eo2RQgcMlXxFzEBZqRbfAx4Kzk896q/RxC1hRVtAj
r9t47y4IophQjc9xqPbq3Y/zc3DM9mtaNCwqbbZCkC+YNJZWHm/DHF8cM/u96JcjbHceT8mhI8k3
ove0ox/KEWNqsFddWGfINVN1bK6txQEG5lSIja1fQSifCcgkdzz4ZjdCHG+sessIsvRUsGhq53cN
CSObDkcurE89ng3EboJ8PZIb1l74qWEm7H3g2trXNA1WR0kWBob7qXBTTX/++tfG1Rmhk4W5x8RX
1Yj8N+KiGvvHDuqqBIX0GU9ldpVq3WVABX/Fk8fkV+jnIsxEkKJjP0OHZjx0pcSELphiTm3xDRbg
zHnn86JKxAQ4QkuL+BuCkplLxm/Un7KRns0GZNCZSAHn4iydeU9AAJAP1P53T51immiFlsdbb5Ts
sq9HwR/EZHulFr23BWRaBdWXrRABd/X6Tvorc9JHFCwn9e2w+AAFsvZ9I0GJ+zQBhu1QHaHcYkPV
8nrsLpGN4SYnxifuba+mbLHoP5ZNeK/2rbrebRj5Tb7APZq0W5rK6R5rkAy16oVEAhoejZBzRHqv
C8EzMym0Bc6ZWAe9lPDS8xc4kHzytD8OtHbDAt1erM2xZ4iL1Ag/vRMkEfDTs3b0Ke+tgrxTOb+h
e2SjT+UqsoP9JnuQctYY0RH19FQP2LnBXqlzz1js54fCVReXvV02xIa/L5MPn5X5laIy4q3rpX4N
uFzrvaXu+YTKw86HyltBmcEW44zeQcO1ZKf9h22VIqUthg8RukYngLBzMY2BBaDaFmZ+alNE5jwj
Wa6XNqI/I5CLh/DiKuFAzVpQKGJF5rYwg3qJGz1UkR4sKn1xNVs9QO2mmzEVxzFwogZ5croQTgjc
OFeLzBlunVhjdlBLLqUcjKuaHo4pzZzENhIpo11Up+6tb0H61TS2HEh9p/SEUfUW3vKZM5mGAAfp
STBZC3Ia//oNnpYBNK+UGkN3fIimQXZ4X99fnHRzWCXWIoL/z8Zgiync6HLKMMcSMHfVq1OWgpiv
vX0CHgeT97xFjh1+LpMr3qy6uJuESp3Howt9xmlGhbTADXvvuNJajyiq9p7P3GfHnthTjy2aGAD6
ahjxP7+9yIv7Y60si6b/G+fHqRjhe8HlbgtFFWzkDezkJnskwxbnAY4Bs90OpB5MGZULCXIXRcgZ
3EQWSyNgBe+1BPwi+5/4F04kWc3Caug1hrQTsUyO10Jk2jvqUVyhnMh8sNC9n/M2RDiSNT5bwJTi
84SRUYB8MYx7hWnvGs8TUa4c/l0MALuxPrqjAgshAJU8od72ASZkk0Ep2ttmU1K2W7M+t9rjR1Dj
ngL0KeLPN7WqUdHCQk9m32+JRqrM2/rAOUxFM6KDoa/se+J1DC4fEDlV8nJa6KG6pYhYvkhFayaT
sztreP1JtrYUXCj2Ot1iiiTgugOal1L/K/i1byMX4IuqI6cBgy9ztenhBPSrZqjCDT7xWW/PbgX4
zFx5RB8dNVCOJqcAPCbaAW4Swiwnu6fnhbS4c857C44f/Tb+Cqn5NXVNE8/WNBYYBhI1p6jmCE1Y
6YycWv9XDvcZB5+SK3XupKmyizwCUgxtMxv1J3HGuir0i/j28JfaaqiEjilpWB7lbq/nrgGBYErh
eoEyliWtBdAdH9olaeXc51J1UW4AMqy3mplCVf6LD4utmXCiFwOarYpoZTcBaSKRhYh+Kz3n9XKm
8rD1cUE0u5tod0oEKmsivEo9Cm7uVB7jG2YiD5oBZNMDsEYyuR2Mm17uU+/tijlKoFQxi2bwBlCS
yieXAtvuYzh/j1iTbd2CeBnCfw4M+ryM2yKCV6oh8KeKuGsvCf8daZ6EWQicOpbGSNQfJCB/1M56
Pb5FWpOoqzRJvj3mjenr2Rz7yhqhsgji3Bu6br2jyCDVimgr2CM1na6gc55+bysgD5ta9URG68xH
hx1890ISCFQyxialzVFR8FCSExf6ZfAJlXPZbPUsRpstpqPQowpV6PRbI+F+ZGCC+TD1IHf/ccSM
ZQniKap0riqQsckwjH/G/xNJK6RgJEn/zmhR1uPpU/lU7PwGThgi5NPcAdcyaZZ/h+g25ZIwm2TQ
aG3pqCQI1koRAOfDsh3HcACozxPSMCa14PNStNedS6s6z2jMwcaYcNjJqivRzwU0OBnjGH1NII+4
utJhx5Wd/Yqa2RV9aB9b2NnvsFyrRoQRoY/jKDJFkoowlPP025nKJ6v0wnO+C0De/ZUoOTHe9G2W
dVoYny/bIJwPQ9EA62T3PjiEo/LGy38jdriUb1SAD+uufScKIMniHgxyWe6KC1YZVWiATntrPtis
gVGKTNex+vrItwcMJwztA1P0H38UgscoIjy/3x4qy49eUFFfRvlQGR5xCYX2huSJPTFhTsBuaL+k
Nf0Oy9FhGJ4kM5iQwO7EMvza3tt78EgDHDYsrZ9OAiQmC5Kxe62bcv+HC2z3dCNFfTMqK+p4tZtQ
am1ijZHqRntmphb6Ec8usuFrd9zVgwzfNlpIoAUnxYMhBnizZ4WHkGbpJJo2q9dz6nqm+4EiS1Cg
/7u8fe1vLkrV74SCvpiWWN3s7kylD54iL8Fd0p7ng+aLtjP451b+ZMK1d4oO2tTTnMfntz6X4FBd
g60vxdpYem1rPyHndCCISlHahhV/MbfoS848gafpkpRPIun9IyEXibRsrZgb8rVnxE5LIv7MVxVd
aZ7NlEIO0jbxX3HdfVCaahdm9emZcOziuv9/zeR2Mi2NjQpXj68hvq4aHqW59hB5brbykPXH7TrR
Ry0yeP1T94WKLFNcxA4ZpNZBiyZemioVaHJJOcREKHMcGp+Mr2L9k8a1aRtTWIagE4Vr7PBoS1u8
uusmEaLX5QUkOV+rISe1FQFfrtBc7cWFQISRNPIa3SmlJ+n6i0vShomNHQ/uoi/vTSx6PY/1jZYK
OXvUq7JABxZpXP3GMH3SQulGTb3t+KxOASLECDfteMiNTRCh6+VUkt2InX0Xt7lMWJF5+K875Iqd
qybyFMwB1UzB+Mj1oeTMZSEtwk6/5pd2GixvBEad/S7u1hYGGrLcVnjMM1Ek5NfPZWTSTnpAZSIz
zn3Cf8TnLC1CbSZJA5P/IDY4eEU8BuSkEGdlsvjdeCn2LElaShj9b/RQg8FZKGWESH95RWLqijNx
zup13QcSdS/Z1y+D/ITx7ruZyg+6Y+XA2nK00cDHydDWYMxpzr5OYpk5QWaa784rtJUpGRDso0h7
VRhMStmbUS0sKSPpYPUJwXtWUOcSJHVE1KslOREbppAla7fuSCI3NEradHveyxR5FRcAVV/nOhKo
vI55DQXasorI0a3Wwuy4PP5D4DcuzrawStWilbcH0u8AvblPPtU/TQUNYeyh33onAvjW5XZaN2y5
t2ZNAl3ovTWeNOuyoQKKR5I1qO4j/c2WwnPewNqnWl4V3oZ6k7sbaJZXN5XPdbbxY2fVzlbONJ4L
gETGQ+sX6Ci5UjIRLieKHB1A8+I/JlvNqcBJIf+gGURT9C2ZpZMdn43wtLWD/aHinJ67oQE9O5qs
/0ziW9m//Didj5kZ3LL+Lt6+I9D9MnDBIykeFyO38bzhQjVws4bSVArNMffEImAEy4LdFPBta48p
SI2bVjU/MBtjjYs/zRo08luvfeuif/HyjpWCvD3b8EgMB0Pk/8qoZzIUdEk7gUci6XYQSA/Xbq74
A/rCi8bF3Hi5aBqr2cZFODM0rz24ZDSPR+2tLrYe7+SHVA0auZJOiFXw2oofQV/HSMpP85toHEsp
35He5VlDwlqr04xNbOHWDykwNgUsGlzYKJs7+JM7tPA2LBI7yld1C0fJMW/wlXnfTub5K82Hp/T9
oW594ijVTL22nnzcWpRhJObRPLKpym/PKsBv66ywCprtWZyLJaFhGBn/bRMzy4/heh7YKCfU6zl5
3UEjbPyvHeafzZStSJDJqYumZEGpYtQGKxydsZHXNKzBk55OWvqZGNlLXBhvKoa20WF/EHEu4H/T
T0QwtqdplpeFkF+8RDCL4nFEMFqILBmusjSzQs/J7AcfKP/mMI+WH/Lk+zEtBxjX3G2o6p3UQM0l
2cqNCXPIISIV28cQphtia713JjCa3EgS7ox2xxJle1Mt3z3xexuD3/D7fC/hOPmzoLssKW4kjmta
PZC0q2NC3MTT/emK6JUy7nIhaSFQ2W2PYxN0sz9s86v3daOj8g+YJCS2UAVJ4SOns/jmqLQksf6U
ENo3+tVTGWS26sKSDUlDDmTb6TJKea8LG+2XnQKX5+mr53DuMic8upyUKVkRlU3Pxg26ToVSooVx
HuXKKrb0h2ZVnhmkDybzGQsH1ogvDEA7ZOSOxpRegQMCUwhhPADxOphM9YOLMLg2KTKsK9vhize6
Eit7QBipAQotmPlP1IzfZqRrUS08E3Vf3uKt1cyUeF9Xa9Pp3WZtlAy6YvcQjGPU5eb1rL9s37TW
+4WrMZ6LRKl55YQtTQ9bCHOKbo0kVyPf0IPODBLsG5Rf9EwOXhUwIklr9lNtBa+9mBLy2WucH4S9
FuGVhug5jh2qhf5/TDEOrGi+eEV/WcvOWjki/pu+L8OuGFOJ82uLTmAdumoSdXE9hav3SWhBciGm
pMoGMpdb+ECafuuc9yYyBaW5+bPikrSAgdmprSVx6RSsHIY+fbHBUxehfdiONVffrcJRAT1om/DB
5dfUxfFtznT2COxEvKo7No4S66W6/e49CkbfqHGSKtAF20zHj1rv5ApYPMR/X+vaHhmQFMP9A6z0
k7OLrvB+5kp7nIKEamQRRuu6cnDzmkef+P2CLUxGeQKlrLAs7cByXlT/sI1yUEGAine1dQU1GHEY
Ejwr0y1QjN6x2ZVY+gfXcik7qxIqqEyqR5Qv7By4uqKx8OYfrK6QgrZbBsWDVsEffJdsAtbC3Ne5
AKRtXVMtN0YuFeTEXaXiJ4DBlQSp0rfGN6T/51XvQojRECSk61NcZ4jvRDmLrzwSESFzh2P167yw
7C1k+jya6A1kZS5/wzcWQ9I2pRBDJY+eb2EYNESCNkE059zhoLeEgTOaD6EHn+wrzHloPuEomHgL
ZHDHpFlG+ue40bPaLQvGBToiT9A2Iipv8b4In2RdYn3AjG2HFBz3+8IDpRiGq6KzbY3RYHfY4HKf
dJ9QaA2AE8/7WLy6Q6RH4dI0HEGd8fOeAusrbcV4QabE66piTqrRYl4+s1ewvm6ls1JZ3E+ZWHfc
0s4qbCH7/dgB3ds1VeaD9rH1tP3qWttZYIZ/jeQMX41rldtzEGQhYRPA73qFV/tJlZoyQ+ofiksZ
VAggmoXUnx/Ko4rlto+/kzQVUN28CDfBQVCjm4R2jooskLYj8Kkf/NVyXACeQmPSFDvxHtgp/AaI
xbvYUWSdEh+Bn0J2fM0L4+zutb/yWE7MtuLVNSFdGYj7S6cswqVpq5aOGx9HPyy5jD4eMmzRg/AR
4pj7qu/mpy/Df/iiTZp0REknffsj1nzvpspGhFq91wGXmDDnUUCOYcgqXlI3bj0PtIlsU4ZkIiBH
zDAULBZTXEuOdZQVeI87hTGJSlrhk0qV3CYusks09haGUUnnt9tUqBLYEPXOjWoyEEBaal/tX45r
c3xYHcp6MhxuaybDlyKkTClI5jL0NAsxUK951jlVRiQhhwbeIoW/Vy7+YBO2ZzZha8KqPiCWFAm5
HLMh2aRY6irPtgd0Gl+JLnbEszCo/YSYPMko9EVsJ0teeIwpXRIasx1n1B29JcGzjSck8WF/iAwa
NdzthcPOV0tECHLNojM7LjcB+lCakDZaj+4vmEQkn2uO5C20MTn6qlquFjUmdDSSa/PoAZnvX8Zr
b8PhNufJD+OMcjL8r1ETbjQOpPWYDJIGz/HJ0OBelTxvRSkGzNbQviphlUC/ewAfQblITbDWH4tp
hXBJfU2gdl9HZiY0UVbkc5dtPUNFxsZuJP3SyNSmO7yRGuPKg3gUuix5B5u2Iy9oLAvOEBeDgGbj
0LLAYV1GrBmeLa84X6bzklHahFddIAgMt/uHzuYI76pQH7dt6w6VMBsutLhOc+95YheX8zXgi+jV
OSEpxucce9a2kLq/1XlBa6lTk6qsmx3hk3wErsUx1xQyuhzLQh3KcXuj4HWjBWKlF8LEtpS/W4Jv
8HXnlTOaCQvNhhxAE1tEXNc5qdWfMJDTdf+IlcgZFW5lapAdG6F5W+oBiSw7JZP7J6jgWMCKgQB5
lYQCdcWdf1tmALTuBzHaSZNpJMQhvCpufwMwPqutdBTpAwT/TtzMWcDEaidSR1r69L6443DN8Jfo
P/Cwwpg1vWiFdIMUwHFu7F+PF4xxTZe/QG9PBs85Qgvd3N0bgMbq8Wc8WXeRrcq2QZ+xj9t/Rm5d
oFpogz63XNYudq+cC8i875qsYd667dDGxBmfEU39xvLKNDwnA6y5DfWym3t2xxLbWk5PCCzRCTgg
88siBKYqD9jrnv9bvgwilGX4ZK1cvOVy36u53QyfjahNADgOjmqQHQc6xrRM/8UY4rUwSLDZ4hgC
Kiq+PHGhxOhY7VJi0H4LZZGHV53tuNLnD6QMn/EesGtB1mxEuGdFJLkppNJT1ydFO9xNcBmf/SCZ
xxk8SkCoFNnpk3Uo9sTohPwutvERbqxtBCj/LtbXv+cm8vOoMQaQUDHWfXzm5dBN4FgZpOOmkn7x
Fow6mj7zp6anKsYiB1vSzsl6uE+jkU15EvCXFo22psq8iIrCOBolyXSs71nuFah3FVpwUyRfXbLk
S7RfvBhnUybJd1C6cLSCq0Z/Ojygc14vkzlrOv6RlciIh3oaMuM785lVwmhN4avkTcSed7imVDc8
6q2Ptwkm24zfJFGfvoIkFtAsCJ9JQOA7sK22jqBxEoeIOanA02YK9hVyzNQKqDyV4FTeoLnbNYO+
RMeLE9zmU5CR1F2Ys3nzqoIp4vJB7RMDJ+2uuH1gG7vufu4XsPmEuLW5Vb+vqr1MjsnSRX2OadM1
9uLTvGFN+RTV56iP+KjD3ClEtUn3mEcTIpSwG9iUFaZvR+mhPqogIIxHkZOSpE0ZlWWncZNBSoZK
pikVhjXWETkAiiMzaGT7T7QXKCQ7D05XwoxuOqfxEgGaeMdkCEW0Ucgdjm2rC0ZGhMhD5JMjrldd
WI1YCRjTVeZeTMsiurAbtYD1TnCe49yme8lSmojN/8e21gpixf0V1sIcyWYoSLQGU/DTsTFp8acy
PE7GiildMnGQpA78OrbhKmHhqiF8VnuD/94ANRRPAm/CmKPz5qOJ/97NhKcnVi+IyrUIOU836dDC
TCtxTL/UUPvNTipOmXex7pThUEQO/t7NcxsHttBAZ5nrDJqDRCkzx5JmphUesbO5RkJl3qUgPOu4
1kZ0ATeL8sK1udA9RQFyJZy+fUWayEuN50PC1BnN5AO+zLWNfRHAgCqRwh2xhtcgdMsHxQE0XtpM
csjglLhZFlNHzyRXfzo7EMfTM6Qc9UhIrJ2ndQyk+02zszptfJCE7Zmbe0vvbugj1F6gbFdv6LW2
plvixVCcGLE5t+Gt19qQeuzO1wkdxqVe0rDAi1xKMVqynQdFydOFJc2ekS0c/IRt4ilHkXR64ji/
1aO/QopMZY7WEG42JMu08ga7S683v2r52pFzUsmv9Y8tgJYVFWricqglUZmT2UV6r/1v9SAHfF8t
5pq63P95PPnvz7iSpk96CGr91kUIPePSds8qu+vBvmkJOg0CnHubZpk9zKE1Iiqo6jj2CFOcfK+p
/p63hkbEDctngI1U2XfA+10dh2afY2eNxPPVsxkz/8L+3ovQq5s+cPUIF9wnHXgsnsStxrRXvq5W
5Pym/1wXb78mMNV3YEzWPJMIimkKTMP1hcWwmAJjKthHTbglDFDv8wQm+rXgGnja//tKWaRMb23O
ZmnVG6mfHe+bLNBf5KW/OVbP+DOvShoY794hPTpgJ0sXYsrvZY44ZWF2jIEdwoAt2X85QwcXSluJ
SzmTlDiGVQpumqFltr9UgvydmSxhnxhgSzXRcs1aSqAeRQEezC3qJq20StoZ4OhK4hvkrcstquhw
pcXPnKfRbxUUxTKahg1sTjguUcnq54fdN/BpBDSnJMk/ooqFJyw4SjhenA4qNds6wFEe7RPfvYLN
UavmWWySJM7zr6QDVVm/YfZScSCwcz7E+aRpLW3cLlcdQga/yhmuaeF+Q8lxxjLal/qUV3avTrz2
i1wGfkVKHoP+paATug01EpoyuUa+f6kkgr6gFsco6TxFpk9BBFFpsCimlNq23wyrWIgMok5w0pM4
Tyjwqyu3xoePlGL5Bvkk80z3wrUFYvPnrvCiIoAFtU8O+j+NNoxS4WSww+Fl2cGe2PgLtYY3wshd
wq9jSFgiZbc7wTyJVRwbP1b8NV8wX7THdvbLbaMfuEHD/+UcloZdBxVoziosaeIsEfnmTXyvWEZO
shdVmxUUrfzcfxVmzpx5cSoWifom8Bx3oqv1OG5turnBzKalz8dvWwbLYv6QDFbX+twWw7S9E50/
w10ad5l3PUJ8OY9qptmzWRGdK+3E3ouCFtlQv+aon6yMnQmuCnLzoml+sKHYbzKio/45VJpChoj+
AjQkR8hn/ql73rUoSUrb0fTjAO4FpEBUkgA4CLKv/9mzH8yhQMbXYu8iWrJ5ihjwQysH10CQgwje
+cPd03BkCCdZB4gBwWcz8KK7socTqWYH7m+0p5bjYnAfFcZKsOCfQ6e0AABi3NR9xVAU6s490ZPk
p21kzIsaqsYEUUfxkCxDwcMDh4rsPb4Jbmd/o85i86XY9382PEleDhyO6nrZVZi1AlL2JgUFhp7Z
bVKnpp3J6pOQJ98bHg6EeBDBb69/IagVVFQA7LubTg93KAEifjujcfgUnVehfPIDbaApeHqOTDJn
ygHc2OOoO3XBQwV4lLMdmkDg/9rgCeOdE6w6pRUklK5eOkXFZlJtZfyaiXKoz8H++N5Seel77Bi4
BbH86Bh7rJqhX1PkoNBchQJwPzErebQ1/TNDVUDEV/5k+b2pu4i6BmKOc1F8RiLLObRnF81fvCZP
fIHy+3DN5ej95lT21LrznKCK+B6rtpGSASJgSIKqrGC7waHa5SU/pP18eNZCinU/xh2f7GbDZyDX
2pBlfvC7UQ7xelUj4CaFkWLyX/HF4+b60TqgwqfLFiTwVcbCy2xOhw294HGvtxiOBN1e5QzTdL40
TCCeXEsKpLtvyslmBR1eSn5mDOwG0c9IRX8+YdfYBpWGV1pnJv8pli5kJLZLZHCUCsGHbaUKNLPJ
DWsZewO0GalU17ekPN6N6fS8dumwZaYGNO2hUkz6rzm8OfyXemu+XMOamj/N1xNtD5H9tTNRfp1m
8bLhrDslxZkX9G5ySWUrT0j+07qKwwqHAT+GU05GO5EyMfTOCWTvzRyjzXTztiv69iRm6z3gb04U
7KL79HmC/WWFj+8dMgxlfJIET4w49w5HEu4tIFA2FfMDW10YOH5lOsbHK0yVk3w0dTbk30yhDDQh
wwnV7FLo3go9mX2+vpOpgyechfgMELYvyhfXFIO2rwxLn46x/ZcL8GG4S/WFy4NaQ38u8GHosLMy
EGtl+zNq/zrhPJp3VkgObe9wG4kS1LYULGhl+2xOL5hhPEmoC050XCP/RR8EgY6BnA5AU+l/TdDS
vW4XwkMCbIOVqWrita4hXNTT0SScYl3t6hGh3cPvDjotYjUMf4xyIOn+i0ys93r1A4UpbH4+Qlqy
LPMs7X5QZ1mayVAvlfjrwJaBIUfRIoGfTrFYcpo2m+I5pJJDsLf0GmpA7PBLmQey2nTtOk41scms
AIpD511hL1bVce8ydIx9OlZW445e21KZhbOljoMlN5xHYBABSygjc/jDz59AZhtCh+UbteoZ3oLM
/ER9sTefmRW2f10ZyNepMpUwb1N4CTqmKJ0rFv5/P8XvYDbsUnWxPyirMDlt8c6FyG5AHl8UOVFT
cMQmR3/QdZ1YSn3jUl3qucYvTfMuvFM9rJ5R9HGP4/9sOeam/dJB5jKIodNG7smgVD0kBXLV/6fo
lTQgCHiVAj7b0i0qDheF/AvN4pOxHQiJ/My81p61g9HYvkADLByqaCF6LB5EQB4Zq3Mk/39ASXA+
YScWOUTh/IZ1fIQ3zXLxlCzYYvbO3dyG+/PxIPntrmpg1J2Zc90zpLyyUz+4KxiLVXZa9FnNHm46
tB0wXPiemyNAOaHdhv0f4S4n4Yeinio44h93LY0F+0VnGVPExPFQlfjwywbQxD1DDOuIqtHufhde
n4/NYVINZMOHAWIsakG2mZEbGyErC8g50fWmJaqOaxstdsIiX1UjqmpKAslY+Qk+AEKYqThhdrcT
RJuvOFrUoLuWhcGrGD2DaijJMOiqNZa5wk4BwQaJlr4cRLvXXAmRDs7IpilQV8FhahV5SoVWttl4
Ne89JLuTq+z44qrdXLXA3gNNCG+ilGf2vLg9wJG4S0QgscDxUcrxHktTQDXbA0+MpzQFEa4XumeE
6dN6fHiYtzlVvIRKBEyJk9OVpukbEvqMmVU4Y8KxPU6KptvdkgMZVDUA2/dBWL+pkqzo66N8my+h
a/b/NYg7X5Al8YlSO6scPEBN3Ag3gww2qWyZFwWPAyXc6vIy+yHaW4Ji4vyd3yWwQJy81pw67cSW
VdwGqgY6KGvZESwVQyQUcOwnXxgjG4hdtUkCE+DxqtJnH3F5YQITdSbVLEUG05Ohzrc+F4TibP7Z
SRlIOv3SetomRtV0bzmej5KgTI8ZIk+iyshBesOKOTMJaXBBx4E/1aQk7bQ1qZq7kDal7Z/XVVny
WYyy7zm0B3FGrSoKV+LiXiDkNmd4LuQeh4bFdfIDNWw82EKk+hJbZ/r+ljFD5ImS/y5EWx5Tan2l
TbsMugLDXYkh+wPocS7iyszA9wgDDQIuUh13Q3I6nofwDm7ugvkRzP/UdcNChO7km0RGwolEOfP5
5LurKcpkpbOQqd/fDTvtuXBiFRTqrT7cAjAEhs6IQL5PH6UTECl2QLPj/GuIQDp/bZEpyZ4MaXjZ
MdMm4CDS3VRNCiij5g/XdagROPTKeyVvJbCKqkSAiudV+UvwFGzeU/JRt66f1SbHv0/XuKVgSeGr
zOKNbqD39BdiiDi1mEtgWQuZ1awrf+yWAgISPohyb0QqH5XMd5HYkN/su4C4BCyHLL7RYaHq33AP
SracraVWkR8/QWHdYzYUDQTDthyDFSMJ4eL4XHoJI5HB4EsF0kUr1HaqpIEoInQGPejtbYMcyn3S
GJUkRNMQUq/pax1OeLw/DDdcPNHQ/M7QGZap8MM/7VT0Z8S4VU7wTz9YjYHTg/adpobZI1cIVgrg
ZsoVfrCPB8wQwzkXG2xQp5/43+hzqR5HGfsiIO7X57YUhhKvyg/fFBT33eJkewAhNLW6RuFgsmfl
xTHqqo7qj3U7+y7MuQqufwy55H51pz5kP8EbvQ3lutEcStajMBcVJ6jFbMrFrJTskLI+8oAYh9nG
ZeEKkDBrrgX6/ibzM6/pGaDj9Pui/11vbxYZbAiTHpUYlpr8OIFeySBqff8gLEM0PFHRNcWTEwp6
BYIA/Bs02LaJbmWo/xvv9G+k3GQ7Jq0n+s/Pv4iqa5KN70TlMGRt+RcSS8WSfMBBugypUGN+QFCG
TZjl/yrhV6WnEl5e50wQ9ajvMSLBNpgEGiAcC1eYmrg0Hjljx17c+rlmu90rrsFiL/cyxtSJejbA
RfxL9oiUr3t4qs8+fBn8BGjy7iFCJKAXMa2XGfLqyKS9Tht29fMT/efAFsnV9nXb/EPcPe1/EaA8
U1QcxVR2HDz9h7aBgIK3eIajyPKFtyk2hQRrkckaM6PdsJqoj78TGCUVPHj8P2HyBg2Epcw7YplD
cqR6UzUztHzohu1JxC4d8YOWAp/D9obopdVm3f5FO1OTdlBQGNhIVp7fwHouPDmvrkNb9WruPddk
xZg/zMEiLAC/b41Pa5MXI2fgZz8VJE5BX/lQV3Dqq/SXHWH3BAkFd+HsVoP/8oC/0EgNtrYCaIPo
p5qvdlSChsfOETTdiXdB091CURnvppAyNeyBCfiuiwf+ZQVHMhVXhyWqynKHkMFL6sHcbteFQBU4
Q1KMLUgzpHyywicksjzLalWqfQy8K1zxEk5frL5iD9MetLS4Y6YOyahy+bD/Zc9T4GvNVCusRWno
yU7bYDS76ocHuMHtNOw970rbCbRpnalOAhRHgFbahHTIsiS2ZWvF/t8jItq1HpKzMtLu46c1B1I4
nlRNSdBuZ4VfplEl3mq0OpbEeX1V2UwJpAD7Mldh1bB1KMcxSN8/+v7/lQtIQr1E5hndZkajglLj
zVk+IhRrtGy97F3lEoH0k8Oc4HDtxpbFEXuPB6yGk57xENGAjucHtsAR35hNX80w7UL9Bq6Z731/
Zt77UlA45RTFsjpXO1wYHxF7wmbUZnLaz3w4vluiMh7xcyvsDBqFNzIxDV1r5BfBC5VpFcOuLqbO
yPcGjuNK1kXX91QHxZwKI21sPrIGoTFSQYQTGcpYfcddnblpDfVUDoYb5TqOYp/rlvwpNfOZS2xM
U65WYuHYvmwTQt8Fm3HyBRSPsXsSaccgk7b6kPPiouiWnS4ApdXxY8IjrKN7wZr326UdCR1sN2yV
m8EwH7ERnhNfZlnDZjgDoE7SRgUaHsKcE5FYCqq9qSuSPAYNW2369IT7fmnOfhlUTt4/JQvXMMBN
qWdQg+/b3K+4J2OKUza/+eeDY0on1x0HQeG5qxpafTSx03Ga6VQiJDjK/glRZrLgDOmp7cYUIFig
J+4prmmF4Su170RyyWmvzIvNpeiefIOr3bAgSOQZXt24iOiPhSzKID5ITZULP6rmML91fLuinppe
Ut9Y9j8F790LMD7RZk3aYCxuyJqPE8M39Z+lYYGamvx2qXW9IkKrQLA9G2f5KIsVXnOgL8stmFr6
z5Iz5Nyvh+S/1gKeirXRhjeZxpDijvntQn5O+cQg0I66yvvIE1djQHzhwxST+j1Xwl/vi9zNREdo
a/J7fNebzsejhfhGAh9RyqQc5XEDBnaSenFd2Ktk+6BUBgaPyS8PgSIsd4THBCmb8ELCRpu6a/bv
dps/51QpIuWB2kFsR1AbHA1tyWS2DCV/jg15pZQVqy1hFbqxON4OyyF1fDwOLhlFrI8Wlwl87Y24
o1A+9EkJaBIzAz06+jYu7S73h+C340/5GWRFJZZVG92woOCjJIjIi69sFUFYUFmpbOwxpblYFT5N
XHzK2UJ9Mz6f5tlgeqFhbAHXz5lSOK/DH0CYmsZSfZB4NYdfmW77bNlw0Vhp/9dmD+KyB+wFQQQQ
Zw5TXK3bLH1/irc3vvIuWNGW+HMl7PXLuOObi/jPLjJhzDb1tgj2Aw3kV9hs0ZfAUvoeosThppKn
N2WplPt3yU/P1yA6MZjIsUvMtyH2u9C1b2ocRC/fe0XDz1+xBXSWbAZ14jGKG7Df2V11A0P0MIO8
hKEb9cMvKXW/vhWi14ZBX9RMJlAObeFHk7xou6mtS2MjRS540Y0YUgmMST8OPrQKTBxBaFaUlVLZ
ZZAYskhdIQuSD4HWW2ZMLGD4CnreDmPUgQRasvKbfN9BYJfkqD6hZqMSXSgA4NEKgd+sp2sLbHWy
l/CcDLv1eJIAGzv+6xuh2Ab67tQJH24D3WpEPERyp2lJib7RGw7+fThFo9dn7dtS1YX1T+fWxmyY
VXziugeAal106NYqTGzkPQrPyXDT1S1gjSGZEhWKD+SK2HJTkU0mcEScFvSHspIpTe925o/pFEH1
Uass6TJ6XV0/I/jsnIRXhNGgmKPSaMTndP6C77h7mHZih0+PF0aS4CVULp/mf84CXAeqbZnzUllE
yF6QkxrRsj68QMZM2dW+qQ5cU4dBKjIKwfAHPPKYtTat5cB1GzV3BjFLCnlkgje+T1FqSZmOcNtk
f6jBSKnT8ccTFETFW2H5mQBryBo7TY8HmWYzP9eTHFrer+xVIS/uhKdWc6QK9DVGRBi1vwOIrySD
dKkOW/WcsZDvHV4JeqIBBDQSl4SYXrxnP9iT0DhH4uRnFZ3TgKu3U4YUvIEhxGD5S1YqRwcUJpR3
FZmlXBcy79bxyCBN2M5tjqSveN3edlWrmUYvV17ACscdgTPMwmd6WB8LPgZWCIhuyWD0ZIrXJJ0A
1nJzYtWf2IfqEAiF0CJM/GmxkoBUN35ZzJqmE7nUHOOrwq4ru7wqo5X/KvEkioEz0nBK8+c3KlSa
qun+2UhuPO2llXuXMM4IQaj3NxQlUZ4lMl7YtErmaD/O1kdagrc9HA0StySsRqy9MlG0fjBMAC0U
UmxMlCLB72DnjULYluBC+mFzzk+rngFi6k7od+N0PCIPJF/Z1XbNpQgpZEl2ItqoTVEEbQ/PNMzG
Y0xksicunoc74rq5iXZOwum6EH+M7y+G/pdpatzXFuEVOx0Sx/8uUa4xdW1HHLiQPqbIb8h8kwpO
YgAxHs5QIXtmsyOyItiTDMwurVT1d+HDVagua2oTa61KCufSzhD3mxAmPVvLzeVbcY2xKjgN+3ba
Ilj7HNmnQGqlPDkBDW1nfC/zShUsUDjf8Ips+VNhQbV5cDfV2kx3V7O/wqJEEtOC78theuC3wySF
6K8kkIIhsnto1DP62nF0aIeqQ1v+bgUOuM9Eg1/mtq/5dVP/Er+rPXOecy82OuyLIIKlbREtwJyC
wj1lRSWsHosW3pofxA/fU4N1ZKz8ysxRNyfFe1MWOyMF9fqXNGPL3/PhzK3HgAZwTmhFqyfy4lim
CZZBEni6Q+TWfLWrPVXg0M7O13GoJmffy5DZRl5vQSGGcP1duRn/k4DAeJMtdzeN+8Zmfno7/Vw4
uyveT0osPNZBWuR+KydISdKW6EkQ3FRA0LhM6dKimVLQMsYOfLx6lVhO5PEscJVwkWR71Xz99ujt
wAtklpqdc5W1keTMhy+4wUWSxxke0/q78AmnVgLH/6TFw6zpxlSCA0Cxyu/BDS+GncqIWu2R6HYA
U8HlBjAtg/Q5gtg+2khvRgMCtrv+NyMARR/V8xEfD+XEnQy8wkQdDFNtKSD8OtvilT7asCe1P2o3
fzjwz6WuOerb9ne02/OvJqzYxePcgOs8egXH5MQan1xunzdHVCmt0RhTTGVi+qtlDrybzQRsbsFo
srTMvT5klkY7Ci8YG/zLkBvb6QJQ27CpaMX8tLqY/S61ZKfAGCkrkzwjXdTvDLq+Tfu7BfOZrWxy
6eq6GRdjkJP/Vvs+laYsngWpAhymlpQME3Mt/Z1SJZJB6sjFkK8gDXTh72Lxhf52OynkpkOivlJV
FGgliMWzTsRWBATwaCDOmVIITnHM9ip2WCIzgBjb3q2HvJ1mvLQciLj0SnwfoLNzB/de+vV5iCno
xxigxR7Oei/pWg8K2adnHsSE344zlWir5zw/RCs7cF9Rga06lc9TZtjqxN+5rDHhbWLrKwlicdoI
o9B4IjuwfQD03+C6M4pR7pz44ficpCoKFZa0MgKMnNW5+gQmfGWqmJBtgtYfgAhuerIeHnQmrGe5
gF7N/D8lp0MmXsl52DqZiSxbrbpIKmbmU4WkbE5VIglaJnBcDJ/t1FLiBsMUBVB5VbH1h4qNPXMV
24WQd2qNReh1GJtWY5e4gKoLi+WLePyr2OE1G7MZGfZWOIueKmyQnTC+eNp6N6eH11mFpNoIya3O
l5yv25mMR6HyZ5j9oBd5a0H1Gt8UJ+swGzHS6oRPIyupY8H508TB7SwlQyCuD5oRpI3W/b8cupX/
sNbu6gFOkTQiqhq8IVyVEZVhHuJESGQOSHHLN+sV6lnMhQEtcXqIdET8KjPYbiZGy5N7nR8M9vpB
WEoIck++0i6/oYVJ/nXzxRjfNT4f702wrBLfECjRqOaVtX0rPV/IvY6Ir/0jhx92+uO0OscEkI5l
hapuK2y6b+7DFnz+uXVQJ2+5X/CtDL0dssl8O101qrUwlCsdBam5okaijPpHRNXaFP65uzgcOhUG
agxxateiC/HA9qlXVKRNSTerxd0RFJ7xnE9TZ+kna0NDa4pnuA4YWZa7SrXPSFPAIoPbXIOGi0At
uqBeBsmgBWT/sON67rJplAQSszYa8/QixDSpjAF48O2jhoh83uC7zHlkquNfl7nOm9KrGdRP1a3L
iIlxfKYMiAQOkVPeHsjrCKWCjxdnMrXkRxDprUStIR3v46mGEe80jp1do0LDvQQ7+x6+lMR/oGCt
ZuhLwFI77OnxZDTjxL4qtaAriM17m+1mTreqzHHtOBdr55YpZKBQy1NcttKSBQkzkYm+0CuTVGNz
uReS+MkkYrDY/xu1zQ17RbCP0qlHF7qtqWSB9agyJMS+yCmJvLFl/Bd4yS0gsqghyxpZt2MAadus
YC26x54NC1qns5KlBQmCUZUTqHSVd0VK5AHGGQu8f+THbgofNQC+/ASUcDPNGztLgGwyPnPS+7iM
y16CFxda36ec7/blQ+KOlq8oBNoN1oM5cmql+O30rSWTiTjoWLMjNIFy73v2akrTkEdvw/HBtEB7
RFUJDzar/ig7MKpxhiAygqIrMnsWflsgh3pS0Ne3nmU0ZhltIzbHVEQxYbo/rCB7jafbJMKfVoZq
6ITcouYTxltHeD0pXbQaOShjfbnSSLIbh9144MbrZVFbYMUtMiRCOV1XbEYbvuC7b76sKEYBzWLm
iZbcVAXcimm3i57Aq8uAVn1twMRgty09OCg2qeXqtVQ6BU7qZBBQ43AxBX6khQXGNmx7Ny9Zf4+V
KiqkXcD6ySYSmxvcl495HOhkmoTSupbxn8+/m/QE7i6ykTXMk15ESIY4noj0J3MEWpaVu3rrV/Rs
RHhVAmiTrG7ZGFHjTwF+NnNa9nPHKUd0ekQhVzyQpkipeNMrVIcHKc2/mMLdL6jo4fh4egRHE829
Gc2HqY0+uRUdmiTsNR9CcipiPJeCtplxpiyKN0lGDPP8/5H/DBXcBw4vp91I1lpeTVmZ7iQ0O6ue
4ZIwR7JDWNI0LqKkbewrEAVHL7pw2VXLpqXbbpqRRJ5uc72LTBZ0+wR+OezZaJvQCnJO8buLOEB6
HjMeA8RqvrJz10Uvucqz/T1lCcvpMBeBUXgfR1HQUXmu+otNSYq7v+0g6euIQtM8CIWM4uhMSjxH
oLXvCG+Knb8IQxUezfQTAa87Ih5y6i0RVfZG8oQgkSf8Iy2Zc48WIQM8pjc2RiLoR3Yaq/8wqM6l
rnbz8nBUu0XcXLxwWPxEG4S4BM7TyowcnQzBhjDb+mGRprUWaHKr5/q+hMICMFNEpUUTnoJgCUTV
bEdUYFanvgts0pkFtQSJFTvjV4mddtNLPWHo2mOu2NLfetGC4PS3VLAacvnZ7PcjcMHV9yH2qMep
5Uc3DJHvFL+KNLLQfAWq83PHQszd5tGNCmpi5FDcdiMiUFsTCUY5xt37s3dHPhkGEgRX6gDIS5Ez
PJqYLk36TM5OLpNobwFOaB46DdShtMXFRiQ+yg1IwnTD9eti1vB8rNRqvqWMrDQGlOldxkGha2P4
xpjNAtlyFJGbAl+Zbzg+Pkh1UtTF/Y/aH+jCDbbbzB2Ea760LwvGDW2kb3yy0lo88klqYf87Z40d
tDgrNsfpfq/MNh+By4cDMXTsJMq6kAFahSm8helD1NWjCK+0qRlO9PqXMpFNJc0McBfDhxj/Ke4t
P/VG4x2A9ZCt7U/7/h56VRLfw18Ta3q31Saf590VbHdsqj2XogaVIfZTTsI7CWjkahIY8TUTwxkS
B73c/k6qtr+dkvniZLeFMz6Di8xQQiNH9eHSg8zEHFBIxFMMXZnIA4GiNbT+F5eS13OaNLgI1BBp
EVIjhPE49C41kZxyeYPALSDICJo2+oTIO4XHfGWWsD0OS6p3OTifbOGL83ycT5x7EuKr+q34sUJr
bgEj5kd3nakIdqkd5l4gi3uKrVKCtAIrvJkkXCwnXbKWpa+oP0NyRZ/5oCOeWi64SD+3M4cryEa5
sefzrene/ocOmDCBojH+jsWu5BOf2FFQIWLqm9dmj0M3tOnuhnBHuIP0Qgvi67V/fpWkF+m4ixtf
XogO7x+aqKwUEBNHWihHLbfyO+FAbNB86bsNcvb0qh91eHYiY2xAvnObGWm7xZp1IzNpmtZUQWU5
SltsrgtOVSk0gCSra9RYB3M2dTN7FXfLxZ2HgzVpB4LIk0BpwYBiGIRGqNRnv7h5At3o+LnUlFM/
ogwSZrNatyHLUF1UcWEBvm9MQon/MoReiFVXdUx4/PbJgFB4nj0WlECQ4y7krLC4B3x/WQfIu8RS
JRMAn8Jz5DoX3ls/NWY7O2v/vxG7FlQo86xuCO/BrMhdQB0QqB3fuZN74H+AL6HtZhS2Sxq0BHpy
k+IKzza8a/vBbEa+/Wz5WnHL0ttEVAoFZijZ45qTUB4KSHNFnI1V6ydxd9ZKyzGVqqzlmIBltHIL
UJlraiGr5XhLku6EnFk1Beod0BSCjog8DDzhtd2ydOd6ufSlPFqOOovEUbVJZkBJ7zAwnT5nm/nx
vYBwcLO4qjjM2IE6BEtOOr967UhlYbynflb5geci6qloDYIFnu9EClmPWMLSHWViukgznxWAXvsQ
NWxCCEyJ5m5q2tyso6KEWHULoUmJ+6+/rHW855owAYO59d8brUgHVCOd7JVptM6PRRQoFXaSTUWL
GkNEFV9IAJ1FJNZqs+DnF/W72EvwG5/aq7D6gf6b4fco43o6i7MzN+jdUx+p7KvtR+iab5VUre5y
c5B/vD6L/R6T1DQYSkSi1ytZfVU21RUZW6CRruuhEKj6ekDBxeLYCY7qgd8Ppc1UbXIcNa5JtawI
MDSkJTck7+GaRSQhCE7Uqxj/Wod8+GlrgtmEiz+U1JH+lZR+IC/Olm3RpY2UFhtRdhKs67vnsKlR
JcrRYo4PPUCJmw7YkFbZohfQEoVysLl60rSCdhJcGHtxJbRhiNSmb2tT24vhjwStKFWtat2Ibl1n
xsWilWktlrEXD1mp4aQMM+1b44fKEsCHm/mmcWzzJ+2Xj8Zy8bHOQTRdVxpal932huN8TmTBGM37
08QwCT6xgTq1AkphaN4WgzQcFGMAtrIPCYWiHlZWn/NFA+Bh4IlM2BcJyyZSNEOpzKT/ca7jmWsL
XEz4cKR91W1xdQZqQDYgSMvAvWN2aB8iMoywNiIQoi41ypW85UQHF8QyXGwPTU1iOcIXbMXmnrbk
+8EaHq1jAZG8EZueR/dSbDr3idj/8VNMBDKONppxKrBRfhIRHgelMhD8qkepKKTXs4wV7oKuUKtS
pPk++04pX5xFUANJ7o5PcSpq4TlpTiJlGazr8aY1l5VAFenvYgIkYheNiE04rmeDZqwYNwcGCb75
Ttg92aAhXrb19YlaqaeYw1jFXgvHDeJIy5nHyihpU9GE3WhCMqLI35wC32r52nAfq5ntpm3hwXmx
tuFgmJAIxyJ1YvxDqP6jOakdFOsuYz5pucHqGqCeZ6+PzQJ/Bjv9BXRVL+0yvbDWsqwCuStDQL5L
Or9hM+qasJDt2C8TOdJbrktP6uCTWkPEfjtyjon0w8CZfYgOjrXj/IZKBrrN+R4iWXNJ3ZhOARsn
ronNih8iuewKG8aWRRIwaCUiLMBczyDCavjWS9CSI90siE9zmJUiMwriVF4MsjNrvRh4CTp/xYv0
Z5eLtbXFuUwD4/qvRw7e+UFvuidF/NqV9P1xkecn6ga32aVoaqTUJ7JbPvrHog2yVtq7xovIRtVB
Ha7S1OJ5SsVBdAH3MAe5Oqao9NecGDpL5Zv7NhUHg3LNdcV4F+tDNZ4pAih91jCBliUJjW4f/wbZ
ej7HPslB8kD1++UbcnOoL+V6q/Et7jPeUDbvmcjTStXNBSUbTPPo6lBEPkPhHMAhVW8A7P4r0S6u
1LEgwCY5c19rUM8lqNU1VjPMTMTPMcvA15NA1UQNVBD4NCuLXhCV1JyTBSELb2URL1mkjIGbrTY4
8LXOfhSDuRAdX6PjYWPep/yHD2mf9VA1ejrsydnCAmRg0gKWL5bvKRCaUt8+nuoSBafs1C0cONEa
Gw/2gM3lhw1XlGnGJYBVGGjmosxfiwYSbJ/13yym8vXJmXxX/2218lzAVU2RAeIxbBewuoQ5c6L1
sKBYpapuZLYv7LyogxNChRC+pOWU8OuK4bA1QhinSVEFieLiR60gvxnA8nKlrgWemVfYXr+DDTIl
2k9BDLTzNyoqZl1IK3dmEvBiH1YK84xqo1GbiJcnxabMNfJuRITwdTi1Wa9u+UHTWxJrUtKwLJuX
q8b8ZWWCB7sy+VI8f4VGWsXUf4zhTRJyPPIUoBTSszl7CVKhUtaDYYx+yoho5O1OTNYW6wAwlvp1
wt5n2SHy5H3OUkU5wcxk4UfJMAM9+Ujl3+aJ3XDn+pAaVKs2/OZNQrDcJGnLUgLsCbCgnU0G/Njk
jAXAolss9JBu9Q2aWOJU0q/3FC3utV8ClJSbZI5r7IugphG3NQm08o7e9SsEcCYJMJONgYYUUlM4
xTcu5Y3Vajj3GpT1tuPaIQb1q1g848nPVs5VWDLkgsIU/Rt5SamSAXHWHPSY1Kqv2Jjkcuq8WWnB
ux6btXgT1qgup63d0u6jaIpfSLeNEFUm6mIr413HX3IcGYe/0LraADxZudc2f/VoJbxmktBNllnk
5/M3s7Q6Q2amcCF4BUnlHEUU5S/mA5VMelXTR0Rk8dcpcg1AB4rmg2/xfhZFx7YuVscfSHhBR3Vn
waK5MqjVG6I//Nq5WOnOijp3716gE+RgXUIAqdW533HyE6TfUyjTj9Sk8NJYjVr9LmX1N5HJUNTC
P8V73eqan61NFpvyXWJPxMT8gJU5joj88KwREZ2fc1p8AqUDjemITnLsMT2s3jeXldA6VZUgLgZL
uuR/YlUX12ScQuUHunlmPllIc7kVXl7dy7+rGVXyD5u8lSRSidgYopnj97k/lAA0+E0MTiIwgCMe
lFMq51j8JU6Qq8O1UWwN3CH6fCHdAkyvROrUNfvIvtmVyXYNCWl7dKKPRbuG+sNQzm1sRu5U6UFK
VK1vnUE/POg6sBxKpW7N7AL503Y0CaCnkktum5b+H82TzW8eP9gy4TGmNzdsua7XyQYYxYAdkH15
lmY5KO+Zn811gNclIDhFDEOmaHvVe2PTULEfnKpuT4PGAvyc4eX/bJZ6qnZh3sv21kz+DpPLTngE
tRevnJnddwJHNyvxz3oBMpSsm4BDfZpFyzY3IOBxybNRQSKIBIp+VLr5DRTAaTHBxV6URP3ulY9M
LDN/b4i/15n6W2sS7KvbCCHwWmvc3tr67sg3vahh2DDFGfvtv+3RDRjITuDI0BD7jwMJSYNpEfWv
KoX+7jczOz2bYWS1hB1QMdvfGYSGCGbYfms/N+I9LxYsVnHeiAwIASGNuS9qfW1H5EScoWAQJvfN
JSvPWmX/YoFOwk2O8YJ8ApPbjiql0BLE1JtL4KCYts5O0C7PLbMDZX1qFJiuxQpLLFyS45TDgz2I
M/kFo1FFWLmtuXKtoqKonO+DwnVD7KPANIPnaK7H5NHbOon7C2K4ixRafIJH75vLs10kw5tWm4K0
3uwxXGg+cAWczhFuB+GYYG1NolyvqGe0znULSzCO7mi+l9hCVAvMh4TrSjBE6nURbqB+6V6nyTjk
gdHobetDXE8EQhG9tbQ0AJ6DuHtmBLl0TtzyEahfxNnXMFSahLwelNDvOgIT6OYkCPjQY47qMbF1
cf9g7TdnGf1zHOFi5KYM/OwlTVHAylFSvBTuqUhP03TW7OXIsjoqd5wyOeHSTg0fXXa6gFdlkz5M
f163P1gu/nJVTnaJdftMKkWqRZhI4IA4BlgyLWPh/U2Yj6RMpbS6Os46pJXBNJqXUKiPlZb2V0C8
X5Pm+SN79wPWuVDUwAlbpNgr8D9s9t+abQiP2QfxfMnqThfP4PHufHkzsJzSXfWAuxZwVBbBiSoV
2wmTngieo0650Kn0KiFCrtNxChQnqfyCjy4BQaB3k9J+G9/lFjmI2vmJrhgg9MnZQRh5Upm+z1NM
4hJx7GXnwBLK8wm/m1qE1+8deUKU8iy/+e5O5A/hIhy1yPXWGNjvskcf8g507eUp4K581FEGksNu
d9AG8pB2NMnz3v+mcZBGSe2fqHY3ihe686c5cTxcJ26DjHff8mAzfgxxNkGZ5FT60uVdz8rRgNtW
arAnOORX3LZkLYDuDSE6R1sV/UANNo7cypNrJKASOp04bfWBduT+FznP38vgMOgK4obA9/XBnZ7W
TX9dMwlhdO9Fp3KDi45k2LxjNVmvsLEYhLKB2zhtqtqkDxk6tJhMTsRs65cz7sh2fXgIySj67T+c
1HEXC9Idiu+Y/v6vIFt36adbiD1iCNEhhxo9+YrPYEMC4FNYY+YLHpSxDa0mok9dAPeW6j7gRwxW
+LI/7dvOlHnCqHLIiJr6nBp0rFco75qfKzqyquKtrycyIRnCBOTPBFbxw9eGw4+mznTfGgxUgKhu
YnWPp2cCs8Jws3AIdX/JtVF6YDkSTxKPG7ByX7WiCL1TBfSxEtyFBSdVS1NuNLlZLOZq1pRiZAYb
TiHMyEmCKkY8FgX7yvKPg6DopHCC5nF3S4D6OalmY6VUtPsOo6G58MKCqSfTMG7iN4ms17MdtT9y
JA04oZtAdg0sFeLxniuKKeTbsPcWtLELvVP/XbNpyQqo6EQF/QTtoOVw6+5qv6ru6RucOr4+IPIS
90btEw1nvsB5r2ksBbBsZvnotVlfqpsQqdAKHLW5NbypEbXbzcYE/BM0yPxTlIJ9/xcWb9kePFTU
kSb8gurQImvCwEfX79WHVmjQCLDEsOg9oMSOYEmz+wR7bDWKq2hWSzS+L1ubJcR17mjTpnR+Rwpi
ZIX8LZqfk9aTSuVuWvlSjBn63mg7G7w1ZR/xEfPChAlASvwD4ng7y7TKdpAnXqTBbL/KCFB9dL5d
7+e0PQaf+mtKLqsb7m5npGgJqp2SgtvL783g/aGciRTczQ0GGBRJPr/DzclJVa2h27EWpX2LZMuR
/pFbfiL/qnL94Tdp3XZssC1cxoBrthaltRa3lY8/vYZYDfW6SyghWWWm7WgKZt/HDQyaJD5wrXlY
ovUT56NIZr+E3QpdTBSrJ1MAeP6sj9FNkOHmeYeRbrVp18M+QpGLwrcwiY4NceVLF+rRMTJyb0Xw
jbbTSpTYuvs4K6Ng6kzkfLrkoGhRysB/hf/7dxxyBcBvl0UWSqMi6ZSmrDRCcv5tlzHaAKfJHmgd
80jCFjf661iXTLaLC3Lkdal8dhrAJjzTnkV2JH8R3HIBn0KNPSNiH1m+7YkR8x2EnjopDI33ojCr
uXBPm9My6RDzr0HifnHt6CVDN9LECPjTk53j9njwIDxZEQe3rcy+iKDBKm7WhGuiWcINq33AX3Lf
WdKDkdo85JlLIDyuE2Pi54vVd5l3o19y8ji0pzJPYHXr1R0Z4fMhOx1XbhLzslJMYC/nsnf93Ze8
LGRk+H6ze5u8JbFgrGeIzR+p45/Z485bHt+WQ+3rvhKxmnhG6citqEmiir4tzSac1VhOfR4higb3
JPrkDIjQMBeUFtaznzec7qiEu2uFdAIakSgcc3zhR1IoVlwtmEbVgIeR2oUPgPqcni8m8lT9dXs3
46fvCVUqsp/yuW5oyIst3CCB2+Ns0LFQFuLqzWANCtqQulFNsj1AlWC1tozF+2+Z2i6h9c9ohbKf
VFA+6lUm5kLE1HXNo0qRuRjYUPIoHyl+DX9iuVTIx16LtFX2dX8hI6dFzGn8qvysPQO/yjFXcsUa
BJdau1oCJuMBJzVmHIVvjnBNOMSRAsi8gW3zrYb2RwlpWjfO/8LCGEAQhKi7s0IAhebG9Nf6l+Vf
RMyD43lQQe30MoIW9TU4p8dLJyuuEKI4AB8GALbLZqMCAl8+EAcS81RTilsSfUeziRQaqWTBE3c/
4pPa/IKsoKOfIOsVMO/aA5QQPjonmMLVl17L4p5SOAEttFZQEy5ZyrMoeh6qX5e7PF92x0P7c3t9
8A7IkvxYRCI0uWKFRlVNI9xVDNA6KGRAB0UEubiJMrxSGs8Um5Ct4HbmXZJhAN9IHCse2rXX4Pg9
C7C+2AsvDhYLO1YHG38j3pdrOKR8559X0237a/+RqzXDYuhKsyc0ni4BVTZ04UVUuTqBnOSRccdZ
WPqXkFDWJNr1mPQcueg1DAo8h1LeIW4l5j3i3AHvX/QytjV4uyZoc41OWJObZocdwfVPXmH5Cxnb
9kujvDmtGoD8uo83INDScnN7l+UQIIwsnpHOLZKptv/1FJIY/bgtObQoctEHo1GCJhTfmnfa8nmu
KVoMFeK0LwnfszsncL5A5dNzYYkmcM9Eo5g326JR98QxNbWcJdAjqampxY/ReEq0Nko6UvXOSv/m
0ktjO+Y6i/DGjEp/49uWtfI/noryP24w+wuKQGht6WZZgT/t0vGKmywQlAjxxqMhB1lfpR1tN1nt
hKUuyOBXlZAx/wLKuvlwQT2Wi8k1ff45pKmsd8CihZvpxnDV9PIH2+lgzwuFGVoVUwRsZgdODR8a
ZyXfW8lcObJ0KLIlxlOvTHd1vwd14S9NszqdGsIdj4Sc/C1TqIO9zkrCgVS9nG9gR8daike82H7p
rTCowdIgXkTR1ko/HSOdp6XIYP1Wg/t9nsCpDWthiAfiUcl9uIWrs+LhbZj5j7PTDEt/UnXAWpl2
mt7PgtPABDI/seumpBHv6Nfdnt795ixtvalJf7T+bw9sNyqFBTO0kpXzNtng4gQHAA3bgSwLvavo
k1xP3/zWM84hoOp4zgOsOZyN4jwD4yrDDawBClD5QE8JlbLOpO5QmHmeYHYmDGUj6tFKb/+44vzD
aimayO7rp5qTKeefEP+nQ70fCBBIDX8HpkOwQxgq98tmSU+F9E1kfT8XcmZedrBbI6YcGNNd69dW
mC/Y+WgVaHXAi8bbTsEnW0dVoJphj5RIcyXYHla0J+lqZQNmSutEQ572Xi1HCuiT8UjQKGBwcXs5
C1PXCEIe53hx30/Fra9aWZk8nvfA91J+G8Xjct6wCM7tluatNavjcYgRuLVnbhAwlO5q23fg36XN
Di5z5anSGrgbf3ixOQtXMi1yy9LioC3hycyhuvJCOWp9CH2OrQYqq6UjtrrP18GNjM7zAXmQLWGo
gRqk4Wutgq10nDnds6Hp4yJHI8HI/g/uCmNh71H26tZrcZum8vwZkkGAUCTw5y3NCaysDY/PYPhL
/MCml9Nn1yeIPg0dB679N+ep/VqlYwUAcyGCkfji2lr1os+dSFZF5soVQYE+cs2rPcyHQC0jbVYm
d3IupM0tTk7nok4maieoQx39MK+wn3tcS/ICHxxhGrGEXvPoQq3yJjBN/2WuoZR+IM/082wN/pn/
LetJwC6DKm3aclLcTWgoohEOMOTDmz8K0LAzpswjgHDsZB4uqheAJ7g+JeOQx9ETgvmY4KEcVWdp
Duxp4nNtfPY/WFIz7Bn7ElIikAp6pzRzxLyqydIosBM2O214oXnkaGYA8ohPetjBf/ED3xhLTcOO
X9jdf79qAEQWWrgsxlmUrOk72YAmiEPMCqXwEfxRWRxQiQSLFWpgYZLl/yspO0XY8jmuAZLZ3/G4
jMv4JLC0HRfOXnA+9B5YCMOYvKGlt1waj9v+sU3BaoJvuvZj1aiU0h5n5ynHWEq9rQotHBEUp5Fe
gJrMSk5MGoZ2Fk9FO/eotpeMQKW099rLkY8c3H0F0f9YEN7lbJRHHYabqmROIaXzHBLVZ7L87l5F
YYEHEbJyJ8k0ji3zP8LbTr5bsSMdn7YLwiHiSyhF0u8oe+c9R+3dVfEDQUU62cROUNSDUR8ICf0u
yPxwTiamtTQct93CgaVTxIM1uHNcyUC9Fon4AqLgXtCMhjDVMIQgnUWHFXHS1eUYZ8Ojs+mseZnV
2JS6J0MwsI6oqeQ7w3G13ftyy9s4Dl7OoVvuKxrH+1Vtx9hdp6rM5+8t/QrzAJCJfpBPo64GZnq4
qqzha0qWFoPUsQ67rXnX4jOHJyqxrXMDpxOWJQ4wsclZPkuGnKXceQe0g8YAnynUeyLJLo3rjBYa
A8Msccy/deitxjC9mTweGJjA0ZIyTxVsnw+Tzz78VavK3e5KeQbI5TvW/YFeom+wygUFHkqMMEry
imht1tY3QpUsT2wYcmJtVhVXtbxLB8EuIsUR3zTpnBsoOP9Y1ODg6TYj/mTf2HVhTEZu5zb4p28n
JHtj4mQeFLP80vQ1CnOXNQlWvr+szHBZ2qLM4ITCET8eeIXQSN6BumvXS/8EY1nB4J1Bl4aOfUec
5lCfswM0Scv3tLHPUgVIFKcHFqCGgzQnfsNjQ54xlVozdGTKYhHJVRi9K/eCi0vUE8qcP86mvnyP
IO8FfqUvHKHY4+8via3LJojluChu45SE6rPDljm36jJswLSLCPYcQs8BQ/CNQNsqGmEXKnZ+U9Iy
gtyzMeVypJUssVM0XMsk/Z8NECIvL/CmbdceM/O+I3kmL0bGJuHTWxRaBz+U5TXIWAFbpP3GRaJl
Gz6MTptTIPRJ0tsy2XghndjOheQAOhgAej/f4e/bBbQ4jOftHc6br7TKsTz58Bb26CgkH2CtMpSK
y+1E80bY4mrHLRvpLxQJRRqRp/hUa3hxUIr0ouV++F7/2ja7pXL1AghoUJy8Sqgydq3mhkgu0tXv
mrk1Aas4lRsVusM0gQMrRgQ7alnBkeTSO/04g/SY2VzmgH2ZHUT5s8klTnE1EDFJUMkRdxbnDhK3
p4awSNPtBCVkHHn2t1qYRjchp6O4BTrqd9BCaO2so+fyUaotSjsYe0zsAazFyJMbEIjvIgm+p+T2
EtRmT8o6ZIkf77uKfbisUYu3FSG70hJHuBzVado8EYA9pFHP8kqPYIsGMzUxTchjEaSo844zTtXR
Uu79rBgG51IC7U8byZNlFTirhZ27JKlty5tn5nyJafvg0oFbGIpRO8C3dviS6B/V/dU/Jjbj2Hm1
g7ZmPKLkxOxtTrQ73W9kbPiJPjICOF/y4UqKBFQnised7t+rppkNIxGKPhKCn7kE4KOwI/1biAnR
e99BDjoKTtBJbOUnmrJfZBMb03oxSdXYUjlO3ir1y7p8ZXHlDByF/YjXk6eDtFHjk0007jqiSmeb
eUWdPXnMFKuDZf1KALB1CbwhEMuFEZJOKBamD9S9s1N3mF+KLW5bLxUC0OG5uWfIYk6nsaGZrySr
WqAv5vAydp3M3rcNeMPAOOSZqjzPWGbe9D+7zlcmPl270YrYu4VSXYattVX4rkYRkllzVyNG02j4
cx2mislf+7hy8KoE8tZoTo9MF9bhxeaapG0L/h+/b/KIG01Y6XsWK23ZPRBHAIDB8m9eyp6QNZYf
gqrnVjynPKrdH2krG9KfkgIeZXkV0iQJqcI1ZEw4IaQN7oZ1o3y8Yy7kJWmkyu4pnElrvP5tod1G
8d6Nxd9cKrTD6XE4ERC9S4AjCkKFxfQZeJZHofEWFvBGTKthQ1XOAHUBFcgtHLPP4yz61zVIbWsF
xpJv8uqW94L5j4F5W8EYIvHOIvCUN1yAdiLFUpOs9KdNmzTaXLCKmqJDLiYnt4bWhzcBdb8mMwmv
186HbWVoqXchv+GL1bAI0k7lbPncn4OPGX5vnHEzDIfObWVNFjdxt72rWhZmuuXy+1zkzl6a7bT2
J5ZXBQXc8lU1aVuL5rGd+PYFe3QTrDJB8gNZa6+i9srBpH70Vog2lK4rRJzXCa3aEoxeaeLzBvsF
7YI/RlwKK3qQQtkjUzbw9oMBEO9uaPex8yrlMpysfTQktsw5OAi86GUfQAT6t83vECobtnN3f0LG
TT5Js8sujKZSLZMmkx2Vh9BWOEpD52F2bpv979R147xBcdwC8HcIHtG5SsfrOngqIPyaD8IHxJaq
aCAxyXsr+GTsWG1euPk42ebUtNChs92WwqpK73Myeo8ene1eBQlgivT8gOwPseBMXYNz40bVi2rN
GaV81XZ2pmpmEjG2Xdd+ddm4q4s3X97MJoGGJBbhItItQLms36G7/EZbTq3t0QY8wSwXwx2w26tp
1RlwF29uVkBvR8FB31zL21UThL1v4h2UIoX45ce4lKmQJSHN4RTKqG5fxIeiXn3z529ekz9Fx4Qw
ZTnq1KJncwYmv+dlWCXaMreWQJFM2sbTvbQ0ZpKrZF0KmUlopel/kapN9BQYZ6DihUR8fmueFOuW
mZM+WVVtCxxJau9KGQGSP43hrjKMv0gexxwpzeb4w7wy2t6+lNZEL6P8ii4he//8XsSNmpO+ibnl
GeJcyzt2qgtrFfL0wEqzPl2/TFpu929SdN20KKbO8eiNit75hFqR2PRmNwrK6A/x6+Xs1VjKA2qf
WkeSeLXLrsPXCKVxZECNYwa9gFVEpS8QrB+K6KArhEcI69JEdy+KpjufO11B4HD3JC8N3oVB2vPW
tr/cBXqlYyW06nh9GHh+Ea6bdaZHCrNSpZoeytOfmHjgrDXdtlRDaSZ38s9pa7u+HQ/cKVM77JNV
JAnHUCXnB+G7FVbqQnkjz6tS1NtFpPity4bK5NRB8xVmtWBMRG/oF8ZQl8mnb/S0xX+0RMoC2PQe
vUYJmDUAWce724EXtAx3poHKt34eawz+Ebeuyt71rY04oGcPILrVCk0mAQ2fKVy9Agmv8WYDOoWV
agaJiQtYwaN+G30QQc1LFMOsYOwzP2fDkusbcfJTdUjvxYegwzCswN8L4NZB83BrDTQf9Himwj/V
pKYHCgxi5ObfiiJNY6RmP0qTuiod3dwXG+eIPl1kFrlqVXGdAEcD35bNF+09MmEmto4M4Hd92+5E
c1uIf5LiDEoZBv7R93oXwx1eaZWT4m9obSXDS4YdaDypj1JZgn6vCOQvTlPoW+mmsrE7MhMXGkbS
JEtyKEkP/zkbw0xZ+2IZR8/oIkew8dMonyLA87JyOT41P+Qt/awIXaAfaG8cM9RErA7gH0e1hgah
gEC1vLEdu5ePop6VXRo56BFo8Y/Ba+GHGXjAY9lM7rFScfnDyzHkKsavQ7iWorVC6b2TR9a/6m8f
lAa/vfP7zClOEzhcXkocfpS6VX4seLEKgPt05zvTXjQZDNyTEpEBi+9t1ZXamUyxr76zllHSznR9
dfi8Ly6wMG71IGArbdpgjPccn4lsZ2lA3V/ygmUm1YxwX3I//cOaL+0Fldcs1QZlOkP6N0kC1q/O
I6uqpFCqC3EsG70vxUCw++MTa7VhjkBgHa3OFrLwVWjLlxjOGzXSIg23yUFC72mHVjx63BHLL7+d
fa2QKyO0Orhn+ikdiqjGppMdNQkFIjzIeHIct2eIQMqfaYcNEVEzjHl6v48WsBJGn9AMQ4hQf8yV
vpsJaN0FLvOoT9koepcLZfYbqLMK/S+vO+DtEfIQRG89mAGAidbnB0StRv7PtksH1PaHW1bmDWbf
7H3Reo7CFEUzTJEzoMm2kRiVg9lAIERDuyhq9VaYlj+joulxS3QZhjVgovtDqtM3onskEHs4I9kY
Qfju05yLLSgWWaIputIIVXy1cpOnfE617j6w+vbC65GsOLTlKR7Tk/PLzi6EnFaMeHK5WpN9Lb+b
jxAoLPCYJ1LqhOeinIlyQJpLya/0K2bYmacndEtNnIdmXN2IcnG8rXgsO/jP9qCCHRDoOuh0lslH
dfmxcy4QENGceN23hbvxZgNJcyzd4PysvJc2VVDmaiVFIB27XHhvjX0wd0NmZAE2AW1RHCe04aHz
zltZdOlfD8qds/1TI6K+SMrt2Q2T7U3JG0RuTEHltPr7ZiM214vZMSoxw/42pymOUaRLVvVYw7Zd
0+EeY+pBQPPqbmISqge9ZYWNBkkOUMNmgvW/nJFbzkfMCmQNidZB2v+xCA0W1AYS7ZBXTW4jBp1z
gUv530KxJWrHAjrrCIs85aRM7q9qc736T/OqKHDuLlRtHiqNsJYYOTmyiTIgkZ8wibhG19UyK2aG
VJfC7m8JUTZQatfXReQqVd1Ja2a/+23+3vzhQTQxif2HfmO9zEfNHASMnfeRXQKnvaY5dTYYLZ/E
IMk1tnoo+NMHcDxJXjutrZa6s0AzUcBnWpTF/dpiOadTiDPMH2FGP3HdrhkAyNT1s/XuvmsyPthC
paAmtjJpadPHpsNU8FtD0xpWRLV4j5F5UhjX6kJgACD3H/SvriNAChyNwOfPmH59/4z2SUMpOyEa
3zt8w9V8GnDw7wL/6HTvwahSuAReavJbfc94mpTbPDI65SX6CvDN/QS8AjlCJSSoWIV8zI+snOeW
EsM08+xvA4ArrI/0XIGkEaEdn70gHtS+65ktDErnwWGLtg7wqIosdo91yTRU2yMe+f6p9SG1D9yH
Ko5m0FJJln1VY1UhvFMvb+aKYCobF4Ug0q5fAfKxZVju8idB6EinoFF2/WMXkfRVU+W3HSMNLu2N
I1DiBnYeky77vQjlhzcluWhGnDkJRhTj6+mo3YOmSBXD8LnKbcZkMevxRBY5tDWtnf/xXn1lh31t
ZjnS+tVokyylX+WEc++IWhqsYXi7azYT3bWR3W40z/iN49tx60eiFSRGoywvw+k+E2Mi4l55DKIU
QXIE75ZJZQBKvcKi8df/Nafx4enKhX/z/0lmZhGxxIIeAMXGyNmxmoR6BzQPNrmbWlb/mLO9Xl5s
F/ogv5YwAG2MtNcF0oroDwUg+voQMkmBvKuDwkeesup50SspYwzK76MQ9adtCRBYKqwQtvyucHXK
vZ3dfLOloMvmYdYjL36Ep4btGgV3FZRAeiuV9yTUOyKTCyzIlV0xNbsJune2hRtF2Ba6KSITwjHi
sBPiYREovdlKRKdbvBL1KPlC1WOMNZGjfn8lmyu2HlXyrbGtDj8AWoFhn9WSctOuIjEw5JUakTtj
fILVOoIXXq5qhp5fYV2iMVnCLPSIhT/UjqQvejIqBXoudmqZJwbcsmUnZIHA7QGc0aiwez5AjOYg
TaK3aCFFiblUddm1Fjmxue+GoNIAwSXvqMfM2vU+Uows53agtscAQj70zB1vJbqUw17C6d9IXPTT
PCCoMqBoCxfhaMgZKJI7pRtOBnC+nN80TNzF7sJJQ6kCwsZ7ogKswN5ihZJv8cqpC0KqnFVS4aSg
B3e05a4vlW1/CBYgovW54Jmjj//HczptfUA+FDvpD/ZBbrqr1ob8OWiV7vDN2gFVG25C7R6FdGDR
Awiikg9MggZWFWcnq0jfRR+Xtw6D3/sKbO1VRqJOUlbGQLk+sN+Dz6t7o9ssq4tiOJV/6v1UAysl
K59GHYrl2PgTVOw+bOqGgzN6HrkZI/5U4QptM+vUhH8I93I2Pz3i9OYQptZ2L4wvSBFaA8yg1akv
5LzQvfYELkzerhJgLolZO0noMYGEGVOk64yWxnjXrQbWk0Aa0Bb8HnhNYW2byzYBLUy6i0X9JGb0
uRfelk02l0zyzTXIub52Y6tVeMPvKXgqhN9EwjKyg/GRAdzcziImOZ8unPElsxswCPeUxyKhTeGJ
B3CUDKzYRvjWT76YcxokYvz4UBXOnVyzC1K5eY3XMjmJ+60hKbm7LQYeXH+Ds83UbAQXX0l1v02a
wlRyuF765qM6Glq8GdODVbHS3ydvQlr7Dg5LaArxJDO+wlb8Sgl2DpISSwkK1dMCSFLpocigxKmT
Lt1jNjrnHAQilEdKkEBvmmzOV7P0WPaqQNX5FmhkFCgFqk/SjmAP/I2WrDOfaAw0qlV60wDnv1dL
cKvQlc1JN2KyIHibcbF0PRbY+jLPFGwvaYHYQlepNFFkLcPQqGqhPngLtEvZytfARb7sdpw7/Dyy
jzzIENPbJCLUF+wHqZ47OQfbGQwcBFF39L1dPDiXSYxTbOWUqhqIBngYynvwb+El22IGdkMSAT53
PFaYyKJ0+x1OAYD+P4UBiGT8BXKyIVCAg+GY9WsBIRb15wjTf/rNKKhcJM//GK19oV0/rjt4rUp/
+5PHuCIIgPoQonfTfiW6HNy0JA+3ehh6eB+aqGZx14v7xvyE+hDAOYMm4HA6itVelsW6h76P9VQY
BZa8Qy1W+cBMkMMsV4Q48BduUAciGNwX+9akwqWZXzcoS+su55SJu8m7/HpWT1fu2W40DKBIwOtl
WwkHBagW9F8RUCTTe9ieHxleDcn0aPMVrZim/ABI7B3yey7GQ3KXD9X2LWR0FSsXBcNZtYeQR72F
cf1kEIOW//WU2hY2aU5VYuE55+/uEx0y3vJklF2Zgxp01ZNrdfWN7zs3J4k4Fw1sVAQydzlTwW33
dg+Ec9IjFlmebNd0v87UXfmA6OVMgdj+pS37Nm3z7hLTfmmMfgqbXUGBSQBaHft9Tk+n7ReNeTRH
81XI8mgMR5//ButjNnKtqw1Y75LzhIc1rRTCjnEKhhkVqIBBqZDhwrh2WyHyygpKQGKbH65tFII7
lRfJ/O7lklpW7C/TfqdhtlWMjEBtwVF8zMIVzMACGW5knRfL+aCVD4Fsd8LlRtRi5YNRoGfx8SMS
Rl9EsMZRhN4qNoq909lnbHmryMaFOd2W34CSWa4/X9P9xghnyiO5aHNhM88CD2SZ4cD/oo7IBa/s
ieS2Chh3PHmmaKsFOH5xByfUs+Q53q7BFKgFjWwBoF/gT87Eu9PSUO6668nWO54+IE+ZoHbnIMCl
aiugF7mSU0x2P5BMBJW89WoZ9dECYD/FbpjYjuToV90bMT84DUI5DIwdW0UjPinR8FY6WIkEvu9q
O/0P47FRovyM6aC3RszmGnpHciIpsmKny4w39kxtlIE0IUJabTeB5t9NvwMTq1Fhs8ykMHrERrtU
2OBq67NsMfbBq849iKq+eWgK66eRVC7+bP7EB9daCanSe3/Nodv/RE+Q5UvUPT/XWvuVAZ3+Cx2i
+ntoZAGA375ZamiUrw1tq+0r/rUiM8nhw3B9GTF6rql/AaXE6qPQfHo7dNN8iAS5bRcn+ycGWHny
MnYE27gtM9EN6vEfGW1H/tbWZTxVR1l/I9B6WU8h0Us0LD7G5DIZSIIJZm79tD8N2KVybpDfxzvx
Md3cLgzdzRLvDMhOkQU15/vZAcveAdiQoWO9Jn2wCAQmno91kJnuMif2CNj1pXRuWGFSODV5wQAd
ZGJxKPLTNH434MU2+efgrShNLrAM7IRua3Su2cFG808w4OQ52NUoaPQvEumXDlskyK6xvOR6eNiS
DyigPdiqicjUHe+y/wnzdHiT0jRAQDadVTqHF7OIbu8IWK/irEAwDNVyMzMZzA9CDUPqZJrFn9oI
SXHOLxwP8B+X450PLsxa46nWIv2TgQtEHcy8nWg3MfkpPHAEsuYx0ab6C4y4GQ6vwhmyZ+Wst+NP
Rby7iociK0iCE1XKKWnIrGjx7A98nzZnNMUf8AYqY8H9yWlafsEfevBBmR3mpM6YGD8ZplrQv+pv
VTejMSKSAdLrAPOvHYzV4Uy7F0GYe9AyisWIB7Bzs6hr6jpeF3AyAT7X3FiGv0SqkePqwlvgC1eO
/tb9bJXO36X/bFJNI6O5Jhaws6ob/3BgqtZSFf01n7qK7BCOxuBBTRg9ojmAvq0GfjXCl2Rf5rvp
Ls3YnAeHHaURPJxDWGk54CTlsD+IG2YUckBpD5hdhwYf37LQQf3CORIqZYditBllacf8z8u/1H21
MwUihuHYPnBTr3GegyIEocVEcIx3gg80H+ecdpRvhSRF7+db0UP7txtY48KTItM0vfpatpWN77zP
jPNrKLwJuPpuzFMcZlzEHWvfcVoonBQgcJclUEWryeiILQKRbOkTca8TpH9YS44RbiwEoDYa85/U
jawp4l97SoBcGTBgdmRP1GojyILu0gbufLS02Dd7iSxKwpI54wawBadoYO27saN4JnoYcP/TnoZc
VR1Phve09KIfbKu5p58FTwepNSdKDfLdxnbLpWEUwKHqfIBUOBXAYJtvOfTRKyGp25k1fXvxKuPJ
Wo1Xji3QGzYVLTCTwLK7uBGCPNlAozMVS2fMdfua4ZcvW2n4a2QfjpRd9DZrZAR5NTArHKLG7tAv
ZOKpVLurZY5AYwBw0tkbmkOpFjEtJcJgg6sIgkrWVqKcNGErDQKKgJccXC9sW9LupsFpO9uOGaLW
mvqKGiaoz7lu4CRirKRclMctrbY1XT0UYbBTmPxljURAcafBsA1noNutFcYmBP3a27otlX0DfZjS
JiVWpDzyAQK/QK/rva9iP5GC3sFn0tGGSUqJ67VYd/dO7pf393VFXcxP1na16TTqTEMmd2HBCCIC
sWJ6n1ez7i04B6DKZ/+Y1fbBffl/V93D++HlMLMIyWo9QbLHZR293yoc9aOAPYFo3ix2Bv3jDSE3
IPYT3uaoNRFHuLPyivzMKfO8TRNTlrcUG0DM2gIpMOh6tq7jn7uM/PrIDD7SB4ZvA0x5o/1wlI/G
Q8oE5AQZhBZnj+YoUd4z62KEx2ZgOGlDpr4p2AcefBLw63nHx0UCfHNoLvKBaLljDHQdq4UtV8wh
eqFRF0RjLAyqlIYpiwvJcATp45udtfCmBXt4/Y5CVozIJ7wo1vM4KqtEgCrpYhI2X2GosLXYLzSj
a3RbOPqflpuTPo84UpUjezsJw8HqI3Haislw1RI4C9JylFwQqJ4TvNt3YKysTczURtUh1MjTHPTg
kdMyEs8s+7goxL7k1nu4d6kK2CKO+AaWA3bafnsoVlhIjZN7eFrEOrktlGgLcFs+Mcy1/qeKg0pe
YwElQey7sXhW7NeD+16QxzJe2m4bJERFdsKQirNpzpR32k12kqEf5yeyGhjIxax6SDnzn0v4rLBK
uKAOjObghvCw3dpx1tzcGeu1aCVR1QyJ9rtFCAAh0zKEra6M34FUFdwyyAaJwK0BOHKZbHj+PdNN
az1dqJXBx7iruz9D926cmOn1+MfvPX39QGFzB5Sfk4/W0eAOcK6dKWXk7hM/i5I4b+rN2A0BEc19
Mx435/zfaP4CRqy7HPz4sH9VmllC8mWKkXqY/OcOiQYhERgLxbgCFKvhQsxvUCmmsXPrNColccao
OyAQt5DS2o/SkGvR35CNwnBBZUv8LseVUDUmCWkM3Fyba1dVR1BxrLlFx9B92/rg/26JX33ZIla5
SOQFySuf9uL1+G6eHoDzuFFwy8TR+hyJV6L+Ume4vuMPx3Bv47ojoqi2xLscgjed7WS1VZ/3NSRL
cRKTDeMbNj5wgZBPAauzvAO1m5PWznR0Et4GvIIPFr8vVdaV5DCSu8LpOshmD7oWHh4qJ5lEQdPQ
wkoGlNx7zbmpc4u6alMsM/rVvpAdyDZxcujFCGgbNkd+22r4/dyuyKA6wWDjDUFbddcTF0KM+yHi
P9VFK5nailjolwBSXY8BvfkWtKcKuVrssVdjUtCwAh0PthjOpIBsa/PZ05ynIHjtNs6rLKvqSU9z
mKFHA08t0EXB2vbDNFTuozTWdZ1fu9Ru2DAjipATWFoTWnT8qpA9o6aL7DL9bA2Qzh0RGewaGV75
np2utvYKWHC4WnbIaUWo94LWAEVcsCDGOnbHcslcsarAZdXO9mG7hIII5qa0k/Zk6rPqo6Vr65s0
ON7Xx+qBgkJicD9f/ZY3XAqx0VtDWbcvGjlf7PO+ah/iRVEGNWN8W1rIVmrXDaJ2AWUGo51XhsPb
IvE85oEl2OJqipnqvFctXUvletOrTVkLTaYPV0oul/iSGRxtBn+vOfr3fjE4bveSD77YIziEu2eK
7Z3CRWxIC6RsmOkHmOWYwGW+RjQxkGiX/MIIH60K72IFwxIqikIqmdcuy/9nzx4BOWEAvniZIcF0
cqgxN/exYLqvdGTJdOQFklbZz9cr5ki01DcqBgA7dPSjbD2er9bMxcDqr3G0oXdG0zZrnjyDQQFZ
jY/eBxW7tltRZf23QoW8iQ1Igi1kfrNkWn79/fiJR8xpaTg6RHG2eAr/eaePWYvHNDgCDZu6Ijv9
pGZgKUNFTCrY/u2xsMqAv5zFwp++TjoKHB073RczhcGA1waejQtcftECoVyjZZ6Nm1HD8vDn++8N
vGIc5LVzWIAl10/4+nEvlrXz/E4R6uFviYC5dgPCrgvpJeyCI3Ned5bpr48wXoTFpnsgTEyhO/oZ
QNTf9L1RQrdO2bLbliNhKTSL4jHuEUkOMLITY1miXJyhXLfhHShIqDpRmiwjptoFZ8DPZq0spozd
zxoIQU+JWYGIgLYzVZBY2+L2Oq8FykYtWf0fstYGXQSUa5fq1M03IufHXt71y4/dbjUFcPdJh3oN
39FcwwnPpQAXG8IXz1dUsCSt4H7/I6/C6/3THFYDXr+s8XYSGapNpoYZojh3EeF2O43XJCASaVTu
CkEPGLckvBHSe6kMNumJt4ryeU7UE8Yn3wEmRvxx21P7/k4PYcOT3uDLlwyXRGTNImLkBabLf4je
Sdf4ygXHnEVoOPEV2EPw+LQaifpnRx3kWOFrtlUOjg3OF/cekPkNHs/l21Mw8phdTuy0dXQiQrCL
Eav1i0Kno9lkez0o/VplbgQqQ3aNE/E/mOAML/9LAI7CtvIcM6cwfbNe1fhqkPzBDErHwTVbVByW
J62AZ/6AcnHYnhSgpiw9R/rKQ5eJRVo7BEgAj8h1K0Od0y5TzC2n0Dcwtoasq1up679432U8Hcd+
KKCW3vqF6OOOTJ+tUqYtQNZote/sqDMqvtjLqPv3LymhqP9ZZ8D3jRCc4Jhdn1HrT7IBFQJ5cGcC
FR+7UvoKx2ehbKO3mH1GYVFrrjSgquhFV9EupNVJGA579P4pSep7ltf7AGazOr2HP3ULoexHHkpQ
gwUBJGJqtu5ikMsKay+dncnkwjKcUn3oIZl69NWlFoPpKTXd5C2ON7AO/wVloC564dePpElbQpSk
dHGqHOUc5n3gD4Nc+x+SdJdWeiH9EQmneCohJGin0YyT8N0yHEcAIyiJlFxt9zIHdxPjnfqI5wUf
oZnc50Riedn9Koa7aG7yfGAkjjuDIykhlnOEgmQSVri0Mj+LWkNGWHkZ8DD3xDhbNbsTQeZxkl7F
aXRNb9LWyl1/mtyJUEK8wvsH/q5IvlOTvYhwyjAeTC/tcbxQaHbqCNFi8ZeaABCqcWGiUgB2vi0m
v2IpQ15Ve9zrXTYMzo34MQTOjd7BcR1A8bpQoZSFvd1+My+2hgjJoKXS6J6ZFa4kmPfYyY3cBoCe
1Xye5mtwmuJY5AnZtEKq6PRJHk3jn1z/rWvYAGzC2cT9V314225p+DO0GEVmO9bR50tYEYLX3WK0
sz5HXMYFY5Piu+Qsv08XL3CaUF1FNkWC4+pgtvGXZsaLBk04uBDRXjtw39rRiHQGaELymaUUBGDb
4KvJk5IkO4+n27FSI6QCYlZux1N4kBqM9DizhXobA2wVIcDHS4hgxM6vyzSVJgEI9T/Alzig+fW9
yeciK+i7U4Cl2e7iRavZqXZ3uJi0qxoS0oQoxcTSw0gyqJRjuv776QbnHT2DKvVG+o2iyzPZVeTL
MEbHaYUQ8OEy75pbr4HEKEZTaDPXuIlEnOH/YUTCdzaUlYeVOxOS2RPnnhmPavOWa3ELZs+v/m2I
YcAeA8lUzH2k8dNA7XSSXpzJzGGX4+7FkNSrXJmSNDFiBbBqxIWHdCKodp0urqr/B4XUpJRkTOES
RtuQZwgnhQQleJa+BTZnztLnNOQ9YWxS2qbLUDliDK42MnPCDpBSI54o/5YCM1APtR1Zku0s7qZ5
sWtdoRcy2de32ZrWBk3vqsXBmdiRWckVpCyWsknuoeX4G53mYS05/EzYn4FNz5/EfLwQfawKU56Y
fer8xvxwf8fPYIlaeN/Ni93LgMQOcccfwhnJ8odAoBSNj8BtU66YSOi0oL82HW9yD9TndtBtnzBE
6wm0BACYwFdJswq51V7SMmQbXmQnqpg/ZzvPfVGw3gAlhaW6lAcdAQd5j7JPiEIFB5k0+qzubCMY
eQCyBlDcFtNwVenqfL5byX6+1pQP07MZ8neaFJrAEv0dSi2pyd7+v+W1AvuKHI3w39draLxioc1A
rJrnaL6k4N/myAbs2g3vHhKAWkVAI5roVKXBDdzTQLzo4ihohG/zPVB6wcOzrV6n/pr3BNHsc7CN
pYtJu7bGyJZ+BcF3G5yK6WCn1LdkZ3EY1KidoUZy9Bpqd+tLNbkAgpDVc8GSNulBaAjUyZt/9rXZ
5/k6WgROobFSehPe5bNL+lMJwSxWxthFrizcUbrMoO//NKudHbg1MSXSRQx6cqB9r6s3J+x5PeFN
boBNGmA3Im8ogts8QSPE0paLWUKiY+KWOmntnHhNl2ef7AP1JtKTj1hwA4GFG/dW6SHl88ZB8yg3
e+yrPJ1LBcVE4tH0byOhAENFVm2P+ccnkGp2ZOqOZIzRiwyJqUcKxwNxsUYgt/Z9A06+wzIIe++o
hwc/GyhrT722O3co+Lbq7hGBKuqL8wB5J0/i+ltBrBvHk2vSqWlMh3qc+oJaw6VLf1GHj3eUp6TL
FMBt0D0Lp4JfmRzB9jfKBpdgb4VQVXjql3+XF3+UvYyIbp8S+nFZpTWbpE6Y0eQNGuFxtm6mHVHa
vRV4Jwij7pi5t6vjxf2Y8kXEN2BnBFu0CdcsE1wLJkXLy9vcqG11+YcLAsKgNqVrlwqqVINPuNsX
A9zE29FmlMcoHj7Drx0opwoGbOHYwV60E5z+TRYl0R0mCGnEdTN+gmxfxPpxxpA5eQRkq1dkMgJ5
pUl4/YMDbnKPFnHxmloQY1ioYrgjYJQKE0dv3wcwFbY8rkVt2bvzAu82jerJ/lVU3NMi8k5p1AeH
GecrDHGU63K7oF1GaPWlq0orlvt3Ywq3cGrU6t4scis7wM7xGt17hHVWksrBGeSI6l0+505URROP
jz9Dr85Bg+FvDg9jdH5xUSBWuws9oATMtCV37PZiaj4Oe4HgBmoaTNTFkbj2ZpmAT79xZZkIP8t9
fb6ztVGSjO/mZj4udGTOYAKEM5dwMEQW72aiLwAwxjAjL7We9tOAvb0DAQ+Nc9kSkQm3SA2Z0SV9
6GcxIo/qsVNiKJ+0eYJePc89dZjAb5PmGTr1zTaHNUiBtLA/FmNcqlBFH3WPEs3qMPQRR5GoNdG/
Kj3c3swAP7nODhl7LkfquPz0/v36Gq0nHfaUjA1qNSGlMHFm9xxR0sSvo+uAG5uhqLMrfaRXe8UL
vwfnwi6Y4QjaCEaQkuQKS2QjD0HDGm/YosTK7rM8rA8RwM2/FBWsukEixeIHMIT4S5Tk7kvPkoTP
RAOj7BwxWrenASdVM0xkF0m+VOR1yzvxxETleZbUDYG4zb4QfbVIXYjbwzASm5B8VjmVisPmUj1I
mrcUHvpIHW3Yuk49y3hIvb2F2u2oh85N6ZLUKlaYktshZuQJMTKz5WUJNejMUfWLF2CS0+tFNbIK
YDuhqIVZBRJEh0AUYIyCrHb4haBLLFSpjzOsxNHndzAo2Ae4xBeed6AV/iTAg5WYnBpdudGIBABD
ssrgwSkRswoS2GU1RoyZGdL4WKbmAXNHJaQ2hLJ6x4FW9kjMVlxacE2i8Fh3uaTb78HljmBfOSYa
JvizDScSHr9+lr3/uIcc7trzUoK7db/oDqGyFyzx2BkUoG406Cqv8y4pxjL+i/Wocnyq0II/IIYi
oC44E770CC8LtIBYJ1QR0E1jgMav/UdjfxNNr6liWy0qdIl2V/xgKhVV3aE7JpwiyWE4OtRBbsRf
a4ZoEVIlI99xB2sTG4Pwz8hUKaLlPHgcUXe4s/wogNn0nCmdNQh/DKV+5cbCUkUgBbjqDG7QZnc3
lQJgZ0NQH+0Y7fy6//C7Jp+6z22jT/WGTiA8VF1bx5u/KoSHaJdCI02sHM8tBvyLlOa5ijJXCoD2
XuUhHC7QMLQIk9uoC3xRB+yfQor8z6hJNhZl+g08RlyGiNGLcROtQk5/bi/j5e+C7uSlytSwLyAg
RfOwAomG7LSaMZ6R45d/g7JGAgoFEMII6RpYCSPm9JHdQ/D0gPXj24zf6OGpzrx/yOSraBjnxEL3
f+v9yVhoLPe8m59pqN9mYCpatOSXOPuOGVMEJqDo8qMor7hUDyS5un/csx0825TsBKECj8q7PLr/
Pywg6/SZFlOa0PskkYBuPkHIhoc/RvmGMj+XvC8n6RPhbfiY58sdhdOTvp6LeNecAxlOD3rWKjzK
bOaHXBq4wnIZwMrELg08d9hqTbfF1O1gNGeR4+ck7KUt1opC8OT8dVptoMq6YsYh0jpPuBf/T41E
2aeJq+Fhehq4Ij2/x8hZMYSDLRn2uzYa7/WejUUuvbSYcNerksSibS66gOS5YqpXZO2jdI8IIAbv
GoPQynNeIun/O3TaWCg/T4NJYZIvQoIFcnF/UDTVEpcx77Oy6faDzx7iyRgrTuWwUwBWpYvUWm/Z
+ZOGQZBxluGo4HukpFiNqqVYDJ6lRvPha+UPC0VJKsujyv9dVFDnXydAFF7UkePVgP+s1l7flbPL
XkoVaQtsKlzOx72tg9nDoSAlB2FDBk2DR4FMBnaFomlaGWWd6mykH13dEZAreJypVIQs2TO6d4AC
MJKV3QRDioc7Tm3qFlR1dtko8lpRa9FUJgj2sKLfUb6WLsUDc5ibGTqeLD+BYy0SWgDzbSIRVfwP
Cok4qr/IMYdv8N+TmB2KHNV2UbvONpTXh42+n7wp1rq6zxIjBU5p5gRP7Q+nRpEWQwRmawzF67Em
YgiQh0iRq3BexocUUYDFis3AopqOh12t3zd2Uyw5UEB+zW46SjW+YpvXek0DrDDQmK0CkJI/KYN6
4ixfSEgh0HPuOerj9kkuAnivxK1r47VU7AFFNsUIIs/t7XcooIqC/W/l7fsd7GI67RCOm2REiDs0
ZvY7lJ3a93Wj9hXntn/pWMDKHiyXM6szHrOQmSjm5ccpNW+5FwEBu4C6XUJcmbXqeRBi9H7qlYbf
8ZZPHI8DdTy5018Yji/tcB4NGDDlhGb647ED8P6mZf5Ui9pBxb/DDBNlEsBvZdEGEODf2768mtAK
gMsvF4MKf/VvPMQhQ9B/f82RcfLaq7qFD7GMMNG9kAzV8AQmBfziejeeNQsTuLhgsGaEPQLT9dW2
VlNDV0i7gEkXRqOIob4wdyuCbFovLHOGq9Z4CwLiMiyMFqwk3ax6/14yzjKcDa8D8sm2pfhZFGMT
mabk+bkhp4Rr/XAZcZrduFhD36wD9PquB0ozwSviDq//z1nMfcD31QRXXit4FOIt8KNOB4+K/tyz
1o2Gy8O0nhCLVdnHwXunXZeK8A86T2wWEDpfC2ABqsTAQwk62rvoJ41sFhMp7WYk91cZHAPDlwlA
V6JbC4vZ949aLTeZLXbEHmIHaQbZpV71T2Htp45kUdJ5K2/p4TpUUg8/dakjWpf6sNTW3SnQG98K
bY3imGtBuMRv2ZdJAUXyMh5A1mFyn/6S/RkNMMqjnBtRF4FQoZbqmog7xOqP+og+VpwZeWKjZEgG
CuUS7wfuW+pcPDONgSCUsGoBhaR/k5EVNi+A2o01iRDsHiu1T22Ga0SnvJJ6b831iSkL3MA1Qlg0
tQBIxzPjcZ4vSiLzm49Or3URSW16PUYKJpRA95P5gn3KJ/Ccrj++dD0mgvwrzkRMLt+SYQaJHZiR
a3wS2CMnBwPHTvJSP2D23dOSmVrj5LEC6ZG44T4e0foglkGP65iTDGA5GZHHH+WwuGyp4RziF7Dr
Bzyq6hitI8Fi9QFp5k6GgzUpmrr30zT1UNcdZVAH8jFn1QxjXYbqV8yHHF0oDXTShvolC/dRfNTg
GRTcx57ydSm2U14oCsnN+Q8GhIlETtSdyJWq4AcrHXjjvxaRiqouRMsfg8fzkq88g7Zd6N+lpErH
xG5PIREv4/N1kFeNCi/IrTCaoHMOafKpDz3pg1mP3sc8jyrm18sO/OhELIxlxwXZ5hU79euIXW/Y
P7H1MiXeoIUYCXtn0o5DzZ2IQCnXJ6HeRf1Vkt/izvxuOvHKcwQ/Wt6q1Dz+ksdsR4l4+3+LBntb
5o87qEHMnJ9zY0BD8l9mPPleUPVu8+kKpMjNMynulC7KFr1WG8uvYMo+0s/V33qrh/lztbGkjPTa
SipTEcDzwxzQvv1lAFQQC4qlX/TvPVYDCqIHjeJLdzWDThEHH4ZKMiVMcigTGrScKVF+4MepIg58
hlSB0M2b+tHPbqThSPSTyUY9gIi3CWahBzH1v8RA+hEU3aFAvS2jxBjMQKzXIFZ0Ub/eXtN/3Y/p
qTgUB8gJRXzQivR4aHmGfHUX73ztjMVM8Dc3PVfpUG/SQklwtXFcEFuxpAltjnB3u1RWX3psTqpm
h+q+RsYBg5pNjjW4aPEeCRLfX3seGv4nrnO21j+EbU2gKYQp1N/RDIDaiLwvNWTh5OFRj/SmV99P
d7QlGHcnDXGy2rwxFjqKNeoYK7eOaR+jKREIdryzH7bASdCEMRG45i6Ujd5m7GJkA5XblVW5IQPq
s3UgTCAlgBuQURiy+y6OYlWAX3wYm/xa/PR/VB/3pDxbhf9qoLBbMkwL/qk1edAAz4WUgEIRLRqJ
wTUfE1HSHX77ls26jrYgNbNqAbxFvbJlqIkfAYZx+pIv1/cNQrrFBE6bmACYjqNpERhSYdsbRvaq
2w+tx16fSLIcyWLsA1sLkWZlEUqjTFPn+KB+gOeR1D75cZEwaZD7LhQwfTi9BrVxImh66mbjVbzm
RH78Fe+c+g1qE7+Rcz5JN4zALc2LF2qpn4MLctJ+jPOzIOaZfO1Ffj15sGLZCA5Igvvs8TZs36Y1
2DnwjcW+cW8QV6vfXoKaEBBORvJZdsTxY7vv+DMJqhTaDgm3YZg7k3abQ16+qrKvWFW/cskFse9W
Ht/yol3cLOKhkH3rDNt6R7vB5FP2sfzxh/TVy8rAsCRBJnf6hK80idz6fbp2bw/g6KknbfvBjEY9
2mkr3JW6+RzJq0ttPR7Eh6ZMwtyQ4V5weP9SdojKGKqENiBOGpXsZrgGhsqzwQ+ys3zVcLwLXdsi
94kKGxB/u6z37H5opmgb3PNgPdNvM4TDoqa9VgKUeRfe03aivZ2W5ZXeUgLXso8mpKHkNm2PpIr/
jleB4ShtBHIhWWSaD7rlFzqFcAhiVDPzv4PJABV4gOhKZy1nd6wuqZs5R3SnGNE/W8CP0zsQPkYo
HOfWSSDMFfwLLyDRSEa0WIDo05T/bm1z8bJ8ge4PNjpqfzTwHVDyWiAUo/Zv7QDf3qouQWgOpI+N
wHe/NnT5SNNkHbhcfG/qYydBeVr+870gwHP9qt6G6eZUdBQJQWaDmc/nQzMwQxtWml9+i22BndEW
yw1J/uQHZ/WfzS1p66RfBYBCtcqV2eOgJhiSwwnlY5uLQrisusl7+uRzTBpkL8R6hhpvdHIT0JHG
5FeIKh+hF8nkuyqIPOB5KMumz/uEeiygM5vEa5FPGooX/YTn9lewuXFg5IzTcc9ScA8bdBAszn8F
jMHzv7rxDwJRlHNudUf0ivXPqQ8y12oXhMYTJRkm5zdaBJFWufloiNG2jES7pDHkP2uTwtlgdZ8E
SZ3koCIMY1LbhmjB1IIkvuiYqFEyyge0CD7Bu88N+wFvFM7eaDksvkMpA2RLuIxiQ9y8WPxvXJf1
sOjWbeUmiAe6FkgX6+CsSJQwU6072DuYWThNVNCgJobTh8eT6d0cuDuefz5bMvMlYcoohoFbq+DB
9WCE9+OP8ruA/tKCir7VtVSNCRKDhftisaNeh+OMbQE/0BNB2z0qZpP7KRDXGXE8BpEuOO84SKsQ
C/4ZWrjLtTtBFrWBt13hzlVh0cd1nhLT0eerIg4cNSoU/L7O+gxR/w+gPwvBvNHVpgg9/OgMd66v
69AlICixO2u/JJOcOheG5MEM6+mPV1KS4dWa1V1llE8f5qp13XrZxWfc0jcVfyzuFs3y+Xi7ZBXB
KMrxW2lGymOmCz1LmAnM9S/jCBbPs+zVv/fxwAiY61I/ZQ6Phg99WeSY/EBmvpZkC/0xu0xO4+z+
7bdQ7mDwvyggJ9CsfItPgaCOKtSYd2FatgHKptCcQWAg/qodPfugV9dfe+MeaI+xffrmsNQgFGWZ
kQ4hLXH/KenSbKhbhVvQ7pIOhWgugQh3v2LGuEGy+qdL8mq9jS29/+FBiLV4LmDJkeJ9gGVQmnY6
heubuPM7coSBvxQWEFFIM8Oe9IOkAM4oJGievFvfMTNKkZq1qGlXEnygo48FiCwD9MRYVjAPT1SY
D2eUQ04Vc13OKeM9R5b2+uJx3xjLh0k0xRzusO4EfajVJsPgXE+F+E7ehBSlWxXNTWfs1LauicE5
pPbEsPReGlCJEQ444BAlmNcAezPuZdWykWHDlrQc2ahavxnQFQ2CqCIayI3Hqte/6EJDUABzDQ5N
LpqyOrDisWcizynICRk2R9gstclfc850XhvqdZuFGAy1W6KKlRa0IbUToGWRxT44otVsHKe6nm3G
mTItyXfn5x7EIuaUbN3K+byAZr4CQ0AZb6Y1VGlYeR/bS4qPc+30idQHD+i2FiW59TXoOvT3fH6K
uD/R9GubzoHrYBWa6lbjBPejMIEoJXz5nko7iQKI2vuoA3fuLzBMy70wIEPtuErHs98Y1E6Yx9gE
aWf+3CXcGvZwktt+wwSbZ3OilmRAxwgWps6X9qFF64k+4e++Rctg+1H9L0ZnExp+25IX841A91YV
oDJT9aZ2jl7T6dXTMCgPKA1bSlzcSJng2nzdWxPeBwe5g7Y3iipoeMzpbvKhoLMx/F+ZMQLfXJj8
iSx32/UOgdsJHGtLWzqP2S5kOCIx7j2/pbClSZYaYOkZqe8R0+N3toXWOx4wpvA/o6gOllV5lTqV
2eH4VQMU7IG6ZfuY4MZWt2UMIpyeY8mY6ZXRgS37hsb92IEbdPz4h6m5xpBMOx7u74HucGTG76Ao
ZCApcWxDovsg3G6aR+dV6hbwmZPaRyse6TjDiv+bLfAkBdOeH78aRpVcpEQX/Erjj9rKSFlCDRj5
IFs+saoltA3WypYYxgSO8Va75tSeC3Wy/aSpFcX2TK92exzGpdqcqfk6b/56P7NHyC2ELhogBTQM
QrUdSvuqh+UWg+v69Uxf3lvS3RVkzreuBv0dPkN8vzENaKma1oa8RF1NweuSD+9BhKOz4chbC8ev
9XOo57NjSwmtdPCPk2rUXNhaWnFouEUVDm2tkgqU2sqAiSxYhQTPvFRRoMZ9blv2YRkpaKtDcOFd
HtgMuiz9NJnIwvVataUmUYE4caRcnIh//sWENnZO/9Dgo3l8m0dnAYOaapE6qwP1aUnJdAE+JVmU
BTmmPGWudvDHsHKp1/hjpf3ihWHS7faaCramGY7uChsDjUNhE7q6RvyGDHMlWwv0mGcPtNIoAFNz
fFbKg0ZCzQGa/X29a4M0VsCs2FAgHnleuzWzMPncG5Tzwya0SoehG5qupmdg7whg1hLUrkm5Eskv
6KFCCkyTQja4KV2ayPscDoxcEijLn0/FCI8mH7iZpKWb2dSl+Pymn1WtlVxwDk6Fz4X6o2d208rv
eVfufZiwR4EY74Yws5RZsNx1Ghy+I2T+OWLda1UMV3d/GdkbqYIdPk9m1TAO5qvfkiOCayAFub+c
rHbaiQxBLrPa5UYcNFvRtF9MRsEI4V6Y8eZTFiQoUtKhcS/pZKnclb9tInR7LBd1WNzZCSUEOERY
O7qrgHPg52qwteWAbVFYVQQ4AWDLJbfCPiIesSdYW/bIqGPN/LpxCMDMz///sgg1KyRWTpne4/gK
ygdtD1VV9euS9AwifHF5p+s+GfRMJpKvjkUgTdemTPA1ljb0JlW4484VO33LQUWZJoGP9pRpmFh8
Th0OYoDGShcmyDjXUhmasttaO2X1d1ccKjXHuMLkfkIZFcjYauLLEc0lS22w1eh2V19pkbcQ402H
0Dcet63ATDmqUHZ6ui3fFmt7kxfC8lBi12DV4VmGdAKlSMaG1g2NWq0zA3L3zJlGT3SLDZbrGYPT
IiTxqWSfxoVMJ2kw7fuAAH+fT0rzNwk1B8W0ZuIVwXSPosrX8JcdUA+C/XmjutJZg81XQOEQGpCk
GsUArqO2WASVK3F2HnPpUcPXfmmdjrthr08Q8vN+mKRG8w1Mrb3NQlJd3YOj542SLL0me7P+KIS1
RniZDaIJG/Ne25dJZsmS28f2TvFvhzY2iH94gq+nSv7mHaH3QFGbzEjONQFEMNOR/tBOp+y8j+i/
j/cBDgDpBA1EO5cXWZpTPjAAsoJaXJTeBk9YOAI0fv3vFvNXU1Lv8RciadyVSx8epx8Ae6Ojoc3B
1dSmxfBbdvkZ9xH/eAHbZNCYwxsqY3E3KLLYSwZasDePBbXmmJu/yM3ZYGHUrkg40atjmiNr8fub
pk2wsSeRgIStZ/zFIRon8xv2HZtYNvslW+Zw7OkEuxDr6BS3rAF6JcuX/yboQBLNLFxcyK/8TGTX
5ICbi/VpGLpoEkPJL3irBRWcEKDDBq2AI3IdivteS+tx32HxbNFU3CZMHrPISPm9Ey8V2JNEPUWV
maZvxxOc35ij4ks5oLFvTSvlRtYDVEwnv4H7RuprqRIptdewVv+hQ7oVIYD41To4NGKRyPYydDw9
sxIJXOHTQ5OKh6tJXfxxRrPL3pk6hibK6z54xydttvRzsm5v7EIpjIrOblqN73WvyiBZ7SNPjRWi
afeR/fCNKrd6FA6W+tFu6GP9Hq0YGSt652zVW9ZxysyCYsNrQFr18n7mI65gLBGa9ZUIpyqDZP/u
bV1yUZ9PEvo+o5cktK+XiGK3zEauMVxfJVzSJ6bm+3U+L+yXqvA7wa5X6cTJRUGxE99gPRLYqKbE
+H/u1XPuJPbbPbo9PNmLRACtGvZLUSAYVZOPdQ9V5InJHC9mVSaaUQS6IhxKM9ly6FwyGxCw50g1
p2kbOzjmYKRFzl45DqQYJjEBIqW43edZzGHeSvYThucofSHz8yPwh5/9Qhe08Sz9NcN7KcHo2D7m
eFKimir+7KUh7NYGWBRd5PBl4Npm7TQdoMQn9806sAHvYfOVn7WZ+VrRKoI31o1ghifJR+V7kVhK
gPY6cwOncqN6K0d+MfhAbd6M3ctMgtz2jNQB0q5T8wUjQJJ/G+8d2TEy9F/7ULEOmpJLQnL/SupV
bWb46Q9qN3EkeVgWuoEuROtL27aLYjPSMUf0CkvgcmhQUDt7vuhySrlKOcx+YHnY/Z2pcz9Rb2fA
i2tj747uPRBB2EzHvjGCMKQaiE/Odd3OiDY+a0tB6EY6eyarglSg0V9OKKZioAv9juyvIjb4MitF
DF8IlPBW6kCzwkxNVDITgPy4m8ENhRIPRGWxISQU915rgb7rVxK8QWYbfc4d2uNpITBAkQ9z3sUT
t6/DVR9FrT/CZ88S28T37+sd3PeSzsndQwNfJpgzLB5b1fy+iMRC0zzR0D2EQ02kRhZKInHghs2W
V2K0F7z7HqjgsSfCkdYgE3gjkOGFB9CpLb7rpRQ/s8RWBg0ylkTS2SVrFjwx4Bo/qyY1XOK4RTAD
5FR4xoEQLkrCkL70FeylKP/6z2kLDH+QcvwSzfGukV/BDEqUHF+0bAhU3viMIUKfKDcD5/A15n+w
hh0RuSOC59FJXRlhYm1yyBUeFxWPXRnQ67yTKp5FQ9F2lt4s/oOtyqb3CC6s0lmEGcKtznXPOwG+
TqnXp/cFyxlwkmDKWNz2NcEZgQaXgMX0PQPqCzaHKfc/xTJry6e6B1nqaoi1Ybh3TuDAarFLn4fO
dX1G693JvnCmzUEMpi2rpbn265Gil8iojASGQwIL8fRWBw6qpxSmk4XXXOVHRFPd/5H0RvhOdeyW
9kYJknpq+GHbApXCDIYCIMWE8VqenWZ9AduUjpUY7IKQIU+241+bMpBhH7A/BBkqQtWNgbR6Ax8l
EwXANOg7TwECI8p8F/DZWeE7kHom2yt75RHoGSYuNCylmDrJCHEq06UwufQ3C2nlaP7Bez1tkBqu
p+jqzJrzUKoGLvEwo2Lb6ERZB1cS4TaNz0NGBwHe9VSIhPN+5FfthzZFD/ycgwglvDf4NkI5w12y
oGgRk53AKCVU5kK3S/rqBUs47Ezho9ha5TYXWP7VOf2QoiHqoNor+ScpX1Z0Qoq609RFtX+TEIj8
BFzqXNurPaSggkeQ61TlZ+A+Hilgr6vAs0/kg7fikNhu2HQ31AFHM/58KGSnO6FlEDFW/IN0CDzb
yfzass6iFqgOEYa/y6FF4MEMYarv2M7POFP6JtgKvFmZZ5F1s3xBpI96Q5Q2FF4SNRh2M1iXlkYr
BEvACi5PRwooYLN32fy6eLGa6lEDJa1udlPG/RaCYx625L15v3ftkJnFsTq3qaEyacYwOxfOXGrJ
dzixdHLgqcn1SZumnMhNZ4A+C9pAYXzSRo1H2zvMlYdUpV0mTWEAiNhdHFvCkFdA48KcfviyJuHf
hc42kVlawvKCqAtBLIkxzCKQBCz20lxsle5DkVip2kAIO01yYb8i0ZVeOh2IFxSY7w2O+OLIrN1o
Csq1YxR+C2ZTmiDqWvi95CqMUno9bZKrEgbaTW70uiJPwXJWxQRyYW4mxpYJ+5ebkXLk4jelZ8qq
K2N7544ExDb+zq8zD3TKw+pDSm9KQuKkw4t6zu8qmrGT9ybK6GU3T2WybCWn2boy6mGy9aieMUxK
vcuHO2NfKJyt3Ckzbe/LQ/fyFCm9sdTOaoDTd6o9SpsD42hCCLlKRHAMHMDIGrisU1uOVHop0BcH
ZV1B3Q1EI1r/8OCwKU254n+vAi49RTlsR4ln1f4qIchtD7uKaq8WMySyhorR0x4d7ExWQbRzGyaf
tzSwhNQQRm2yRQMbLxHI1QKTJPCVH10dwEEeIuan5lqT4icLBPD/eD6GTLv3IAIFgSN2WRwrYSV+
hdd/VHOVUUUGPRnqRhqEYngSeKB9//cJrNbBmkgfP+idrVudLf8h1s5DI5BueXwd6FUG7quPddas
0yOhLRYiiYUw8GHB+6r9Ev7QCgEsaa66Wv05IYDLbrSlyjiHpg/RC2zTogv5NarYgEXvBm9AcOcg
wg7CgTMpMMpVQiXh49L5zq8sawIUCUvMp68Uo3rLOw0qVW0NQQEwGnTSapr9thXTqevpjJh60J6e
DalNdFr7cjr4WrEGRe+UimKPUkGIG9vK5s9Kpz91RberhdYMkNbDho/y2iUlBnmQkNdhM66oOs6m
tB5B9yOya4lknAy62t9n7ssRSeJWNrEio/ZQLcf0bZu1nld5x+vvmNCm/y6e7feBlNi5K9MorMi3
fPHrrs9aj9zDVWCzCZQPzSwTJ6set79xO28M1Kw4CF3HS8yuhtAa7CDy7AhZtdQqs8iQhNnAJ+d7
1oQhqhaquVM3/+N3LJVJVZoF9/hGziqFXnAtZyZCmakW7+nSblWIn8hLjHg8WSTsMDL5Ik4GGzEt
KLOfW2IF55QbJVTikTng6OA19PG6OxXZUQFN6AgzzcHzat7HAsFyh5DJ2/NbBxv89mKBHqsfFHLW
Whky+WzQnS6AAE+78slqi7pr6V8tgroJ2Epn09y6dhdYQpXRHfcBaYb1z+4YGhrltBu8v1U+CZ9m
L0TLd5X79uBvMYtsu+w8BSKbh4m3kZGrufnWzbJyYIK3peKnN5E/P4v9WMwCVKWY+V4Gjyt+A2oN
Cm/pxZklAiMw2OBjOPJzE0/dIRSjjxqxzp/DbT7j0IGv4ru0lc08tlF4oit5jTgQl68j7zcsZszn
PrbkTh4ad99maZnXctgcoZ4vuelEUReMnoKT5tT42lBh+KnsW6W5v2OvGIYNNU7c9v8fJg0mtCth
5VgstPMTT2smn9ek222zMGz26A8xupPf2vT7Z/1DMnJwgkYZuwEclVTTFG2nzWQE+BgiZpXOQtWa
wfEOh+BKdyFwEbQFKLGVuRPgwaybkJMiTk3Uix5eIYFfl94JDZn82wVL509GbBTwBXLDE7xVX0Gm
HR3gYQ0/d61jTT4Z2uJGq+MGmzgNX7BAK2FbuahRmbr4V1QfNG2H6ZhjIP2ZS/6HO7Owg1MC851i
fgXMpOvEqlOuH2HYae8Zp927jHtTc6XHm7vm7RVqfsqomR82grUESYAI3hP7sUmHNekrdwPi5Hz0
ikCv+oVvp47b81b4JlMTUGg5VBiyOGadGGexW4vm9SOZ0J0kKC3NGH0Cn3Qh75VJUjVMSM3NnmTO
hrvex91u+Bp6gJJU8DkiMmjkZwHcemdkdJQ5npDHubkZrybCt7KNtjs46VEQDs/hUgePLopPcHxi
nnRmP4hQ/xvb90B17ur/TMhZio4PX9mylGMYbpe+JUGDWCOMjDfmsyflr8ag9pQHAnTF+UDm2XOr
tlWCEdVJL0j/WhSPRMgziLOr0LLuvFeRhP12SP3saQp5bPRc8cbTpgQy8uZtPnUZLV0nQqLqvm5h
pDNosx5CuRQfVHpyWTedLX8wTj26mjCjsmERsdd1kFx8oAx1d8hlnZlHzYFxbLam+V9HLcFiOQwF
eAZhvCse6iovvZdgM79zm6R06fa466XmRNSdPcd42YsgBNmWH8Vob100GTMKhzymteWw92CYed9j
CGjz5FfT4V/0CeOGTri8bA4LXdcCyRtthp5cX889k3mwLknRYi/G6YiFDW3l9u/tZYKSNR3MjvLU
xGDVOTQHGFVbpWX0dXzkTK3pw4ExLipatlIx7sHJOwux8cuWz5Rguhvy7l2pdir19mmiTaqv1o+p
2w69pmi+M63YMJmpcKZEx/zQmOUrhUO2qvvZq9tOR53KVxHyNnPq0L9vApQy5tGXOs0orA7tc8vb
gC6Lvx/B2/dKtLjiS6YD+hiM4O08YRcfEZXIsLgRyf6oJ0V9xynA4XP6rXlkVlVy0dfEMDwm3Fit
IqicJMERraXWSTR+/wr0ZwOhkoPBEpCclzrZOfQADa8vK8mafy3qft/+1w/MzP8apzcGYtFMdeia
oHwvSMOXTv0KB6T9bo0cihkoKeD+JZE5RDwy88ufjW3oYWf/PrL2JA70lioZBbaw9uqhC3bSwLI4
TnYqrR+GeK1HT0aXdb74PbDPJ5QJaaKUQ2jvoFHxbcdLr9waWgVsF0LVEwFVRrO4iUHJel6kXJ4L
oE33ntEFhCiyyiXQ7Os6+Jwpyj5VmeqSHBN+Q8O2afO+LvR4a74VSdum8+svMuKHoBMWvt2axXXw
MDuWQUGZe217EQg0sFClQadcmJok3KMp4R8VwOp16s0W8lGKO6rnXOBK39pEyJoDn0/EKIRZGaNi
GsWCi+dk/TJQh/ecxTv7mw4t/oeLjevB57NCVF0128IAkca2+8zVnqYeZdUGM+pZuKs0AoYPYLgc
vqSfJHNjNnsGs+tWSnhRRVqHPYEYzlRyesWn1Y8TDfKIElbdtszdsmwJTYf3WiD6Xw7Nzn2pV/Zk
p9Hn6k1Mm+B/WI5fvkdKP1ZBujopd2BCBkvcZyW2kmawjZYmQ7SSSclzzafvjPytrXlzNGuUVRtZ
/Ai+ZIi1tRBZE0BzznSYwkQgEGeGaQRXrOIg3CoU6CsqqXrtRufahgW+On5MeAs5+KyOevVRszCi
DA9fwfoIaHB57BJ6+a4rpokTtNR5fobu5c8ZQWUhDGucnyFMAovYTzW3Xeh6t9uQyC6e3903BOuM
lwk47JAakAMZXGEoxoIQi1SArnCNp0/Bg+FWVURyGeNoyhBYYlFhDjzuMrvKUULbJpU+7yVMNkgb
tKFHwPx2e3NhoRuZZUsRm8g6AFD//4+bD6M6s/XBHTfTtavwsk0G2wMg1azmpiBGy2hFFXj7dw3I
c2h/sOXKm+PN5Eyy+Wa9HigpX1im5Px0RqNc9dTO7CoFJ5IU3F+X2+c4LM98vznEwldRpTh1AdZc
96zf+2v08RyIJ9o5p7AIJy/3Wxn+tUbSjwZLiO/ZOhMXVTGEDHBe5pa20Y4EBXwb6CJHR0SorZbR
kmR2/9uIJ/HzbgB/XJCrPEGaEithD0RFERWKdsI7r5bq4evmm8rBEVxuLooxNzaLvev+fU+MBoGt
9zEqGot34EtGuQAZy4UIzogrwlFgLLf1Vkktg/Hqzpnk6Vjhfpi1+7S+8xIC42kUucD20/adkNOl
3mG2uc4aBRJsWXijZq9jzbW4rxNPsRr8dMCrfaXt4DfArB2rsiCuCeKjIx8ZdBQMIcAI2c4crBNX
6jZF2X9Ho0sPckWHgk53iX/QzF+9DT0ewnDw74fKqnxDT5NH93HiOvUIu0ioGE+eJCWLbAmBUrno
gUyo1oiiaA+MQhTN+8tSd3eOV+ctZ07dlQgX7aW9PAGBvep0l0KZ01CdQEk/d+6oCyoqrHnxuF4L
Zt389jlnAKX3ktkNJXWZFwVwJf3scjrXHgbqpL8PY8GKif/B017yfkWJaJAmCzbVsJndB/nVbXix
WjdlC+gZbV4ni7J2QXoQcucYTPZQYtBrIlBvpRo7TYcFWEmSDyDrzxHMRu+KmOCicVzFq/p7gqAO
7Gjfg6QxD9lYUYXUvvzaG2iZrLgGFg3cQ7vm+Ty/XIBk9TtFFI4Hru8SbkB5iQbLrzsjLA+yayf5
W1S9siQjcEAVr4NDLxXXz4oG6G8DmcDiXTI6maMP3Pk+uz8/sdrhilDt4eaYMa06TCavepPqGZC+
GblR3EYbp/tQPGSKFV3b96SMRI53uF/IYlrWRniWIlJxx6vyJSry9lwXDp78wJyT4geqsSpCcWoL
W0SVJSNrEjsDXGRj3MINVEJt7uw9quiNxWrQtM02+HH0eMAMmvnUWwReuboIut+XZ47xpewl7TV9
cbsjrQ0gFLLnkMtZ/fRaKbJcVBzhSYwJWvduY2j6cy1XXUvqRRRz3X+YEiBWKkiqwGJthRkQFzY8
m/Hvif7n7iYtUb3y5xTd9yINvmkpE1Z3gGCD7Rmp5BHadTUzqAD3bzBUp+NibWTH3h/3zI/f1ech
AmXSG9IDYrZu0YreESyMdeDmpx7DLa1BylQiDfJ3ndBdf/R1EwgQXsbx7E8J4f1iq3b6c74r75/A
wZUxBj5wA7/yfrKmOHNH/6Eblnyb0lphVzy7ybosbS2ZKs8uXmAD2eLtJFxee5DbTji9Z01snK52
nO2Cz/kq2UtSwvEzL75LvpbVIb+U7BFyKdz1sWaiTdThOh6LvKI74enKB45lF+aDPfqTA8auGWwJ
10A6Cd8SvASu+ncM2/xGS2dQmdvJZa/OCmMD50krflVSrCZuOpTdf+BTrb0LBlk68yG4ERqLByUO
KP2cLWTPKjpGXkWaA9mF9DLT5HDGjzDMZDJRFrx7TX4Lmtv/accKcuVvRgqWyzlNmu9XclNPmFa0
63vD3uAfBQFoEOpqtflz0uU4QW+VrMRHt1LdBNfjuGF63ajeYX1RrOVlWpskJyxhKnX6lqNJvvaA
o9i8nLY03aNoE/J3nh8BTJo/K209N18I51s3YOh+L2AUoOgx0Ha1d2TS1dT2dYxFjeqvTLfwo3UW
nuCdUxrWjWvJ3u7OEoPX1zdt3pusKyRZexvixkNiN/o6I1ddUuwc7JLDH6z75VuGoPfdDIMDqlMW
ramsl8CUOp7VjnHaLPGWVPyGSaGZGULmg9K2CknAZJVS5FdCTguJ5vqLsf9p/wkaUC11Zhd+vC51
g0RB6o373GtpKqLULsoNKBNnFdVsi5rRl9Qa877Gicr4AWk73FfGLZjrQd9RvrySwnArOcaWnZCp
9TiprCzHBeX6UpwqubSksoBHzSHzXxyqU2pcOW9yyyuNyOHZL/eIH6jPMFqodgWE59QfrZlA/kI9
L9bLVt1cJ5d1HQpBfzxiNJKdQ7QjG2PP+cVQ7NQQuj7I1lvhJQ/Znsw/8NlMTwLiuZZ6Qr8XpYKy
BiWJieCNXd+bti6gl8Y57ZNb1na0a00L7XPPIx3jZc0E+5lNYSqmQ3Kej8vKib5ijXaNnvz0dZhr
NITwsXZcQrZUKPT7K7DgyE48NTwzYy4avkgrsddKPwX0zWHMhMbDXcMf4rT0lYcGecEnh6gPjkbs
Lb58eEoqaHMXpIgsffHz4axUDks394lTC0UruBisjuO6ThwKT8TC333d20awpD2/X0/fkjgBmtah
LHOo4bFwvYTENN2kPXzHQkVmzDO5eGw/4yHjC88xnRW55TEkGECza9G4+tWpns/JMdxs3XuqyqlS
Uo/XxTh4FaM9Bx4ApHXLPJ+S7F8+6P0whCFcP43r+xIvOGF6obZ7RBhu2lYOyhi0+NjmQOam5UyS
NTPcjXdo45vl9AQ6BZ0feLBWMUtr4XaxIOITCJfQTZ6/Lc9VPPMquJsn5BHqHmj74b3rUmfDedUl
c4x4DD+UVq4+VreZHSLF0aAm8+WN0J2Hg7V6RajENvrZG8RNqQXUG++fOvCEtqdQfAHvtUpD0s12
+jY76gBiJAj2BqyRiG7/RJUQ8fO6M604ODvpwb5fmNkN4WMfWB0PhJkP1YLWaDdOg2+rJ3xe+EOp
5+twBYJyG2WTXwzZtNA5VIMVnVwtGR7nhIy6Nu5+8zSMRrpNxU2zxt14pbnQLN1IAGwfHtmDnlqM
HFGD+WR3knsDt/FSJn9p6XqHImUbqRNIhrb6+mV/6SdRlDlOEo/TEgTzsH+FfOnitfSoKA4HYUUF
lUcjUfL3nm57llCdyGesXl/snFwrDk1KKm7bu6D7SJqLbBwvPE5ZcBCtU3OehbwgKl4sDVpp4PA7
US96U0/qYvbST7LxeW4CybWp7dXC8p4yrtKyceqNVyhdM53jv/YKU3IEejrqL6V27sINzr84PyF+
YumsESJ/4vLWcBwqKmidOTWs1xzXfsf2NOymOAu7BW6eQtyUYPcD5R7VdoB7KUivLSSM4oPbHC4P
k4egUPfw6zhQKAlX67+/VGqIxNgfzZid4dH9VOu3gGV5qC5rJXjIbJmoL0MvvDm6kcsylB2CaUEd
4nxL4G1sVK+TOM27pXYHDZWdaWmei9eZMET3lfP1KOPO8bRbaI6CMfhBjIb1wp+ZH/shD1DOuZ0/
LlKFKsNw94IRGJepC//k8op8Fqam6T0gJOFYLAibBdkIV0qglXAKHq7RZrZjxZ6Z4rGw3O6EDDHW
8hBBRRB7Hr9v2wIXvYNdEUzS0OWj64d2p6ISWsuL+tLJUvsqBHX8U6JM1qQteZIMXLUsVI1OBR42
U/Qi1OXmjJfv4+HjtCarsQ+JpCJBM2TVl+RRLM+JJkmqFmBgE7cMk8T8ycKPVvVxxSNYPPBgc0NZ
YA9+GSoKSqxPODFxX0LaQSw9AM1UCg6Ftvjbz7K3JNrESWCbMUv5JlQcqUq0s5qxNUxQNkkyu46X
q/QF4lBrdb85gsr0CZ40Cr4cty77Szw18xerSGkxSsjwYMRxjlQrH8zfCBJ35NrQNXfBd9KKTFpy
MWYAHfvGsMsfiYNHUPxRQ1LYfs/fIHpaiRgK3xirQ2qzJAN/++22TwQgeDaG4i99xdDkIRNz9f5E
unKrOCKPvKNbaZVT49x2zoRufM5GSzuJ0L6+xqZLegawg2EONpoqAfzAY9NVAjsWWcaafXBiJmk9
OlyRqbzFQGPXdlxyVGEXJo5Stj0FVs9vMPS4HHsSYun658rraWpAW+owlkyEKY9jHkwbFS0SFipN
McRcYLO5bXugqN0C4+4FwTZAFAfCIkSyHaU5172XmMBlUE1eN6f9vrteq/ePRFeETtKgIVIqltC5
+FzFelNRCP5lVHdlXOHWTTuXMk6m9uAfADiN2oBzL4oFejdAxWjDChqdskw6WbO0hdWqxwiKX6Pf
8Zc3Cqsbu90V05pGHX8RPpsd5q2cAzoPFlf5EVvisTfWauQbD/Dg7+REzN7+gWTMM5q5U00wwed6
WYdduUKo760hgMswHBdRlLYA7cxcJlrkPTHm2FE5X6CS0rle8HezMhXoqNIZGG9EtC1u+9asCouS
/W8r+2T3Rd1NdNHffbPZKWvD8iVaCRByWotpDpjeRkq0dKT8PsZQ13yoMyw1BSY7fCECm82Rffcp
+eimmvBll7SQ0sDc9hrU2IPY8ZxQpBqx9hh3GPTM5/oVXsUWLxpSSn5G8FMZTGP9+U8EMHITe2ni
YtFpkY6ac57yV01TtgO9FHh6U/vLogopULLZTgDyo4MBqRjdEmXaGTJ6Qx9EGmrHeoSivNLs/Avs
AjKEUpZMklDlL48chvfIITm55jydIUO7c/phKaPrU+Y72P36bgUevFZpgBaN/bHqq3sY/DEVxULG
J294WKbEhtOXGFZHTdk/AYIJwBNe2bX2tpVMVIGq9R/vX4If23O4JqSX0ukD4HNdiTrWXoVtFGSy
nTlVIyrbiJ5ztXsOBlgDg6hz9/rrjpdQf+ei1IJ98kEESL49Wr6Zy/v6Z35RGdaYZFYB8vWr/z5q
GS43l7dqpBUnJV50ABqdMeGPoRuVm8Xsgo6vJy444TGB8lQRf9Hr4Wo6et25JTfmXnpEvWP2tNQA
c2zgXky28GeaZ3EvXG+bSfGsThMqQXeHMCgnAOnR4xqIo8Cm2jSBLY5jTvWMAsGyf6Bv0ql5CrUs
RA6dDpg9ubrLCrFfLLYAQwSUfKFeIPM2HOpERZw48tfP2ym1Fguah66F+ZIotY5WRyeSQE4AYD5D
rAS/LaVGt2Wk/PF37+Y4/wlrQhHZ8RS9JutzdYB9GB8AUCww7dXwk9G1ptIruNJ2goEEtDS7AAjK
qrZFjNAV4Z7JxcxcOy/ENv2rQWaquv+6SVKUEDIm59sSpoNqPHYV/c2A2VsC4cGGSYwCzmoNbSJO
7VRQmQo7rBLbtvfOkm6+5b3CdILLQGofHCVn5PyzcGcepHHDn077YVXE64cO2Qw1dKckZA4+tcAM
ncVC6Vlzfwcvh/jRG3X+xKweqJGO/xicbPkDDwE5/8ZSF1rGw5azl0/5gDl6ULmHBbo2etyoKa0B
4zkKzjFNcmaQkdsVyIX1SN4gQ7eKLiCE4MDaqUEUwMvQWrzWI6k9/txgXHby5p/GcbjvVwQiLOOs
2PrSOvodUTGgdl0Zc6xxXQI8Mc2XoZPAooSmorw252kbaCiHslXaCmyWMK34w3lm1lAXLWAt8Ju5
dnoksbLkAwBY+9EhBK1tcSzqchh2fkMCEB28ZJGMpQkbybeGJwVkGIZPon0N420FFiBj71tTx+6d
SUcqQHz+oaJ8P1NcR1QinMM5LXfySS1UfgupbtelV889nChCqG+NP8S72N+QCMuJJegKbsSGWjhF
odY2pHrwLvzQR0bP+muRgdHV3q9UizCKs9n0jNMvgRPP+k6TCzO5Z0KuhpB698Aj9nlqUphBuiJB
HqMwkfxisxkO41xSU7NtKOEhbxxhkDzywewiXEAfuzlMu2VLQK9QM/RYyjXCH4LELwwKCdZsznR0
e/r7cAFgdXDhn49kHj3kC6NV9YtMv9rEr5qNGX8CZ60B5MYVzbqg1mIn5VvHaP+Ndo7WYUoLvIUA
kIGC7MS8/DyqS5y44GPibVHR1Gfk8MyCsYgs/7ywei9GuSkLrulGUybQV0IBI7tDvmzB4KKScqLO
fKMPV+pAbjouWPzIZZUkuvR6a44Aruf6ILBRl97KnRZ7hzHNBHPJovz/9V+kQr2JVTxpmK6AZu6k
Dv3C+fE3L2wO+ARgnMauQXemiB/sFBZ0DHRyh+3C0pmifrrL6mQf3D9sm49HtRUphazQ6xLQup+H
yBhZetFUCr6EQlGPQvILtSoo/ye2c7dccZkzDwWRdcQ0HkMkUxmRD0tL2GUIHkYU2vHNzQn56fS7
Jq/8qb62Utp5jwhesBnNR1tmz8d45Z+lHHVoYEQHv10tuxid7FonKom53GHUwwvlmkKAfMSsK8NK
4QMPCowBKdS0OtDxkCCPG+hB+ng0JF50nD/tAL2rzQh1UVzydUbifo7aV342StWjRYZQP8dYPHji
T2E5rObYvQJPxOQz4joBwTF0/kAb03i7BbdVtlnIRpQAJocnUrsDVR/JzdL0BV5dY1ladv5OBA9k
OmlYkgxHgeRStd35+b3+N2N5DbdWQRV3tB0zQZmzky8sjB36wzXUyeYZPJTEuFwBdmZKUkh1avie
o8ewy5ApuPC1D1EdbY0Fa4aAU1QJvanndkmiiYEMb/EP1kLqooZ6w5Cd6/V3nu+TwBFCYEtLUXxv
/hTcH3ZmJULc/9tZqa+yzewWOg/Kg9wSH2KrVrmeRIG6bKXXKckMtYIUMwcgOFHlMjuly43nB8bN
bnOnasbdNnj7T9QMlhO08wZek8cPkCmZr8JJ5fUuVa40E6D1zyW1pJR1BhW0T8Dkaxfp+wIinfSS
kQ3VhhhPDEIGcPkJwausq2xjR2aoSqocasO4bLgz8cy4TEiyLU4JmyOhBS8VHKnE4mH+Ep+Or0fP
K6zOeinYGNU7HmFWHZZWDh804CGW9KL/VJiZwU8hhgRdXelwDCuXtEnRTHs0tc1Wj5kvVyhh5jXJ
Qa6i+/Dnl0Ct61NLEh/fIPxxSz5/QvrPye2DJTfjA+yAtP5lEyykvawMRLmxR0Bqam1/xw3P67oD
hw+P38IfEeg2OcPlvVoWPxvOYfbarumX7/lJWoO9cWb/ruZsznfFVyuYQUgf7ijJ/3yMqXHPHwjh
zVyMRJooT/3UGfy2E/rz9mlsyldD8N0UO2d6UHiLKcuD2AeUz3TKxCS/8C/88OFhsEiDEB0wPBvz
NfNCrkKfEP1QTW8S6mU4/XJxU7Mt9kk+bMbmZx4IpLNoKMQhY9g80keOUrVAhouzIvFf9Tv6g2UX
EyTls8b2+nxwzIjsHGkzgVNYhA6zpyJX/7nxdY2Rl5sxzoe6qQYcyTuLEcxr5XRBvDLlIuwDq9Uw
E2MIDtyzWZz6b2n/y9KZL9xXoUMABrFadzXhSFhhwLZassM0CwshLmwiCApWmqzZnOD2ud2i/WhW
7u72TUweP56paiUrqFqv8bxDteRALUy0ddB5i52sJrUCNh3zoiZ6rEkX5KgwQjJ39CEv8sIhJEBC
3UruMai4Y8N6j4cF8RAACXcZNtfukjP0LJH/KWXVHKahMRyO0GWQUAWGhEb45COM3qUIoeYnFvFV
CTKtdybw2B8iWfPKSzZa/GAKfIb4vhbSFApnIC3zI91ZEppB2dfCluNOIsnBdym91qTdxUcHYu9N
WqYEb33M8lUmMZhXinV8paG1uZLIMGcij5wV4OqqgV/AeP9dnSq/ewkxDWS5fOtEpIvBB5idYGYE
vbGDjuGjbyVeiShJSHHxZYa0Cz8qnFOaiT02Z844RQUVGik6ntdJQ8KT0bdKe+PWHdlnJ0i8oj1w
6Ag48jsfUM2dMoXc8kLqJapVlUKvAOPezlC9XEU+25uQjY4xB3kvud9G0b/Z52bTxDDEx7l9LASC
KSNf0sdoPk7qXZqmhhLRqorZHhzhH3linonKwnnCF5U1F1zV83Fuw5ioYZugYajMcPDcu0FkPJFe
2iGTlwyugAiZyRApVIx9SjIj4MqTONQ1GMJOwF+ce8x2R18SNkYYkjmtx+QdREUqo723zj4NbSN2
jt85ptwyntQmYy0uA2oaTiGwMYXf0jbSIcZGCj9FlfZpYcophcjNLsi3Rk1dokL9dGFRvBXv9i3I
iEOPPmkZdbuXiT2B0jk7feY45NfireM8oKxcK9l8rgmA2BBK4h5W6RUyMKD5cepIWYC/BykAcaGg
++1tx6TuQFY33WEn9L/Sv0+fn4nuoBBBov3E0/yWDOHEvxBrW3D4GxZeNZ7fJD0YUZkJ1oo6J8fr
7DIn/qJR4DzPZ9HRTlzKO9byLsMNkZPS+9V0/GA4fy+WaLQ8ad1jYKOgh2NLAHwLhF7ZFD3zWxjB
bgctu+dK5fR7dY5adYe7SP3WQSiihWQgR+vs4Lx5lcq9/EWcRIA67D0u5SyJ2W6G7+03+sWRj7CD
PAFKbZx/gVoWruPCOfnulUVC+Rocq3BBy/SBWjrKcptR7f9+u0757K39T15URRYERaR/BAMj5swp
DfATgju/vWaJuxvixd93nqOjB1Z9JJVNaT9w3vFRbkG7BfIoy5CVZ82LHe6npKHdEFeDLGxR1s/i
p1EQkN46JF5/2HBkB0xs3XhwjWFTcqJu5tYF94b0H9usoueNnvMp8Oga4RdjdkBA1W33Oh4dfrSQ
rCgwquhKd5nFalD83Ql1jqP4eLnVPX4IuQORw2f5Da6jOW2oENWTH1yuakugTxSk2aYCKvGN1nRV
vL6K7cWu0qklpQsyxNL4A3WnAPCDLjwQ/u6NpIC+g8DSdwGU7FoQrU33WBaxzgkuqoxmnvnDmSJa
zEQnuWt6v71ZqoYrZ/ACbECSu5tN/DNlnpr4YlcrG2ifUdaZuFE7NuW8bFTtuG+h5UwaiBm58rg1
2DDHB08prOA/BRcYlTAMioAToUyUZaJJL+4F9cGjpr+QJ1ohWrTWCx56MwPKEkdv7sVlLQVyvvMI
J+x+pc8nO1X8xChHeBfUqNaAQYfKbyX6Cq7fxqX6L+HwvAQb8jx/nu6GHd6U+ZKT5F3g3iFtF2vR
BtexnJQ3gJHop2yrCOTluKBv5MuqKc427jV8RZlbLEuWAGoJ5NmHgiCrmiGLrcL0FBSIzyGmxOEJ
O5jONmVwZ49T7u5CO1x70AdVpqT94P1Zl6sI4pW13LULxykBVxOyZyrHB7jBxGhdhWbKfWZ44pEo
8EJJnbhi5kTdaeF1fCk2Gz4bniODE9g1K7Wdj3V9Osr9N/M4P+UeLeP40RvbGMKwgunwxgfleLeS
iaX2ZhwJJeuZDg/Mtim0ygxE0Cp/mtZrbILs3TqGeo2U12vu2KsTFLgH8J4UqhFRkE9dUVngFCHK
xbtdu90Mk9iLFEzO1a3mYLEhQ15DyLziFAv9aIecAMbKVSZn593oTMUkno4992XZIKEAgER3xKsZ
5+YBOPf6sZnaYrIDnylvjBy2DB1cnCF7fSV55W4er1w0/RkoS4nB3tfpIIn47bMrxdZWI//p2mvh
Q/kEYRi5e+3Z5ZbVt6heI5zR2xWTvvasLbxrTgGA+tHFxPLNwPzVJfRZyMB/UtGOcTUABdENtD26
csjwcrJwgJ8647X4w5w326HU7TT6bssYF98wz3ILi20rlRIEi7ENY6DnRzlBAhS4jxYxnQn7rU9a
OFzHK8BgLUjTKrNNFtGiHwpkOhtKJ7B7va56kUK7HgwJfR0lc7sW19ZXwtJElB4QsPnxkS34B6pw
yxK944V5DtfL5isFvGy/8VHyJ5DcYpbrEgm0PUGO/iYh5ELAhTLWNbN5Yrl/B/D4+pRE3aCPYq9W
33qjwOhADKy6RX1MJ87IL8hu/qqRuzaQh2WpWUQqSBowXRXDHyE8rEw1rtFm7SchvO/BYUxnMDjJ
r5TLETqX71Q1nzEa0EoiOsZW9k6RkOHzvwMrAvKOvWnUbRRhY+qQUWiydxrXDw9pC/D4uVcpzNcW
rOuBeHI2Ksz9gVPdDM60R5JdDKd9hfDL0r8Lpz/E+WlEhrtuPp9+os0cfO+OwGOMHOacVcqp3rdf
IDGyfckgsnjr9t6q9uFxH1Ia0cMxhMWivq4chJFd3W56fds/DOoqA1wXofDLFdzp1dicEmKOqVEH
yiwG77ZIexoQMAXvF+N51CmG6y/O0Gwvh3JjtrOnxQWTaZP8/rfAwrva98Y8CRR3u+jF6f95V1Md
lTgqBd7ap6MSxM8WCw5iYIhvPj07tHUnJkUHN+H84iuzlTP/30GlA+irTw+9wKFIuEW6FthgTM0w
toI7TsP10v48CpXt60rbKnnBzgltAabZDZfWjAfiniblB1Q/oORtaG7EEcGHLz6GII3wYAcruVdC
7v1VmKdFpIRMhzz+mwcv3vhwD18s4TWMVwktAQ+oWW9gCS/t9xNjDDj7lNrw5nom1sVPC9I18QtY
48sg6zjNY8HCOyn645CnX/5IyC/GDPgPXHJwEpb+rH6GpvZXT+Ov9qxJAf/3DaaXa9abHg9ILvrv
FsdfAnPMPurt0C1UUr9OajmRWZDGe/3fM1eJJdiBPsIxNSIOQUCLrBgI9zNsoI7qMKdXyLltpZUM
8HQYHGSOkD05cIhYW66sY8CEuj2DTaO75GRMg9qnPtAIXxjXvRzVht6kD/FYq/kK9JA/DA2otXa3
Nam5C9noJZ63zvOfmLifY0SBn/0LvgKOv5n28VnDdpc68KFT6aTf97eDrJRj86HMRbj46VKR0arl
kCAlrOeZenwBUzbH89bLkrZ4jmGksvBSeUv3wnUQYQzvjuYiwq+gWu9n5uCkVzfH9tc5nBEe2Tv3
SYsAmeB7Eec5kBwFmJgQglTW/mgD3z6tsphlhwgFmnRDJXWLKYSQObJh/chFquN6dx8+j/J1Tmlm
46i+PPIhOfsLJwuvnrtOSWvo/+QyzWXOoK5HjWGqqwDn1q+b6PdDg2vpQwTBaYF5jSMQk34EIAK6
qy0hUye5wi8AM06ab/AXwWE3CZoCPqqlwk0902sXnTK7J0UC8Eu4caL7FRO/dosZse0pfsTxLLhy
JqZksS5MsFf6ZnC/fwbWHuNTNeNRypC+nojK56xQErdheD7/GeHG3D/NWj3z9h26M/P3NtppIDpT
TiT+KXUVbUh2x4Gxg3k/7WdEuTE4SvHwoGsSA/K3UZDnK/rDxlmAjhMypoi6M0TpEtT3la59DT86
OWR5uyRpLuiSey2DZ1DWseO/wKih8GlEjZ+C/CQ3EsAQ7c7ZpZz5wrErPdcpSpbju6Mc2rPtJNed
PNtIVeDq19bEeeaXI6Ss3EAyBqJVnIaM6EiFa31K2iT0pe0ovu8dM65K/V2gkqpgIiGw9grKNJud
Za6T88HURfYlIURKRAymEj0huy6sbXWUhny1q0Jlkq+YZgD4nn663vP+XAVannB+QBssutIfWraJ
kJBS2W+dBF+HeBKrTWf5mZ7lxP++rINVxW61hdnS0XL8KfmtBVrBwRaKsve6uD97iE/lZ7e5rdcD
jB40mAQAsHw7JX1MtaXVlPMrzB/1ZYoCeL8uZYUHOknRhD30Ufl50XU5nSSNBckz/VIida9Mrafv
fWmMHtNhhOb/DDz6O0bGVHApoSZXnrWjklR5cyCRXtiOv8rWL8My6CePClAN2T6VJTbzq1mgH7i4
rneYcql/lhsj6QhDjoPnCVA9YtcNvDXGSQSD5mUwyfBM4uVRhnsqSajd6gXsk2LeTOaHntRwMgBJ
wNLSTYmmtKrGZRr343c4o3+OUdmNl7mJ87dWhjHzvgShXddj3NZ9xDpqT7EO9D33z/K6eku+Fiw+
EATRtS+WQT/voNrFOWCXFy+LG5YxFMYGIni2PzAEaKt6ju6HUj5cUg0RMlQqZ+etPDOKHfCucMX/
2gji10+tpa0wVuwKGNPZpXDtRyddF/t1ggcrVYYOz0CHD3TodwuAgAcMKwFG3a8WnbXc6xIJ1WmW
ZNpwzqdP7kc8iSos+lxWcdzbLvNjFNy7sg7QOUQbDZAtzuphuRM/8U762D4d/p9TfaF2h5vTBhVu
W5lXlI7dclqPR7Si7Em0kqqLFbPUnffE56MtwiuEJHFi0GVh4upW219YWbNFOoDAXQ9zy0V1FUhU
jSUDx8Wzi34miHAk/FevatCILAL7f2Eqvp5LfdI/3JKb0wSGCd5dxWCU93Bnl1fXz8WdBiru4VJZ
Z9FrVSbjaXWj5EHeHgXj1BD5yGnJw551sSyduV/dMZi+V7/uCVcBbTMO3yD1lq3bMmBpuXkZWXlW
vwkrmaNASz25ykG53l6+LnkLfQFTzt+jhWZOYRHX9Sg8CKdu1G2Gkd2WdvotnhS4+pYwUtEi+rZr
ubzt2dh++U/nH7SLLde5BuqZEISa9gbKNRxd2AJ4jdnsFXdh+POrdTjrJUmgb32PpvLKo7YywaZr
yun+CFP1b1DmCVksPm/goWqcndJbDxjsJi5wTL+abRJMzZftIVQNcdTTQ7oL4zNMgxD3n1yBK0dC
1lIObIc3XbXZaOtAYVtaKU5mTjDLh2KrDmupqerjJXn8LEfQGWbHIggjFkfRebUhQ5xWuqMiEkC8
1x7Zled6mB6mxwUng0iESxCzqPKn8CoX4Pxkbi1Em+/bg0u66ZG3dvSZlhwBcQMixDOoR4/QXc4X
9nUNLxg1s2CdRDSz1ufKWW6CkFJ9u2jfPV0QgGe1eZCcPF2WACGtsmXSGm62gkU3cipzOBpZbKGB
JWQ5i3iLiQC2q/GJRtqn2Q81ovPR4dneBhifthMNgAtGuQWI0r+aE6+Wc+1i3T+4O6isKt5Vn7r6
OdgL4eBGVrdm7H7lPgjKB7DiJbtetYymFHr52wVkngWpVohgPbclw8yyf961zTXg+1OS2q/UlVvM
KzWKU0+vE14dT4YV8Kq9EZISL6lYWAqAKy5NTuh/iB3vLMx6x89s9/fAlts78zDZcy4lqaq8cp4I
gOz65kvq5IbtEXVIc3noVigzPEb1kB1u+fJQuRnaFExDza2pfG2R1T7W9G2y+njdUJ/DKVw3HpZk
t89lbF6hVk5f28WYoBh1IKbWTqIcHYPH39SCUyAzRWVHkiUgbtI9hmV6zm7ptyP0X0tumv+tjdZw
QS7sJPFxJkGaP1bRQM5e7YKRLwcrFOxoN/TJB/wKS4RbuLloemmdiIKo5v5F1Tsz6YPRVYhsfD5y
QRfYXuKT2W+9pIFdBknWcLlXx3j91RR2+Td63AvMGjorwnfYbRNaLM2YtkDg5v/pSyHC2Wx5GMAi
HJ+wk3s61eknUrpjZ5bpGpQPLsY21xPBGsbI/YFDwZQjrGpTvqLU6aUgdgT95nMFnC5cqPaK8CQW
AaFHZhccLxpnSxcGhB+Lo/+k3X7IKTWmU8V7rZsSD3a83kw4GcWrkn65ST1DWeoOq+eWrc/G7L4o
LQdjRnv/cw1cmpsAKz78w7Ew7J1RrGARTvObXo3v/fUoXW5IoIHerOh8OVUIlOjd5vPhJP+CTH/H
O76yE68I0P7+HtSAUvcDOLzBlDEybBD/qmdVRXRJ05Bujn1ijEGimzrXqAP67xiFql8pBlXIOGb8
t5QUqArNUVQsW2zJurffZa6XzNvWK13sPVXGIKXh8Ypubz2WSMKlCPaAlQQQQiQKfGxfRdMDNPtl
6+lTA+LAZtG7nWCxLVqt/RcALCR8srTfKveL9RaMjVfbPFtSmsdBh6xJsZYnAHgzxP3nvpMQ/pDI
lkKjDBqZsQIN+MMngWI8zDTq7JSqMoH/srxQFmU+bEU/fWF88W2JI3RHsYys1kuGHuY7QdD9r4Hg
6E/4esZBROVW7wDM0HsYabmh944QWcJy7uhSgJ05AUxaTUSBtgV0w5Is5pKRczGxIB3TKJLV5YET
uEQc4xzI2vJmHMDkwZfp2aempphKHnj2buyJqKDsYD+xQMdmSLKZRcQvxW8KReJMykLtg4NYZ4U5
R+qLLczOTEgFGPKGenH4HI85p6QO90IxRWbXEZq1IuNng56Ut6ANPuJIeGY9/m3KaxU7ihPLesC3
Jr6wl/ORUITx7NY0mJGoM3XPpgcF5zUMuMsb6RHM5AVM5afohhRyFnKdeX+RVxdqbe8mANgMUn4j
YIJp7NHQVNu2k55CWspGqvtL4HC36IguoefUqOnGtOoPZqCyTK6ZGXzWfSzAiHdOKZ+bBFhg6IlF
dC0Q8bTos/zblLNvReyukEnjugKLtK4ydFaDReIJTHg7mpCJKQ7DNxGuAn8Ok0OBznWtV3+bi5+j
7BgBM4DlbF+bunjBQ0dE5k8fID9xJNcWhoATfriZHfCPNN5A+Frlk2fYIjMcYB6VMDSKQeFeb8Mm
78OlOhx061AuUyx6eegXy86NaalZ0H9F5SUBwzGASVf8J1vpEwIw1bvBSvkhKFvbZdaDpU6mOFJw
dhQkX/N37dKCBHMKtHHmMDot4K+n/M9yOsVXBCHZPfGHH3iYNXlujL6sG+DzwUwTuGxc7wdkFmER
FFY5aiGFXz8AdpeHq76sO5Zn7q5yB1s87XMrRv/90UQWJynMoFtLOK4Z4Klqq05lyBYBKinEQp5n
4i+2AanzLh9V1B5QcnspUterQiJnimqgCUqs3XxjekjK/Xqa4HIZmhj5RrqN+Pf5K+495jRg8hFr
qezeilMTBmoiD00NUPHKi3dAFxz/qx/JVLvNf5Xeu59Vhitckj52gCcLQnDOP4Ve4i/OE/obpwNr
dXgAHHknS9AeOAdpUAV8KEj+DXfvNoyFowNa+nR5YnstMsMyXylR8jzl+nkV4RCcMKFlLx5HKlFi
f6WsxkJCrQmR2SRdI0ByuTnHBvQONIix5ivR1JYoaZtWfGHzuIvNPIitO52FmGfhurjBdVLvPIp4
8OHeYjOEI5nU+lIL3eugeSZNxf4Z2Afg8rxZvlX9CPNGLiGqRQVKkKU8AbqjGbrBIxzKKev+9SUf
NhGDIvLjXIHkSyFgHxePvCS6pH9z/P0DTAbULeL+WtJvqP+4SJmCWbtVUmS/PoM52+7bukFbcHym
5kTunvyx+nbYVEehBoqULXurcwtYVMbaArSDNYfgXgo30LrKpZEDNI9bKHHYuUcNOcIK65enrsD0
R5A1dNlQJ5Rw1z1fhFIgJg9fMEmRXI7WRJ82FlVbuWSFbdKjSk/EmGIE/Rb6yqZb8nvH/APs6v/S
VcV/zicxd+G095bjYAjbFTbssEIdpuo8XE2/6RLh0YgYrYFaw3uQAi6FaGqCXkmJRlLN4D1fuHST
UJ7U5jSMmwdH1/4roqOn1ZROou7K9YmTiVNH5CfpqX5F6EnwfoAHzP7sbU0TK4pxqHvhaZ8DBGZl
zxEQo6T9P0q0qPivjna1l968lhvG8TmnDaDFSU2CEcJYX47tqdtBLnStv4aJm/i2Fg6Alzm6Tn/i
jIMHyk+5yW5ZpiE5k9MQDyNspamDLdU7WFBfKLhj3eRN3O/AGRy4pwPn7+xlPFpdGq2Q25wriqLB
8T0adFKjsvZoURMeQm4ojz1eDMCO2jHEBCDRZEks35AS57w2V4fAHP+UwzlG/Kp5u3UPYsiISbIE
4LMY8nt7qbi1xiCvWyMzTrz+a6XO+AtjxbzGVmrc4TjCByDdTQF9FbQ9SfOw+AKEKLTKIRFOUp4x
wvOyRJ17P8vDoZG8oJdweqoOkzre8WTSKSZVa3sT+eE351WiYjqTQXWpnmZOMMN3hsV56gL/pH/A
3/TYhoGWaaN/5u0ruRUmu4/TSEh35ATbff+scds2of3dZLEa3JDJMJIUdUWr5rH3echTuEzNTlnl
eXXI4Ykpx7VTdbr1g44IK+OdShUBmZuk42lGCFmUx7Sc+uvkLqO6sjEbHTxIzS8WaqOoarBclJg7
5BFmnNw0pYx+ayjC3F8Mf410I0Pu8maQls/y1DskQbta1elAAXFokYegC95QonDs1tULRXRJPag2
9smD1MqVaU+q6MOYIEhp0s5TeCqYNBfaMaqs0f42Hhdja5/VLkPnOYdKWRD0fK7lVMNAj+62y0bs
cDLapXY0tVLRf6qyDjGG/WKo3vH+Yv62sph3Z/gjE+VH/Q9bXosT8ztF349/e5uCngPbwxemKAi0
9JcU0ZJmSVjxK3UTatIJCwyW+tUmfoXb2rmBwu4R2HoYRl0iFgdHc2uHMIUo9o7EVy/3r5Wy5jyd
8KPmvQsAY9NSA9bE5ZThF6QMGrJ+sBH7zklMwM/v1GiIzBflYmbCZyEEhCCMJfk9Ow7JwbuP8RIA
AePWKg3Uu9eG15fz7HhJ0Tmzn2UQVP2wZUt78AYvsh8U7mysOF4ZC++OPbzWgXOHaRSA/XpMAnXF
of/bzZq9X4D2wdI0X/lR/qNWRHCg3IzjMGLlZ6Ei1IV+bsAervPAICAEaNiDhxqTIj94LcuT5XYf
5JFENADBpmfmt2rMDVhLE+gnbt12QC84amALxSJdKCh+ubTuCn2mJFyTMgM7pdE4OZO1d2INqtlk
QBqddkfwRy320+cFvatOjfeyI5KFJeKpttSs3jJcxVx05u9B+WQJWUksrmMvJfHgk+b4q4q/q+9v
rmTjP5Rme+PcJsx0rv6DUw8Ht1bqRu2sjV93aJTnLn9SZpb14G1evbnp5vel7ClDhr7BxyoClevK
ULTho1rfh+CA+kS5jmCbI5SAgBzVbKvRbHUsNfAYe+2Ww/I6RTSMOv6BMPKotk/FSaWLSCw8aBBZ
rxPphKR+FdiOwMcDqd7gPkszuTCStRaHrj62Fv4D3Fln7crc/JBmFhPl45d9EuFv4cbmIF0H4Vmh
rw7c6EXCb+rq6UOLEWS2WDlIzhUkBS4rIk74vszQH6xog9Iz4VLQo8HaLKWZLDbtMIP8Xv97w7gJ
TIckYVMEEToPCN8E0Ix8OjdEDOYMpcsUtIhWReBhxQp4Wm1KghT00+0pN0HJ/c4UvUbKP3Icu2Dd
l3yR8/Zso5/xYcVxYAXjRyIXd2Bk0nTrvJdEMA3zGfzO1TeuN8X9a9SP4xi2aGGUcNMOotfWgbyE
03LdCnrYnBgZO4XaKLoJt7OItzWieAE/4EcorjGsJDqtgNenXgtUDvtF4anV3e7mqDSVCqGhO5dx
5MBYv66czP+HkyizscNBeBuwIY+h+MRu1sNnipEz/ULDKUddOwhdzzZuePKhNhoSUGGZFre+qC/p
7wgR8pxNvj/KwOKJo+ejTphaxYQZyCq7oNxfV5GWLY3OHZaZ07Lz0qguUB0adOscS1dNn+LTMFKG
wSF6ZAv/HQAv/Q6bwhVJkKzJHov5Zl7IxJU+Kmy5x6UBLfbyzwftRZIP3aDRJjhqaxkURJlCScEj
XZU8KLZEb7NhkepAu7qEFixnySQ3QX6PQXj9uQ3H1/VpZFJETnvCyycx2qWX/ZHcCY27oKDbP5pT
0oLdxF0Bm1O1VeDfoDcLfbzv+vVQK+X9SV45kF/oI/miyKmhgOgk0rWmoj84IbyNkWksWyFxIvHm
zVsA2s3Dz+JD7XngvdxyPwc9Aak8J1YhGpsSOy4r27cfLVl/MernacJ+qRzncupgSAqc5m1TmmLQ
66CO4L6t+8n0l63Pr56ePI+LfEe9O/vS09/kJPkk2zBL5M4GcLIyIjm/7IQrqRk+/stc3cvIj3DG
ibueutK3/iMb3+DkAxD9UJrce1QNNZO8NyKCQAxe8FmvldV+1HOErFWhIxYsVFWdJv1ydRjOGFAX
awkZ4Y0knfEwpVpw+fDmMNkNMhcrS0hOxHkJAifnZnwtPKWl84rTPkOb6g68+UCnEsI+VbHRVTWK
pSf66WB7gvZunwQqwEnVFGIBnDIEVDSnpksKFyUMe+UbCFJ9hEgHLkVYPg9Mxs0uMRuZj0MHdxm5
DOdpnt7+clncW4+nGNKV0fA32FmD99sWv6B+XC+zzC2rKTkthaYxKiuInR+2PN581jWftyv25fWZ
3p6HQl3nDY78CnUgEfB9BOwWAoARo1HwXO3frB94+mjbejRGZmcCpu6EINlXfUjwMj6sZl3lKmEG
royFn2CHpNnaM5dnAUmb0D5E8Qni/BSM2yYE6MwPQLfFwwQMU5nwIIpicdUIuWGAnTRtTFPAO6ye
Evj8BLx9RrjHiA8uYZ+Pe6QWCDk95W5mRIr+WrVFhdnKfIEh0PGloN4o+77VCOQ8LbCQUCU30Z/D
CNXENf6yxYF8i89DezkCb4Fr6WtD+BD8xFjZt5aHLfcSD6Hru/Ugn8lTdKSIk5aTFLMHf0GmDf/F
e4ucoJAiYIYPvlH5llWS8MFQuKNxy3khHXAuZUfjfYtp0noZjIZbacdnGamgB+NUKrVQORKWpoyr
d5D/u6OH+eZoi3vkKPr5BmjGYxWPyJqOdRQsVkViTYHd38Ee0MLKcnvLZ6q3A9ZVCSItjIJRpc0z
LQyDbMPkc5rENTnKf7X4uHVHuch4KJ6/8kgaXINYmqD9MEJyQgDYYlSPr+YcHnUXvgbBJ8HcT9Cq
DvlIvi/2VscyPo+ZeiuEeG3n/8B2Ob42NULVGUbIKUclvCJ9hX8QT2F6jj/1jNzYbbj5Epj/V8My
h7vJ4z6FjvnndF2LghCXUly6tD7E2IFQFNlYbS4uIPPlyaLF2AI7fcuug6gFV4/8LyClEXRE93+R
Rha3pS/MAj0sh2zO+0ER0lq0zN74o4GYtVMIpexKz2MY/+gsY1ErLsy23eOBztdOIUjl8qHiwJKo
aUuLWWdbfbL97ttvNi1F7BxVsKnSIlIg4c6CO637TMuGhva7XM14xCSv8j5D0cUCbbssXjAJT0XR
M2aJmrirgW1UP1G6Wd+J9H8BWuS7HpdQxZXo/PHIc0B1XeMHLZDt9dHY73Op0co+pgb2Uo7a0t29
pK0jrssSU2kYWG+AOv4KFi/2NARvD/yLhE+EghV8FR2pGt2BewXsqM9WN9oTSlXuQN3z2YHoofTO
xJ9r+IQOdOAXv8DxSveX2/4/sFytmAFZ1cNdU9hhlYx7l65Ednz+VHWKDMcefVJviuEvfK38Qt+S
Umj9FOLfrwxJReVEnV6wPa+tq83Xir/6me5uJHCOMaYuyCwp2xNPH0IXiZjpz4Td50Tf5H6O+IL0
Kl1SCEyD9JxDK6CMaKYgKjNdOiNTDsBhcgQH33wKCcGGIzMQ6U1vLP6/Xy6GjB3aurFPHbSyDCoy
FixD1Vqq+oPr4T/oe8g8Mn6BUdeTgf48Kw0YUr1HKAsnBZ/L1pACqLpx+ZF5Q4BKHJGETNw2p3sF
PoUgk4i8p8x3QEBtg9cgIaKyTE+6Wemvdqy1rd5d8fazABZAocWgW49ALyAYBwQ+rhb9u/5Cz/dI
xCC4LK7GetuQF1sEtRJ7+8knEAcZDLWbPbkNTarJQj8OxAO4qykemvNMK1QTjX5fEaqjqkA9P+29
gi7M12lDkM3TTkHcMdBczsw7yKLvgK1BIKzPM6OGbD1skR0wGo2N8IKWtXeTkUAkSf1Oq247B63D
Lz681pxpkYufYYk9gXSEZLmlQt2bkYUN3r37SUGHrC/jPU8ytyefmEKmgvBqIBJrwcIUKacxS+YY
Iw4rCBjTsy/vb9+Rwh4op2CCb7LK5SvTyGzK3pSHzEsfUN4tFbojbPo/zzCnoont08gF713RzY/V
Fdd4+YSOQKCSrk1hKQKSmt5YisCvN3vR9wPSAUgc2mYYrAoFvyZVfjKD/AhQqJIDGm1t3O7AcMGy
uApVHiPrHP92zwn79d4qE0nraqH6uTTimZUrdBGc9pGHeGm1zJ0UG/ItNz2GJ2BLtQsdebvxF/RK
JuBlQvJFFeiWuu1XdL/lornWHGKUA96lUxez+xR99JEGYkyv5J2SAx0Ayopw8yFydxVbT70UjBn7
EeTYLB7uFbpCP6cswjPj3QosFQtfjXvu7kjRDxc7HCIQnbh1dTx7cmdZkPuTufuu0mXbhwHbpMrN
xkrZRaC4c8A7lAEjxHVJw6aUK9SRPtfn+rSqIROdCSXgYXPcj0bjZdysKbk0GlOp5MdCHNIZZJwE
jBzYPgb6phvZ4hLgb8EA1du6glYTEGHN9C7c9O2aZwTXJgs8i+KghVIjmatAFqFbmC3f30O66QJP
z36VCwTqYt1QqBsvV/5LGjx3xUuJGn4njox5gnLnfbY+yYKjo/Y4zfXNAOEfedsHvHgoz2GDWFBr
x7qPQcpw43HYGEojApXdiGbFExJzcC6/EQB/AcVXssB7j/EY5RgQHVb6NN2FkrYL8mRNbZQNLGlI
AJqhSpDUyIsIejFKxznhKLATjjAXC2xVpRVGIaTAH5mgQOvvhlDrpiLzJITPvFc+L+OIHioas45p
612pj1JF3Zv8a+arZzqnpPU5xyMbmNAfyRUvh2jIG+oLSVvQRaOHoluB3Js6klA7A8IHQW2ANxdl
AFnlydpWt3J6RldFwCi+nj9aBsHS0hGvpf3I/HmLz76AxD5XCXKzMpbjeGiv/arbzOVDSTLIss45
3+JBpNNMgCxzUTIEDRgHCXS+Zr7PNBbzlYt4PkYd37WXTXxXy2LwCJrKmSodOfvutCAGTvW2ESlj
tmvubRmmY31gNa2N/vCl2DSihJHoCmqyuiGGWsbGVybfNQei0Cjglx91NU0yzLdT6E5ZMSMcuxcJ
VQQnrUDWUyYxOrwd/AJNDIAYHMuiz1yDi8hL4lo0+zv9ZsBXuD4IABX3LEZUrOzG86s7mcLDfGtd
jnLOTslYk8OvYy6NBtvNSXaUmyf1eVkPwHKegX5if7g8f1v40ccz+Jmmfh5AzotYwxVZQq8F7At7
udwd5AwDrf28mi5Ibf864XJlEZxJv6eM2/uCLbnriKDC0mCdRE9G6EY5GVCB/VhXn6WfEyW3kCsv
rCNzNYGlWS8vDMSgqzRDqW4/jUiOEdWhtxCDseoUxMnhd9As+bI7edyCwJ6bPDjWDDkYREIezrI5
OXIft+71p6p0imykSZMZ05zs/g1Fb06Hb5VPECBsuvzARKKGXpSIuKanlFbGZuWl2xzuB6nmjgKr
14zGZPXzej7qhK3dlsmKhm0mboPjLD1t8X4jDIKSJur0hBQiwA4bGe9AYB9pmXZj0rIWbiOWsv+A
wApbTPn6wvOdaRfezQ+MeXTHRNyacx1alu9bnwS10PBvO39NwQQmw56a5sn8JFYacaJu5jINcnau
N9zWTtn+p3UyvBQ5UeD+zNzTfIaMgDLielWvN/GovFeiBooFmMpsPpngCM5rHHqnLwGEhf2dqPaH
tiuS0pIqWvMVgGohQdb7yn9kQXVYb9MPp/y08CGnJ3/wJyKNkgVVuhxENB1y1QaH05LZD6n5b2PN
7MJo+DpogWdFwWwOqA10pIF69ZCHuwZzotYkjEwAA2Qd9hBxV+bsPHtlFl0zGtSmFCPoKRNUpGXM
IorxrIf7MXrlFSA6gxUSqTButIWIvD1zElCRDuT5ikGLACZXoSv1zVZpkJu0Cc3TPI2Wjax3MFFN
+KKalNDP5NYevSaNgqG5oz+2CtlagLwcO5FOJNCF2OBrkzGx1NGmHwCoKzdiGVaTVu9Bs2SnnGEG
J3aY6qDtqyZ+WYzCayxtZofdklzUNWbW28ZlfRUpkJ9rvQTCsA1kUCuh6+Tqk+qk0aiTsr05lbHl
uL3hqJwCy1+p2+jtizqo9wrIyf6jkKOC1dn+fP3FmeG5iZ65zDI8tnpcT1fM9JOsPH/qx28taVEa
mruNBvuagVhjbVRZx+DVBfxKfQOvIYwChMZqLPnjtvoXolaUY8vs8nxeSKNrh8Gme35AKgiqiTAU
bMpfAnuMC2gOqBXgqFkvhvwEwekMvw4/UU0IXMEA5R4nNOlGtMKpAxZAI7nbpUhUpbOQ49j43Sye
u4WZWuGY0XZwQZTySdk9xa1MFNa7tE8JFInFVfIvwCr6of9L+slEhE2YhWnw4oZhh4q34p+OizuK
Sbk7rmSlfkYV9KUaZECELv65nHEYcDBrAnZsOGgfQJpkAmKngrDkAXcObLcU+HNKFdx8PMEvqmrv
NFfZoYBrzkL+/EdCOYBLhGCqh5x8be70jtOJF5z47Q7sgRyW8Joas1WpCe+3/DC9YGrl9unkLsBV
Z95oycY4KEywj/H3/Ek43aO7zM19/y+uJqHPUf7p2ou156HbgVON/cDiIJUfSK1ERgNzbOxYCyhn
vKtp/FlfwALmUldgoKei74FQJQlMpheDe2gYISRuDis8f8AYtCzucea6Bcl5ONvmE/VaOosKAkj/
+1opZ175PHYinBdDRVOunT1ZaFaSF6sy/VDjGe+5hZ0SFm4ycL72eMsR1CWTb3veYZPWY7d+oXl3
1fmuKu/f0O3vSBDoiKxpqUz8qqM6wGDbpznSqYmGzuZdk3x+GDQStl6G5CH+eMCG70ElGN11/coM
Z/SJhvWRgRb9I3sSuICFzGvxTud9uysLDjI5TBWYNddhEP4YhYujCRF7adOCPz4yjokldMGq2Ut+
tZMfm0YZj9rWoYvT921Uds+b9WPY+UzFYiCPXLvhBw5HGyYjJppEP/KEPxeKhhMOiI6HGnzV9q+T
6eVruHoPPbJl6zNLqJczwm2ra8XBbLl/C18eOnxTAl8pdpIPhkwe7k4Q7RuJCah0eDudU0DGjLvB
eo9pUK49vvnP9KPLPKVQfXdjVon5zP/MnBUlboiMvsFfjs9ruHo4c0vsqj1sHiSvT/CaoDze6BaB
DMPapbfgKyDPiRVUpY82XGkuw3tDLplTnuLI/BCev6gLYQ0v79TcPntSNYvPCF10p7BGJudy6zNy
WKIw2SCIuzLV+GxnyGFo4j3O/HUGF4KyWk09jWWVYh5GOyDJAsR6CiZXEEILh+JzT9nN378g40uF
gA3q1q972blydAGeK44ul0RtZ8da3lzk/zqabFwRlACHvNv6IUx7ozB4E6qnDvnro0RJaf+wgP1B
0UXli7j5ONfchgdbm2rJY7OWVxq2SQHZ2qefR9+ab5eKj49rLquh40MCaX4VeX4+zQvV1GDZngc2
bXIvCwIa9pOECVFRuqnVedHUuyziKN0dMNnMJMNN9JBPJ7ZAXAOSuo8EAFw89FcAR46P+t9h7beo
kWB5WYp3jhRnuqRJUcfuRkY/UD3K1AHMZnETu2n4PPI7pfQFfED5X5RjguiUo2ERbF3P0KltNd+2
piAcpKD6Raj3bkE4X3KLKikEYcs7kSsQTDrYLgDLAPcPrh9s+4T64JAb9AmXqgV1eOArue3bMh1L
/c9wKQE/DfH+O5ZI6lUc5lQNz3GP/r+gzJ5ukrg6rd26t5uS3MTdPxRpz9gDjAlfkbXxuKScYUU7
95VddYYrL2k6TGw7kVL46Y/OytCpvn4eTxvQuDXAg1bWuAcoaZzxxcvAmGAfPBTnbBClcmCIrpW3
q5LeWiE7bYsSarYJVBGWxkNBY/7ebA+okKm5EXDEgdlgNU/5UCo6HUB5wX9I1imh9gtGmiug6fVh
C2xrmUymphCy+5rLUjvlpgbaRkJJtoDfLWJmQqFtB2eKiBzACxE5bHXVY+TuPJQYmrQWookUr5mh
Fa5ITthPg5hdb5z/TkzZaU2wH+hXYL+kWLxSjy1AeAaYXUno/H4iBS/Viiqlju4nbf3d678q8dNR
/XNH0dlDqleR3o1UMqDBW3bh/OmQ6NKP2VeutOk9nQK+hxEso8/VPGejvZrUX52cOS4hgTP21eYG
f8Do97uMZznxpSFdREd1u8ZxZPIf/GjjWAuexNfX5sOPAKtopaml0cavq33x/7VhbyGpehx4u5GQ
Vx6Dh4o4smhkVADuQJOC+R9izRx/qZc8IXd7S+ROwYJ92tiXq5eMfdBuE64c/GheqIinesGmig8e
Mv7hcy8uDCzLayVa0tTBu+y+GwFlTnVfgzbO/iFEIM/8QKRD7IvY0Q0h2eOS59Az0htNcNIbiHwb
eFIRssIywTAIRT9Ktp9NyQz7m7dUTQCpv5SLOzItgSSUDSAPUjhPDsw2J46hAzeTS0UQlIzb7Nmk
8wLXLb0vlHl0jieBrqF58/CcNSyjbpuAYTreAGMjJbAiwTu7SFwaGpEezGyZWNiywnaFmXKxJmPL
XLhZC7GjZkYlHerocuqFEjV2GGy4z6CX61YUV0G7gWW5ls+F5C/+UKdeoLtbYWv8GvRTz6Az2PmF
DSdf/IM70Pf7HPggu33lifXUoso3UUP/utWDKVMITNVG6WfpOaur6gKhJQwTO+P2RQVeVmmzzIYb
nW6UC3UqZ0vfVd8bUdyp550q8BmQ6qIyVgzqbGay3nmQ/D0cRT1sdxRHln8wsAjsBHLcSvu233zG
2wd60G4V6gRXpmok7kb1ptCYHjjQBXlRJfIkIHsw9uFE2CxoQ8eVfqg0nSydm1wq/ZYLgjKWE6cu
Ftrl13jSOwEfoAztjdkbEheAS92Op9wwCYbj0YOj+krwU0ErO/XCjRMCRe5UdJrUXWQsClQ2IH7M
nnJJiBGcP9l2UOiqSE6gKWSO1567vONyVpMSXU2XdF988SFEXuK+u/ZrmXv6XTlf1IcjYsL0TLTq
LDbZIRcdKtEtkJJyPxOfH0S03hRA5wTu8zcmjxis6DO2HIEAlSEnNz3TtjJ8nKRJUxP+rLqLlsUJ
LMbqmlUQ7N2O7EBmoYO8Sz4wo/ku6Xn16jVPp6C6+2a0ET9M7SiiHwwGd/OugYdIMei6xtInfhq5
ZanBy4TCmH7M98FXCMd5117gfHcPGgl1MKdR5zmWlxraJecuBa+6LNnzuPY6YmP/ks810JHgkc0C
K6E+hUbRwqmRoycTvSKv8db29vrVYuC4shfr/P0f+m3klzBBJGzA1RgNcrJd3orIq1Z2jlwksT4i
4ugNjPrRIH4hKgs5sSpDQ23cq4I6I8HsHxHmx5UL+EfcvUBXIesLsxkrLGQW8wZD/ms3oJ7UCov0
/haCnY6ifHVxtYbud2zSWPvzHtvqgMVBEhIa3QttnZ0a2t3NvqQZkZPeFMApt2sX0RMkZCjI3EqB
Qs3l96bGFg2KUyW1bfTamhpipo3yOaKN0V6fKKoPhOmZMF1DF1843SrYVma8mliIP5P9Tfs58cUH
wkJfuKW2mGP2JEpJkU4HHDLnX0qN02yfiUranQ4OXU08JP253lH9EVorZTCjt/DfOEp6makROMky
JRN7IBiJVmDpYnxr8dRV12EKJuc05jvXaYD8rYcLJSNaydsAJUN0sZqwyFLib6SGMUGjN1GuGtUS
Ud146xdjlkAWLlsJbmWjicKM8duwZKyBQYsO1c6RuH2SoU/Mznsyd7Ggfqk8KT5xjp78fGFx1vPQ
nqQaeu5Zy93pGoBK57BEKK/Ye4cOpLkCetWVqiEN5WXMhA36UXTOWTlVspuW3HXQxABj/RfndYZg
gOhJyPtbRpcPvlMjmVRkDV1NpP9YRdaSTHGS7MwoyhbjaEdkO+0o25L4vIuD0/5egRqOhhYME1Es
NtYTMi2P2XMfp3swE7L464kpVNM/g/ZVV+WfXt1hRrWhUVKQIRUF+FlePKxwW3QXM6uIPBB9eCAn
d+zyY2k7gNvjEeA0RyALLYmfZnybKrowHXZVwJ9bbNUNszb6bviyxZQ26t4AqzdGC8LIzWLbhBMN
557kmMiaWO2n2aQ5QOFCBTB6c0OmI8T1b63Ib9Sq08H9UM2r7kCJD7yOeeqGO03iZ1fT392FKLOA
3Wey29SXTDen31Tyi2DGTHFVZ8U4a2DiFAll4IGUVCgboxV81rMPvJVZPVpPaJlg9nXZ7lXcGwDg
ioXam7rLviIyDisqHFzASBFDMq/rv/xFEfHFHntj5gN25oRInpkwgPDVc91UQr4dl8fNl/gStG19
zesCeurGNYliM0HUKGeGf3Dw/69WqQzljUYhsn2eI2qPUmbvXplogYnYdqrkaLIF02mhahrpjHGL
WX7me+E0cITFU854BpESkRlEVJxrq854I8uhC5V1mcDwdpQcWXC9lGGF+ZDVMjxo0qXtd9FUVV+W
wKOurGaRIc089D0Ifu5GMYm7s/vOsWe7OhpAV66OAFO9pu+IbdRs/wgW+qxoBQWGXqfbp9YgvHUC
3/3YrLftX1HBBIUzLQ8Q23iw0gpJg03J5RcmGqleAhlEyMg8m47jePWMbLX+zwsxHGlrHd/5k14t
PPANxUuCeD7k9uhEyeF5/p9R3CXxIgEVWBNzbBMpJqTE6nfgPWwH5AifF10be3Ro2ivokx4OXsP7
fx0rBghnw3lW9UkSlJlguBdM1BNP0fMjBALY4PgOjHZduJvT3D8vTBAGST1w9qtJZd8pFG93RPHZ
Dm8E5vIgcwMQoQP3KpPs9uQii7e4Nwf1ay0PBd3bDTdbXywcb08kNLThUNT0q28Tdwq/5TdH7NHA
21i0x7E7QLnfKKiTlMSEO5RTzLBlWcZZ31j+MzWrn0qVcaMez9f1pguoLJ/1lIN6+Mca6a5JTLQ2
nkJiKck01WPSKfIW4jyZvcQyJUS3V2fVyaEsXw1PtJCzGqCCuNNhR4gA06HMu1V8g2Kz/y/3qWHp
Pqn6/oWTQlQsj9kSHtGIm3YxhzAGBxtQMhboSb/1MnQfuMfocueMAwqel6GuxThPAHBBv7tWviY+
0+x5vWvYDgNB+iV5DoyptevCnwPI38UKEqfijITHmg3oXVDAP9rsspK08IgdLGCzDvpMO2iE08gN
cqA4OGzo75FSXEY7OPVI1eJoAweGv9xL2psjX7UMiFfIZPNaNBUzYh+SFrEDsPU76QK/qNn+oD50
Tude1yMoLYk4PyOfCi3cCrs2cK62X/45TxdYJM4Za2h5H25cJit8jDfwlt41wtQu6uxpCuVBKLrU
FWWfOnz+JX61gZ2ALPkLOHWJYcTtS/tZ/Z4YFzf6q9z09wAuGAThnI+iOsPi5ulK36k5FYTDndpC
jxWdHwjtR5N4PLN14zv1Datc85fJv/Wk9Hq2qSMSmktuxocSE/arfJx3Mwl+UjytANsGrwjxlH4n
d0/zHCdfQ/+N8Qi5PG3rSPqJfjHkbcyuZFm7O6A6s+MMAgifhwLNpgpUpmRN208PfmNeLXs/y9WI
p/7ex4Gtam6Bqc0lkhLNIU3UgEaCDF7T5rMCm/gL4s1tAdduTXxLmu+1nDDc/fsVbjLhWr5303SU
vp9JL4aIwPmH//TVqe4IbiLtGrEU8NvxFQZ7k3ADIHx57sodLXSiffk+CNBqhZKII6030tft5oiH
8bjZ30sp6NTFWea4ZNJtnlxdOC/D8i53hIVJmTii0l1NW38cIRAC/htU04iU5Xe2KVnlJHLGPvqu
72O3Wd6Yf275UwG2rYDw+kVUkRtaVn8CAYcZL2vMWTzpeh5mKvFcZxJhsRi1KAk9IYcH/IqGSjMM
k4cUeo28eZmGdY5VSI3ykuVEFmN3iWbwpcjJYizFj/G6j1bSR82ISVyBhq254Hslt2aMJykQ6v56
DQf5S62Mr9AmY3EVd39KC5lP84XIlTk1o2LrdkU4r6CASsR8UziMmDkbKaLOlByrPc6MwQ//6wFj
5HfonN+Jhn0Fm4+Fx3AMprFuxYjwwM1xC10mlqfkEAoTz6HICRq8dYMnvEdWWj1bxfcWOSELG6mL
8Y2I6mVPRgTPNY8Ug2FQ02YxZJYlnp+WXI8WI7uKaLIFBMXHfK1AfIxQ7lGN0N5t3zfO9vXSflWh
r7jPtvTy9THsCV1y2c/LofG1udBblQDkyXKTRATuCfCyxc7pkm+aWc0yUSXjlGQGkUB8DhTAIScu
YB68bkXqcuZWGmljtdZSuYy2W0LMHOWoQgDr9ZES166mIbn+q1XmPOt4Dn73eR4Gh2hTr6jrgCGa
ni/JJ1A/bau6mAM8uawHFhwUsxmcU8Dn0KxEGxY2WG9/OQNW1E/NjgcD+abYXL/sV/IYFtD/l0RF
wO/Jqd3bG3nCnGmYx/7u907lczKRa39oaW/q1cVp825dKlKt1HdFwEOdP5CPhgEg/rLZBZhU1w0U
CCK58mlYTW9EUUzhWjuRC1muwuQwB48LJKSXdn71UMH7H3WYI/UF5G1ILvqAl3olcAgUG2O/t4dG
Di609tAhB/Kcqmq2LxcSCaEc4LVmrnKrvFlh0d9y9pwmGNw3CS04d8S6wz+JvMOg/kXT43uNnkEW
s7EzxIMZqhRQlE8rbS9XrNym8PKhtiMDno2RqA3AFCh4Hl4fmdzO5SCdbDkWYTaH8pvLrQBORRYV
7S50zKwyPI4jjh7oUvkkmBizAxzkQ1wiwEuiofovW1Fxc1HwEPMF5YQMMo/U0IHMnxk07FlUpp39
nUKnzFc1/tjJ78dEVNerSrRTSO9X8FLmiFnanieJ2K6U1LgZyWzyFYW/zXwAvqt5uSnQ0+2qAIhp
v115o5AXyn1B0Sg1DPog5K9rIHN7vwsEGnXv+wWGzKsxO7xRS3hcdzTT+j9ngcDKv0hPvIWwIOX3
qj/ikYRSWFK1jWgGzWZiY4x4NCdjGfJ8UXn+aR+5XRXXadiPzu00xf6B/hmbsRBLzkIE/sb5od0E
AH47ybpBlcWSqpBPrd2CEE3OKSb2KdYvgGGEIJxagoVcyQCzOPj86IZy0CUivsoKi25WTHK3WAHB
qtS64Io9n/8F6mRO8Uq6BgVNqGRibewIohkLiIQh7xfnQjUe5wH5UzAaL2jJh51fB8pfHnX2YNV3
OBN4WkqmbxkQ9vN26hC6h9YBhXsmitFmVn8XRg7+hrDJvo3GnWQ5RMUkd9hkuLjZFHrkeG29Wnad
qi+EBDt5OeZgxd3pUcCndUWTHFwbHyF0TAESR95dI6DX3LotvjpkRteqn2kIer0bUc/1JfDoHMuv
MPi3w2xmXmGmvMo0+K7iuIY/mDkBTvHv4pMMt9MHqGsa9uZ+CXKDuLJq+XQXq3/NrSmpgz/NePGQ
dw72bOsHIb8DodMnhkgwkk6G9D0LWCpFE2NtlrwcDFm9+sieWgijXHCMe6dax+zYUZ/a92aiuVGO
6Jrikrv2dIgabKmeH2wR19Mvs79XuuUHZVvTFETL6M9uSsqikKUiJboxG9NG9JPADYqrmLQ3ODqm
FSy0ZvP4UEcnzm9oP2HVom2VYNKJYhzdMOfv2cnams5dHQ/Xbe/wo7DOGKWUQYDLHnxPaYDJrYC+
8GN7Oq8Kk63KeDzqICuA8eTSrlqfrpPNQC+AZ1XIaJ1T/DFVrzoPYQokpcvm10uU09cE9MKNuI/j
mzNKsKfNoewRASiUk4d2V7a2/YS204IR/+5zmeRfxRImjQULnfSDxI1FPTPlLx3UBK+G3kluefUO
eJeD5QxngyRRyCeRNjbkQFq5GpcNCQqdUrp+hB/A7Kk5Q4kE/rcWziOOMFR/snguoAPj4RXscebr
67/rSJaqAYWnm3o1zPu/sPJTzonsot1vnTP0jqFNYjEAEWWjvieyAMO0lq5UTG7OAWAqm8JHACLI
9ATUYp1PIK6K9jbcl21hl9a0vYXYAqG3T7tFwfjGpAerxJS6+mOHxd8V+A/lIOb6FtOAc8tVC/hj
ZbVMhZM++5wRzjxlHfGq2DVDkvq6HWmcm6TSRoG53rCfvs2qB3Vzo77b+yA+LzEFa3RjvjtV22vr
ry//hzReRf2KTrfzNrA/F/NI4u/kTLgqW+H2JK1XsJDlP1Uxb5HGRo9CPksqxvrzgcEIO4fhwTha
UXsTqx0704KsuC0OTojbAWxtPxD1zwevdIPs94s2nTFMQVbY3HIOf8uuB+xWMNOEstvJBs36mkji
EMk2rnj+YRjgYON5tz750pkA7JsrjDb9v3t/oyEOFUxzIgA8kFw6jKgug9yiiPPcDCYYiVKoPAHZ
Y3Wag0ALRfZYDZ6YY3V7pHEUdvWm9y6ZJvP46+M9FutKTzACZNMuFQMUa+fKmy9zpDIMjxGgpPxH
hFslfrgeVTVbJYiQoMUjq4CArqiTwq6SblmZ5OIuxrZgV9NOyIpbAEQqYBsv84dL06P3w2y5oWmP
rIIxyEj+l5fPDMeUE8r8J/rYWJpEewMwCnU0Shlav32SYBathx7jW4959rxlosWpiF6XdTeqxyEt
4a3n/ihJjEtPiEHY8LFghTLd00pBADRfdNLif+rQspoZXL/gxe9Sli9YUFUlyyZH8w6BqYOVnEyo
/AGP03XuyAtVh4xChD5gfXFhUDVW6R2HOnD14OlL/uoq+Nom0y6ySkbHyWDqkxzEEQfnUuMcGRfp
kfT+TvtYxDZx0f3dzW4VR7A6O29Zr852zCUGUPCW51+crk1guc07qnZKNwlSPELxPphE8uxn1TgK
6JUkx4aMCf66eIbtfi1I+NkxdmpY4RaDCUBoAaROukBj5ulerWOFCGqdJf0YULYumwJQVX0mZB36
y5k2KEi/eUBHbwuYO1gRTuAnKXS4cqeszb01no6ZJSUGapEljuzGAvEq8w9HdfzBq8B6ovzH5t6D
GJbzpaE8AcMs4qAndkPYQKvjnW8RSi8NTe/8/qbPwccj054sa8TLNPT8odAAomDcXwV4BDSSyxN7
13CWSoChgVjRmYOyeTzEr7soDpSHpJreyamxfS/70hh6H8MCATNyCAIKPd6akz1WS0DhIe9izXd7
0UltRtVotAP3Mhh4VTXHXl/IBcFZVB5RRIA19YZt7XJtYjxkdG4oVSpLCtbq6zN2YliVcfo0vgWD
e2p/G6U7YDj9u0eEKf/Z6bc/K+c0XphgD3Tp2tyLp4U+g+Y+AKefogrrnJXNxKVjEjNsnNGaN1HB
PWUhlq+NR0ATzW0C6UMbBQ7sLee+QigZJStzfdgVlIDMPy1MGapm8/PR7TziyjVc520kQa/PyzKt
Xbl1m0+YSIbSOeNtF6KGuq2S+ybjQnY1kdcsA7C+H4+qjkFHyAWUYGz0WsPTVoAXBrfi4Gvxx8aP
WaMEeHCMfiP9xlczOS4mmfN4QfbnLTC9hA4Dx+KgwG3SaDIlnCPsYYDTnl2RzYDTtGyz0z8X7Xof
6rRfr0EhySXUvFrCiIWPXNR70gsD0FQfx1TjxeBHcIR/CcPU7QrxOMUpqv+YZRhnbDCwHaI0pMit
VYjqCudlQS4JZHBxidNASsJ8MO3k/7uHcUPFjy47rPsL1+Woe0B9C5HG1B0S69rm+L/7ySTh3VCs
QhjCnGcTbOJ0XyHgclYJbfihxFykR6q4pesuo/ovNvaqokH35gwW6Rn1/R+vqsqSlN9qCSekvFSk
SdGe6FTumH1/jUG6jAWdx05AAZOwXIE7T6a1783Pqud2jYTpuRZXTekPHBGuotCiMocrzzRHcPqZ
NFPW5tsAsMArTw7hZ+2QQFS8lBnuKPJR7BEBrVYHm9aifRmTyUMmCmKV8CbVtJwyaOVSxzyP2PvV
/ZqXI4F1GN4dW9cKXhuKCHsq9L2TMZa2WwMIxlkxfjxnEQukoHyF5MpuRM1lutJGslelE694L9Z5
9KGchO2iYq8kZz8qm5tSeQHohqesrifKo/2iqQee5qMFlvJ3gqZOmlbYt2w1HQ+CKYGsY5XJouj9
IgzwHutVD2zC+sd4PyDAbSGrz7G8zrE5HYw4BBVaoee70S6tySnn3cw0hkqQMCILwvEnrxq5Gbab
0gHICSSL6SGG+mCdcZptfns6WT5Ivi/4Jz+NeY03DCvj7IfT3aQhqsQqnnw8n3GQ5uyEmtAgvg9u
ecDDDaa3mYzwubleHDvJLLaA0yCgcFV8hT2HsQQgqpzrhRg9JArP+rhwrgogWpw/hsLXRnPhO86u
9SH650+OoB1qtlPDWW00ofgeM+TmP2SI0OqSjIgYJXMzMEh9LqOVstsPcXwYebhhLtdT7KL0oNzb
KwY3DSfx67/aIhYLww+cXxZod+NfUjqClyC97vme3YeXhehZC+s6OfAsBevVUFBylMZHqRQbsIST
orqSskipp/s/DoodqyfPbBfDZfKmbWWtp6LlVVqybQXHTXRTR1jho5a1LETnDnlD7i+xTydA6zgM
e9+Ar0h2YIxFEQ2sRA/KKVhxVRt+t2Of+qsKt9Gm9jxYHMDUIQlBKSWfj/lhT+poHPUcjL/rDjdn
zGk1UBgoG8f3FTxbvQsPLtamKcX+clVkjCWl0fn67KJusGcrlzzyUrm6F9vMwCRzVLDqckhNuEQv
3bESvlVZG+fjajomnyayw2NrqzZxtvpoQRwS180o1IWZiz1WMBndW0Yy3RH8Fqk3pLw8/BnwnBBN
TPf6v6+uUTiTKqZUxR1eWQpkkT+2vVqOKVouDaYlt6Xiw7X/onGzLWP1fNhxFMobsoeDIRWNWZ7m
R/QE6bqSrCg4EIj1fx9Jx5gEetiQTkB+itNugkFQY3OsP3QPJ4ld6beJ22Z5wzv886BeeZqY88al
hZJNIrZIjnSpX6hcScKDwskapDRL+xnfmc0kDEGPztUqfACVBGYYArlPoVEIxIprtJ086JV4OEOZ
Jp3GMYmeQublo76D3RVrY76d2TQEvGsaS7ShTV8T7zSAZooI3zvKj3aKLsIIubwPB7pE2jSWz9rm
GHSbLqukVWp53c/ftkORiRgEPjbu35tKglXLd26hQ1/gHwhayVEfTzW1gvLnhY5xeR8UlaTSHGi0
c0QamDR/FoKje1eSywKEgJUJqLyloD+3HbnJj7zgURh9l+aywe5IrzvdirB0w+zMtD8Oe59y9K1u
e/AJU5qW/Ml9c8UgBJLIpiyt5AJvZRU704piW40mGj17DWDWQf9HoxiTWrtFSCC+/TYyeYxPOHNs
oEm/Bc0KHN67i34miEHpfUXpcN9ny/uDBoQefLNvKrhI7Zffd3KA0Dd41i4WhaPxx8ogvueVtQoi
1rnVkuBv1fEfDGqfrIcsC1CTaP7nrfNPj3sGJlWOpIDuvDS0S3AOww4i5wdByc1csu5Ri8QYqmjY
byLxCp0yV5PBlhb6b8+hq+xGBWsqYLNV7ZCsLSjdQfYcsFcpwPU2jUyEAH7fWi2NSk+TNVJrXy1r
/jUZpckSxrT3HnmjryyB0tFo4V5FZnjdCGB/WXsxBrBqoJAExzkgiHMWTJxtzapVS+zHU/oDqsO2
JLOsXfrQcRmtlYEpWg1BMSjuVGIQ0HlqFaGsskPh5DABzFgsKHUx3X7clLMQt6PG4wGP61uIXqiA
fE0yVQJlhGwHTX9iTxCaHREay9jGSxL0vG7WX3D6DlE4pZc2mLSEt70109MQlJz+3jVMjTovI1D5
VF8SKU8TtQfDZMbQo1pskWXkKpWweBN5qB0jfewIzxFCC+0CdQdWy528HLT5s1/+8ELX38zXM19B
ENNoqEV3KMo/ijr+FLcnc1LAPU79Wbr2p3yyAILK4jo1PqPmoTGKeYLOz5sI2IZjFd005YxGdOuY
33rylo1jSptqh3QE+do14lemQpDXdLOz34YXpj6kUoyOYw3le2qDM259zmT5ZWldBTdcJBthsYir
nqxgySVLiQpvPZ02iUDADx9ec9AIMD7RDaJH1rKWGfxyzVaHZLQ8zGIIxTndpKjlN3khEo2b3bPk
GaNzlxNuaQf4eQvY1pgzvSaLBXKiUHD9i0jxt6sjHQT06sMDV5WHQ9WnXjDTYGcJCgFg4FsMVRdN
EeRyXPMW9sJVcQJOH11zSTgRddBieQTZWHDY+4PK5WK+WqaCu6NGzRqNQLSimJP0YEQHCv+mnQjx
cnSMQR6kn4zssnOAEZYn3YOVaLbr9TI+MhOthgVWzNqicppLsYaGa+WoIpF4pBBqTuhNBv9gY3qw
MWBaenbUfqOugea2uLJQw9+na8mcXo4D3mAqQS3lnWgQiXlw7kdenefU7jqT1eabO8ID/GH+SNYH
RkmH8+rJsO/SrzogG2Pj7TFsJzjtrZvXYOwOJD2Zy0eISxZe1ifeKhMtYCrmtO896DRa2/DEjc0s
NksRvbBwL4iG6LDx39fDluhQfcwj5iV/D7QN3rwRvZ4M0W5uE6C5IW7mtVpULd8ft1NRMjUj7ht2
igcaBuFauPB3FiZ7x6ROhELu9opTMau89tDMgGZEkvARk4ksYVmGTrGpV7cvJcSmY5/2bF3jhPoU
4saJRdrPTyqJaAf0XEfbt9G1eih4dD8xsl+7t+H1Iu7XFHq6Swiy+EVSoW1tJmjzy45X70s1Icq2
SEWnymW6z7xFeRmwaRZlObv+YbLt62T3RLiZ7Y3zTW21+3Tj3R7mI6DX+AHm9JHJM3an+uIdStMf
05bgZ5Tucpkd6KXBXxxMFP01OoDivBy3BMkvtjDm97k5sXK7ntdmm+Tk4/oQKS0rvoDNIw9Y+9v7
nDViPp4tWndNlEjhkc0knmHeHpNYqH0o6F1qkJlIY4i6V+pUpFXhVSNFMOOWrj/ZY6KLjB4IPjGT
6nG8ejq97n+outZV3V8fcX5R6oFOj/KgoTGdTvD9Ud0XsPldvPOMiylwXzTlbXyoCi/DVGC5R+Lz
JtnwKy6g4cLw+xSix/PUt9JApkLiy01leYcpiCwSpS7rDKsXip+6A+j5D4Yov9hen2NKaqGgC91E
7j/U9blDVeqf2694FgODFGE9nI259/cfsm9v+jAy+A0HqwiyCeQMx1maGlzn0MLiJAyvR52iM5jf
X7GV7BSF07mG/yHBBggjxnJovCcWekDkg2/ymmqwATWPtARFVMyLozDSN/Jbh612u3GL1wo0bWjm
O2z2/YB1gWZon9EDBd0zzxvSPYZQQ+en9Z61cQL8U2eNIxFyj+uRf1k5jqg+MnXVDERMA2OKylk6
ELRU0Sy6kSPCZ+lZ30lWP9DcWKdkGckTrVY/YkxjC0gyMbjYCJ3LeRuHw043ZvqNVLXbrw6uNbdf
CfPRkgHgvniUuSGdvurN9TWpP4se7sehp477nmNnSbIUdq0Sk36mWcBaWEx3bV6xt8yC9aiOFvwJ
daCXzt/31CMn/KHIy/JKqaJNkmpGxd1+Htlh8Q0n0l3YtoGmAdDn2PHvkaYoZOzON3FQtzyF3JfY
jgoaqZTcq26wUY++PwgHR2FyoErLzHcoZdbAEpXKrvk5wSWV/EsPd5gXoAjtZsiNzUKWU48wBliu
DnFpiKo7coWpBa8Du9R25EI+9OwAYRJqwAHgLIum7iEIkJAo1pkF6UgTuki3Rf13iXU4F+yjAbO/
iDP4yKO6T6+HaXiGvcMqpBZQDQEppoKKyilvjmvGvesyQ2g48fXFEWL0Sg9uzS7pCdZLwm5KLc02
cu9vWST3//XB3Jb7ywsWXy4BkrIhQrYFQw9SwPV3Gtvl08Sa0QL2HU7DuOsIlIBQ+ttDP+DLsW+8
5iEeVT19e71TWkLJ5ftvmp94PS7omGR+xJuWju9u4wpv+RYrfeXMcTuIyoWMUS5fAG06XvTsIfcX
ZgyQvF1LhrxhbRQJKYM2F48JDzTFPbuFUYnN3rjoO12HdrVDwXwT3lZswzI/9puS4KMwjjrRgpOP
byH8IOWYN7TkC4GtuQZlO8zCpTtODyvoDrrGuwOAf+Hr7NqcOjDuDlmT6lAkPJvVg/nfOCm1wHMZ
fWDAwZToHXi6FlhA30IlMHvurz938gmH+QdoSPWQG96uJofAVFjPs5F/lhYrREA+4TbfK+dgfSRv
RIVrdUxnDrd7gbdlZ24dZzo1EZNZ9kKzyEhlFWz6l3KbyBq/7SGO6KRPA/kc++1KZ+APz1S3nNNg
9Kozy2mUyw4ssK46+ze0SjVOtWi60DAwE7pchOdL2DgGuJQNZ3Jzcl+CQATOEiUEmUKQuKml6chB
vJ5RIuZXeUzU9MMnEJpVxjCAxYRaafChlCDO1GLbo8vC8VEjNf9CBXYG1MmWQlVXpIrtPvT2yQxO
RnP7SHdKqy2dJQ7CR4Z3If8gxW4ttz+khDCHzlobj0oN3Od44JqDk4bZCfkP71vwLehAB6sQYJe7
oPudtWGR6kLtxXTQoO3h3sO6dbkibln5ddJSRFV8scYvJYxNLOTWBy1ZQZ0R3W3nWaWKPw5OxLq6
FrxjE4+OdUS/ufGSfoWALJ2p2XE0YivlM0J8bQJ/c8qqtHT2kADwjnrpyqXSuOt0ytHpnNIMz354
/VOx10AAHKHLQkKQ96BKlZelWhbGX8eM4BOWLmeBBj8ei60s4HFj9bJIo5PacjuobpJ2sYAAYTLY
4qYcieq1gBv3BN12ICVyWSx4sVrJBOqnXOm1tdf8nUcZ1YOcGSuKLASWWkVVFz047TvnmCGVS9yd
mF9rlsD+PnJZumIrjG15Mj+FFt4f84ooDUE/RWn/52SjBg37hjFmkDn/ZCPrSxQU4sMFuLIZX1n8
d3ugaexU0M+InCy5dMsnxwJxJfZwM10X4U+iDZR8EhbApJbR/BE1oOyS3C8+PiAb6SIQOdASdfxT
P1DaLj8B+vvILtp87mzIZ+aLgRpS8vqOG7wKX+JTbUYiJCTzQRaYIbrjKONNaIzN6ahMn/zTKXKU
q6wPl6F393l3RBXY/tC/PQxNkKdLlxa/0sZeUg0xYpMQ7b4Icqn7jhBtqxzxAnoMYGKhXNot5d6s
2DetyQMj+B1WChRVjk6hj809QMNEQq6Mu7hR8vwwCtZQh7uFMqYceZwFDKGSN6/OCTRM2r1cXfz4
REMQBt16y2tzHyN1Tq+YWD+j/MHW+1Kh0sLKafEEpUw6aX84h3QwcKbQqHSjqS6yUh1p7UwVzDtg
tp8TlCMBNB81Eh4h4w0C4iLJn1dYtMRWqnFT4VDg0n0FLMtE+ygI0s2yVI8cNC4YacIDZeeIJYMF
4Xx+O1bQfwxAaI0KnDGC/oybDG9fpjMDu2GTiLwdUgKgIfWB/EWvYc4+/bIlbQH7cdJxA4HRNFG9
IWSrCZXfTR1f+FlE9/pbwl7z1wiSPmyhO9Anie+YaIxTLI1ukTBCyygbW49w8JaLOuEEOW8AYR19
p8iTHRbiU8AsYjTz0YYGMGIECYYadydZfi1rh0NJiOq9CqPvvW1nk4wzraCh4xLwSfkTS71MvEfA
QnCS+Q8oy6iz4e/7fop1/20V99fRseXSBvG4cDNkb9gkeA4Y1NNQ7a6UiHJxJ1qX7Wv6UBxFDDRl
YYEQLyu0/O6Ud78rn+/zitEPQ+Yj269HizMCEvJsmmSftMmXZeS8qHl01weBqzhq5TlrQ3jBQevV
/TwBI4r80eKttIkKdn9paDPJ+PB0QoIv/ypRtL8UUWyYcJgF9SvxoUJK/9e1tsQMBi0Z6NnBqfs5
ez8YhaOdajhtzIxha9knivYnY7tD/cEyjMmzj77kvfOBiflsE96Wi17bnmtvpm2rDOX9r29Bn+s4
YllA7gF2/cx9M+COvquYO5ofwwmA0ZOs9XIgwSbe8YV3nEL3LTga2I2Q6jUg4ARslRI+x10pc8Pt
UZhJi/9Z5SrXLrWTMVKnt6LiCO9moHc5cz+YfXuCxuXe3tiCg0mJ+wuh2AEzo3n6y81/e5FCtZnL
rIQsdPzP2Xc19pz71RJ1Zo0l9MbWuR+mNs1HND8JggMaJecYSP8oOjyiNETWwpWW/fTtmEVwC/kc
EVjM/wr727XnE/7XF6UCY8NgqWltM6ZXBBLDj7QTcEKuIdchYq9eo99zJCkgMJfcPkpjCDeDBo04
tl2Q++9BxkSVtQNLNWSomEP+F9uC0GWI67bKs3YdlBW9ZbKzvuNXFNWjzgRjMJ3ngrXKExLcMRL3
LO/e21ejyCcBoHGzuZ3kcOSjlVSC8jBFshTU/xnDMBW4A7q0pN3PyVK4Tr3HI7b+bRafo0Ds5k/x
65CHTTHyQMlWIqtzt9WVK4ZO8KiCox0U1Aw/SHzS1+JDxZ8vLHe99pDnVkXhBCJwjo/kJw4+WhP1
ngoWVEqbYhh1EQ3YjC1VF8wGCYLxgvuzXbDtBBtvsqtmBNnAnNG9dKQpJNMVbq8ZItMKWZ6yOJbM
4LCdNt4D+iXm0MX3V8gXkqTGHEXKcEWUn4+EKnaSBQiK9aW3TiRmwFsjANjp8MZ9rn9r8k4jsz0S
2+zn1xsuRnO/s1RANkic1Cl4RzQ7U+0HAypFZ81VoIlYsAIDslRG6GC43GO8xVpGm3NrnzbxBWt2
2Hjm+RE/SCPgphrYLfBk9VQAsMTEjCLiTL2+SinT4FB+040PiFSrCGEWaofIBLD8Ym3VaRSgNFjF
Jhwa576rsyjK0Qwb8PU/ER8w7Tav9H8vn00g+vf0WX14H3kHeeQ93jo3isTVBa0pU74ctAUZ/Dlr
0iWXbzkla9MXvHR2emg0/TP9pDJkOdpHtM/zJNXuRSyiM6iqqNN4VZbSUNAfXesXlVWDwzr72QZ7
ZgmULt8luTZhGNKOnadEDpC+3MQvJ8IAIM8KowOeRsiNlsb53e3RcJmznoChk+786LJGH3UzKVRA
7Wq/SEdVSq1LJrOvY1qvn8XQVVmCHPFtB2J1Gi7pap/bg5Z3sTwgPl0GV1igiPcofnmZZllG+dBK
qS6J2It6kiZex4Y9bIbKU9HFd0DELerKyfDeMaBheb7rhkOpY0o74YHaRWzeahiqExNZA9GEAqsE
mVeI4bDA6GzI56To1tWjJfX7iSFF7qbxn59bx9bzSyt+7uBSsA3WYYbv2lByxgLY9w50/nY/K1jl
GFwQcVlLjLgDYPHnWqGcU15dfGHum2z8Q5FeDDf//iVR/Jr9xX/AVHOeeXQwor+OUS5ekj7Fdm6J
12tDzwiLjHrJ46E5dAaLqKcASxCzUt44f27AnghhgMbOM51JILROra+owy1XvLcrvRDtBo0ZtVmv
9bm696pZN8NxDJCBZx8WWmmlMXO638o/I0Gv8/4mBK221ecY8Zz6xCwlsdCK2h9vx6orPFVMclVM
HZOlyDrwc2AsEKOWdjn9hP+GpZkg9fHcKN/r15rdJliZjo66Rb5sUDWadVJ7+FesMX01+HD6EMXp
AX9OS9+ZxoXio9765HFHCvja6ZMrNhUSr6paXGoPSavpSl1gEODq775ADwMTT0Okrzjx+12NuTOi
TOUMexNNCABiksS13/DaGGvZue5G9t1cgg8F8hfr0jp17OsoPbbZGtwk9oCHmpl3qkRIJybCpxa/
mb5IUaxeJp372pZ63G7NqOdEI8Q31HYIKQXAEVC4USr3+e4JnkH9dL2o9ujXtq3Dz/fuWmQuY/GC
w9rMPQIlx+35wrtedP+e/AvtkOfZH3OOYjmsX+ca6f9ppjHyQ6c2PrceCIwANiUj5wzNjUg73g5u
NiwtIe/3jhV51mQxnfiFG5vxvN8KoWb33fv73ueEuKosBlDRW7ZD3VrLBt0iW3BwOH0EvokJTZr/
a3rBwciT061h2eFUsyG2EZtpRQ9rcUdisxVn0MVQmiKxP78KRZVIoH/gBqXrkHiFZHiomBvtWLP5
TMrrRUHPvmYdtGJOmUVeYbeRHYv/2cO+hUScn0GGzHWHb5Dl/95E76TOOn3+wLpyCnn4auGgsgoO
fhm2zclrsvagKPHxhY6go45/mQTGA2DWWElxwF+FbasZZ6744VOOkhOSjbzqsP8+UgeJ6wr8Wep3
ZvxgFK8oFJSQjJqz8J6QgY6kTFnoaMMirK43cUV05ungNAoiF8epbgVq/2FpYyfPjcDRDyzd5AaJ
vufkxF78v0ja2xIuIPUr/kymuKDuYMV3td4cq0pXZIf8efNxAK/HBSqHVpAvoKc0TPYhzh25UC6h
J4JfXpC/eDMeD8BlaJGt8iYzXyz2t7i6CZ9wLzB3PauR8uLufikDHZOenggrEikjUfe03PijRSaN
ilQrNE0YG+86d31HIwwZsXmD5ZKdRxxxEZoWG3ijL+np8YzIyC011V2Sp/iHgNJdNP1zWqgxYe3Y
bKEdXkZKsruSEJmHGDdNlMbUDfk0FgMF6V+Msphz7PMsZw5iDZrXhpa0bQXoO1w1WJFB6YbL3oy9
Y93hrreOJs4o1GG6HSawrnn3jmPPTdgYtZ+CNAR9aEbAgNa6Sl0UuBj/bspvsuA/BY3IteVlMIlH
fMU7u9ie2093LrRcLelNsqaU2AFmNRqMFNXga5w3Z1rUascRDTwYxXCNdO+MKBVHh3yk8LzzhQyC
Q1v/HHFaV259Vt4W7THUQY+0cCMkIi4fFcH4wOr7HFbfPRBiVk7b2MRIb/SLcd/oiytj0vhbRCoV
e3aqumBJsIKuvY6Yr0xLSsPFyNVe8qO2tArm24C5u5bqDfwD49+pXi8GQd+i5mLbV9WZQsmAXiBZ
GWrIl6lqt4Qr0tS4Zu+gg+OqWilDiK7Dxp1OFwY/AOZbRk0Y8EJMafNexjW7UvMMIbGyFSHz4VwV
zaQnu1I02nX5eiQLGvDG4jOxrZA81nBrTTT+j8aF2uyN2dV1s9TKjcN0Uw7IUjDZ83wfKc0XgjiS
a/X1lJmRK2ZAhFr1rOrkKxEqXht8Pz1UlvpueWmrIqf9532S18OJu7tzPQ8+LrDtnk3mivYIAFC2
Ra/UxF9E5CeVVaDXeqMS+qSiamNJ7y0b+LHXjAmATbMNkxQRuEtQ/hFbB6S9/uQm5RaC0NUInfRi
xXJhU9VXUgCDlYWoJ9OG0IwflVjcWoVe3BOUK6xNOl0lO4H0XmvdZNsQa0albrWtiyTiUCGUhBXL
kIEQl3zt4PixwDt8w26Fajt2NP5K3JJHtE3nxoxZfAYox8VVZgIBNYMHKp8XZemeitqcAXJMInry
eWgf2HAc5qPKsfHe2GjXSIz9pgogvCC75eQb1S94hUwK14FfaQ7zuvNfEyGzaVSx1YW/FDe8Ki0y
wpR3Slf1YZRq3jtU0v/6FtIQ2HPrJJtuddxlJo+Sc9y0nk0FGN4MN3YJ5NZdmUv3QS4yOLnpYZ0u
y9O12RRXyGUoFAp/Y/m5VNnr3/PzbahtdwmI+zeIZelstW4oY3ADb9aiAYUUFgCo/dIdYyLDTKv2
RRmACLZox0S8FF3WMCqLXUkrZpuinUVgaGgaYZIB+qhQHYXjZKBSnz9gXzm6Y8Gi/d4lfvgvcov5
o5sCYT58Hx/i3AArJWKAU3DmeMGPDwMJkCiqEJZFNpD8FmbdVwWqM+NvZOHBB0WrvsGkxiRkJLQm
9R5C+t+Fnmz7cyp38VlADsnxb064SBxqmZxKxt1CLxtinC2sT0wuvNNO+drpFPcnsPakpl6u1uv9
5eCrb69572f/sIJqJ4NoVQNjWQqyLpLUVBhC5Tu0S/AaFdyGlcr7hBb7tWqJwoLLJsVk8lT7NB1e
jtLM/lLOi6ak88ETfTuOdq5Cc2j/7Iw8qOvn3+1+wwNndrLX+XjPB2wkrSHNY2DY5GHmGlO2qpe7
UwbdW6VZOzHEfwP9upNqwnzVONZIJhmRhc1jV4BJ/T0OjxZXkGzyfwrBtKbHrpqFOd/td532wCna
0k4jhQWDp1VenLb1jdUnTGUNIEhXqPafzKXdGhwz9mBSgge9/05QBcqhNqGSah2kZIaeHnLeS+7P
igmd9h2cR59FUfW4HdDZWZLkQZhKOIYRR7fjWVNiVuguVsNUQ+7+jzafSNEBSP28x0OHzoyBydd+
Wg5AeKEfyY3DJ/aviGNp8l+kFJi6MgN65D1IVT5FMBmmLeQHH06TTKSS3sh2pfbsQ4Pk3iM2uGTJ
rmlIAkU573tfnx4tB/rHqlXcl8382iSt44uRzHsd6bPh8g3IluU92I9o7Us2JQyBQ2IQDwm7KQdh
4aWKH+hDcKefvOOt+OuL+poyUsSc14JjojLgusUur652zniL029yVQEhkQ0cxjVbloszP446UqvH
u+ViM5W63GNhF85nQE/9BIQWAmu3RHW9fwRgufzb2GmvcZZ4cCArgCQ2PtRA45CvS4LHDGGjH07A
mnAame3PaQIjiXy2TRR6bOoCQV+hY4v3mGs/QyvWVwbTNTRWeRWGx/VpC/TMK4gvUcju1WRI1Cus
Nc+vKuwmapRl6qFlhBRriCKPUc1lRy/Qa1P+kd9u1Wa8o3V2NPgIFjb5ipfNQAqFxNFbJSXC6AiN
CpvryNP19eTz0Gi9wTiv/7zh7aZFmrAiuVkniaSgpilVPaJ7MxjCWqerlvtZPyBu/GpZqiRJt7SZ
cgKxxJ0UMlHN0/agtfwmgG9L5nL5PjJiokttxw1yPg3EfOq4u/HcvAqQmh4E5X2w8Ntz4Wl+mmfa
DP64J0lnomL7LMJWvNPl4FUzHoaqt7yY/EZy1oEYIctZ0+c9BPR4G1EDCHjhhYR7E577maOjQ7DD
LLi4gpTzFh7/8R8FWdPH5nHK0CxIAeoVNuRVcMa7InAQi6LAMYrYuMBusSvl9azCyVNXIo8hftQe
vGdtdO2nfnifgpMQXFOkL5YPw9YkTZjQYGQCcQfU/MxnvZB4+5xeLNe7iUCyg4PhrTz94rMdDnLU
0BkZJxDAhW42Vorjbag9FGx/mJFchI5oVU1D+8eM7g3wu3r8HIStCrH5tGWf01x4R01MzEiDEpCe
KjTW1WkxHLfKlHlTzHnPfRUsaJ7xRT2vPbQ+yz3SnaP1iQYXDJ1nm24Cc2CMv+dm1+yemfL0Y27w
TlcZxPp3ZgzER0nWjma24LFI5arkwaSFF3ZGCJRND6/lrg6A0mXa9Qup3iiYClfz+OCxdSOtyp4u
1du5b4Fm6fXRoNFIhZx33PgjpdoXXDRipNegyI8b98uX528VLATLXH9dmBbkzLa5GddHdk86DEVL
x2VehCOz0RlbfBYfs6RpY1nUNuwozqyUSHgZcjLs2BwTjs8xH8A7lo+Gbg6/rmOYFYjvFzv7QIyv
+cpm+P7M+LhBkikNiUleE1XLo9yRz6rpxqhBXfrCbzAtUPFATbEv5ugWCI7zM5MPHwis4XbSP23U
jK+1QkxvcRFyMU5fo8FrCAnS5jALyIUxVoBr2wHL5DeK3yhoLJYcEQ8GkALuWU2m8GgMm+Z2fUKF
Th1qagiMLgxaOSPcY6/Gq/OWQkEMSN7ZsbFLpJS90txGnNWMOLewDoxzW2+mhXq2RBvILDiDO0tn
tjWXCUayxQzb5gw/IXbMRwaN3TNeVAO9lkKOkpIyCqrbdL1lCJWfDDbam3j2Hl8Bx9w73V3YkMTr
joDowhwBIrPC+0T8Jaca76nlDvV2hWIfQgENvjQsthv6fJClZ6eDKZr0ymiqjiJ37lBzG9nnwCGH
+rYtJeab9mJJEQRFE6ntQV6ayW41VqWN0om659Rej5lNA79w7gw7rlhJR0RER4teorNhbBJx5Pb+
xbf3eq0WBrbgoLBP3/+0b6J083t2I8lsD9vqUb9qe+QOl0182U5G4PR365NNEm2haPJHEtanDMFh
yl+YroNBiz1BkL5pgGFlA6GBeMTHxRbndxwiPMVLJKTzX/ItySlS4L8E7wkHMs6J1RCNiT4o3lpJ
vCYmvo7L1WWfX/dd9rSGTHlm+zjszHZJ7P+9Op5HbUfh9GnOkFdQjJMKsG1qyLi4FX9gtNVvF6h1
bxsK7Eh8p2Bii5ye++yIGF304gL/d/cRk6Emc26tUjx7MxqNeuXcBvK3JbxWzTL6mZqCeQTnbiq5
XXdRw0gQfb0ECOtV/Mnwb/uBdB8turQKguO6mmFxO3TuqqYF8zqrnMuy9ZNCC9xJN0Ys7qjTWfFU
P5cbEyYwmdQ7P6KYtp3Ewhmj6ZX8fmW09aqDZYLoJI5nianNUb2PtwMLonpnLrJZ6l/rjU6GIT6d
oBNtH5fx3EXynz4vOlbL1AUk/EKSeL1X7Q52pADdI8EY6d2h5uWova8WiOuSUwvYiJgkV6IkI8Ri
ciofEBLGnD1awWVoZ98Jha/pUEdSWw8GRO0kHyrwiXwRbMLJS/J382aK2CTiRnd3bFKkSPQTc6oV
ZoP5t135CHCCR5VZgYJagq5r5pDiQEG1jD+s9Xz44ZpmWdfHh/wOYkGHHj83YZngFM95XHS7pA0o
qoXSLVW/M5AxfmHuQMCdpCpqpRemKkol4Tci0BDSsfZUMt6Fvz5aaIZ5pLcBPZ5BOczI80bL9Wo5
sHjaJpahrAUjTdj5Bp7cZSc4a3FMU7t26TQLPm4KReH0TS1tM8iFlVl1AtzJOn5aW/SHps1YdLa2
x2NokzZSQI8nzfOE730RlGB6WB6VCvwvSiZdyo2UbYw36wBPBoknzRy/sskGnUEWNxr7clv2kUZA
17FDnEiBx3+c0Awt/pzd4hMglK8+JkiWygno6aNIgG3tCX34lv+zrcFBXG5gjHJW27ruRw/1NLmY
VPQ1VW8Lr+fZiSNag18vr4M8ZqI1P1MIUmIydhyt5vW3sY7zw4bWwwIpI1+KZ9A/axeN07S3kZMw
81z9/Xx7pDUIxdbgMm826EaN+GJaXfJ7IaIt/HN6pfvkH0mAR51TEXgiVextdcwruPNCh93HQ0Xo
fPH9u5YTFHvFIfv7mYF4SgS09aqd3R7LlTf/ppM4UTVqvimQj5YXq355Q+zhfPWKFBPyjB8fxjtV
oMPQLLQa5GS04HXB7S72md674/qughjzFd8jdYmlI7fiH1PgAsbUI/CLvOJ8kUjE2Vbu8JARXJCy
KpnIrU/velWyKa1rdSWK06mqSS3HloHnNd9h2SY7wdRbeiPfk78DAuJFygcJWv59b0DAMwis542x
olFmM79Z3o2d+X1xK/uYxwwcNLEAuwTrwuDRQ2/UEOBuQJdM8VvDaaBXbPxk3tA2TJdQ/7dsKcaH
AtMHBiW5mOJNumKg8aUMBeQCYAYawWvDbOmMx2jEVmxQAatOTOnuW5x4NP0VOTgUr/hZVDsN0Foz
9zgD0wzseu7GWo0WiAZM/F0wVjcB4fOeLH2U6mk8cx9XBRS4wJ5FUa8x1d4OYmmNiGA/bRCImyqe
BWTfcjJ/KRB0BuJ3cI1MQ8vjPDOKEzhYwT9nMPsHtGRdBkI7oQB+Y9Swbn9S2HDnaQqj0WV7q4LG
/uqZKolC2itLX5/P/FU+24Gr8KtaEq64s3MeHzAkYWSY2vHVlnc8xGy+/pdNMu79sCFj7B3WPf4f
zd6Fjyy8H5Ff+wkLBHjhg3240BFiVtElnowyD4qAhn7848PHffHi9UxX8MvwAj9Mw5eKQz/pfH1A
bFdJ4mt2Y0Oxo4p1DRCImSHKff3Clsv1AIfYkwx8x4NczaXDGOVVPRlV3ei3zfRe7RqsPSDY18z1
xKZ96+5j9NlVnyoOQ1fuAFI0QW58Iy8D1ACgiAY5k0sv0PDdl3jJHg5cOUm2HXR2e98+ewrV9Z3n
SPxIcd0OSUhVxkTEd3ApBTxVMvnKwWnB3rpYFtPLP+OanCea7afMVncrKJciIqF8eDuDEyhwbxOx
BSdb1mcnYGN0uX2/dSJ0rhOSswdkRGplhFYZNRx0tzmpbzqgSNZUouTpT0oZ6FlYcIfm+/f7LpbO
G3QcXdDTitDrJA+T3GeJ2sK6lcYq8lNX48pTvXKdThUid0jTxXQie8Rn70MQLLz3s55Wvz66y7M5
6oN5/ZYF7hV0HD+LEVxiL4v7GbFy1eOI44hYRfeij9TnOnoKrV9fl2d9tat3VBrCA6AlloTseiVB
29LM7szMXU0JF1DhAXxHU0p83u04C7FLPNGUX/fx2GA3TfHrtUtFWhD5PRE8d+GohWX/e/mBpnSY
VCxdOPEBe7B055Pl4YRRknbTAnxhyeRlNP+j5xgGfXVqfPxH0JaIfSMFVi/VztjlHwlFOx0udS2U
QVbYsNHxIr7w7B1De6LayAd22VxwfBL06QMyGNpMKrBKLnoRTsFgD1STNXQKg0nm/EwzTsVwfIxs
2YZOsrp2U2ih4rrNrHpjgWQBv76i7XM/D5CKkbl/FYCMK1Y0N7FQPVmwDSUz4o7QX8TFEB0IoVLR
+uDXrSXw85qqZYTEVXFU00IbpxUXB+3Vj14X+9Z6Ivm0wpyXPWDz2hmG4xjGUqHVGEdnPiOe/rXB
exrZ3vuMqGwM9LM9vuI5RVMuidNj3PoZvj1huXGDUEEKrZeJFlPIwG5JOTljSrDrYS7GfoiPnuLf
i1PPz6t4VE2C3JV+MTvsjcQK9u1k+ZBlt1qyjd3TmxMwty6Y0MAAm+w5+rcOdG0E8d6R2cL3J0MQ
bMObkOc2R26bQAt0Ovao+bJbI3hruDCaGxt0hM4BKgOBb+U8ZE9FG1+UlY4ZFD8ERczpCHRq9xBV
RfwZ2rRESp4tPAEJdgbcUVF5c5RSuxtVCC66veR9FF1EDxRmsZkvehzZaP+spZT2eE14tKOG6I2N
ORNVq2csX+Z3pSZMkp9MngMlTkQgnM9gvWZPDxhoLi/2QJz5q0ODHOa/E0wJieuz9V0KJra3U2Zc
TCWdwiWWmtFgAZodOyGpk/VxIm2AV/qhrwxwU6egm2X1NeXShes3Pv6YtBDkRbSz+X6RcYC/K9Se
KEUKsVxWDW3Z1RSOo6/42bZm40lxA0Okp4m2zmg8ZJQ19VFb6y9Wp/kS9F3JaPbAoahAKOnUlebV
AM+X1l6/xXyuBIENOZRibYkX+WzUWHQUAfiwQqgI8a7g1NCcBWkL8I8OEdJjzN7UN2ez2ClKbnlA
a7ufzRBUaP1LzYkRYg6sS5IxhfjZPiMqjqDpiVHdiWgvXObrpPFkzmwDYoiweKFqIf3h5U5viTi8
u8uPzePKbBZ2vwUaAkNbgjNJZEr8bM73OYw10dqgJg2Mc6nvRz6bLxjaGBspscrrw2uHyKbNr1r5
cEPO2jzsYohpe2toQZKNL1jFKhoaa8B89LkTUH6do5SpmroHHB5MsdkEi4id82da4MCniawUpwt0
fvJPDBLt0IugvX81x3kDAecjivjrQOQGavDx3zHb/LxMNBSbsq0A5u2EhJKgHdY/Fe74QyLQa7Dx
UOOwPBq8fcgY66oBoP7g0CgcDDOqPUThoc+q4NT4X9COQmmMI/MxVuIfD0sFQBD5POt11PjOvyFS
l44q7zXBn8Fku09/SJc2MiPODPMGUdnIKXo4A7P70g1CRQLNI7pNeu8jbgTSCRSyaD62SYbI72TX
3FcbQl5fJ4yTkVv3aEaiSXbMJx/VErmyQsEOtFiq9ZyNkxeF6BQrorypBbAKa/g7KxNvVRFHSdgg
xDY6erBOwP4SFSTjKbQ60QKDrJ24wZwFfAWpt41oKdGOXbhT7CvIOlSaO1ccDiB6Po5PLaMDrk7+
F1axMSrnmriwkaXSz4vPza5s94uu5FxvdVXn0BIcoUZf/E5zqJe6GxZyI18KKZ3b77+rkIRqxSwc
KfKawJnwA4ssy6447uFUynp2R0izHyNfZOvtahep5CRqwFJk0YlvLXyKJvTsE4NeDhSnqHzDlAKp
k/B2Yc7sWj0t7ipvbPBBmBeVRw2WOYmYQEmLWX7b/YcqlrTmrhev9w9H/3h/WWRvGvjJGz3emSWz
HayaLagoSh17xQx1WmBTHIWfwd/s+s4zDsQrYXYxCkomyUbjfTrhfozkdvz9cpZlerC9AZqk94QC
FzfoP00gQrpzjFuXA3WToS9Uqb26p+u5mkZz1fj3sVQvqcU5g6nnnSLCtNoyVh3gzlZ+i0dPhhQd
1G6BmRO39FQCxgypeKj6GtukBw8zQ0rgkLz5Yake90BNGVj8yBdgYlMAw1EZPZm2HrtKO4HgbxzM
tjFZUnCxNMlac9iCtVAjVp7O52W5DY5WrCzGHFViQJuQKqPKUnLLADLd7w1LKRu0h3wQ/Wu2YaA4
bxH1DRgRCgt7Y1uF6D+rPHFjJL2sE/Tv9vZdy5h6T7PTekX6AD3TQA6i9zwdXfc6sR3qvL7MP1yE
snvNUAO+8Xktmz9zbS5MUC3qjr6hGMT5SCdcKn6CfPcvwpUuO0tul5mg/tSF2DK8BoTnsi5fSL3u
MTubPVdxVN8oqKxc0dsXabCad7vVtGfgQV3NqYo/7bAdTYTLzAqOldx68o8mDb4j+d/scjRSi28R
16l/IPI0Xss6EaB7ioK1e2CTNveEy4YOHeYKvlEjjXlXm6u+9B/bqht0wRoQsmsIFBr4crmO5Zng
xF0nfwcjkkxh8karsTNei3rXQNeovPyhEMCM6KTcCGp5LYuW/dLM6Cvk0wg8c5LNdPdISW/5WwmB
LZp5mY+mjo0NrQYgVyDbqRXWtHQl1UvefPMo8BGuFHq4hj96xa0h9EdSzpSSRBbQB0JS2V7vXcgN
nfgW14MF0pRXKvCXW2wvgwSI2ke7BTy/3NhED4t/a8rE9gm5qaEWhq6kQsRDoCm2QWI2oONRdQuy
h+sdDcuQtcr6hp4bbrsMzUWsVxS1BpDFuWEv6a5yHU+3pzzbidyxoL3AuyjIdEdcORV4ekPYhfLH
um0tiU4NUB08y8IFQl9vUGxg7HrxPBW9bTHZKA/maq/JJdCKYrJAi101l+IUGwQlRUBzcBQb3sr+
MmmAu03qsOSHj9wx8ZUxcm4F065wVf35ox0HBrtKdNySTCGcwaqGn9eCyNsg/g1KM3o3WqTkHK6b
eTqCSd5lGGiKL6U8O+pWBMSdGSHo0Pl1muEwdIja0d8Ze2QMyb4ci7mzUqSIHmk7AJ6bRS1wlDDb
celFv3AWjxQuNgv8XRyhR7csVZoXX+KPy5GYWQOPwMCGOTizQBn6zRKqttJMiUe7X2sPk0UCbJPz
qon59tPvyoETjhaePwIlxY4vwFMK9AHm1oRQmTctMtTvRWF15km8AWxBzo8zPo8gsdPMSF+u/dDy
HXX6ID2GRQfdjTyIg09Q3leAZ2HPyZf6wi6npKw43zYYGzVEwk3S33mEZ7Jb8oB1QeMdUh7+6773
whRN2K/7DTfeGQ/BU9dXeyK2w9fveFn/oPSX/Wqn7ZPIV0Fi67Qs4JigQjEBofVEyV/jJ27fuUtT
jmJ6fClL9Y+7p+UV+ba0YPehjP0Hp8/1bd4t5Y4gfJrniAXoxRhoIWpDFc7cDoSIH3aiRBDVJgp9
J8wXtEWeZEsxEHO0IxEd2DLaRJgWyQv98TsOWpH3vdDL4PY/MCl8GwTABV0zPOF8vu7jtDqqzGNv
GpIN3i4hulWkhvL8fBPK13oH4+m58MHo6r83uE9zYCLtTr1PQG+Jm8b+P3KmmoWzlBicGbchyg1W
+IETkJapE6lT+wpADZw0QOiZap1ASi3xIYaCHWZ9CQaMG8f3OkkvN5+R4uEceQN1RLdtf3vFzU42
JDT6SzaGMJXAHS0uXeXaa7gBFPYQ3nbvs1hnJ99aErENw1BjtWcKbimp6LP3YuDJTOz7ADi66ycN
flNcbM9t/4UPJboGLK9PlzEvdBhxlfBtbMaLKJ4sXACMq16JQ1grHfXIash6wd+z8TPbrtZ9NhIP
NLOsYLH+vOUGJDd9epX6rim9L7PI/i8MXUy9vmVsJlvXNKeTo8Ez6fm0x1sHKGaZ+h4Y9BrB2US0
T91bpEI0Ya+Y0REmFT+oj9WBfRRPJjzystHolDDzg0wlbFdPhjScoiCMLpbORWDqM+nheCBubSo4
dbK/3A1UuijPP3XPsVIG1pMQiQUz8QVnlcKRrZ17HHN328L0/p83ToxgKawMq5koR2sZyBsCdpHq
lUxYgIwazwtMLCvM/EpNSdXxvslM46SiOqU3D5kovw9tt3XyJYLBN4crKLmWFJfI5zoRYh7gOWvA
d83L3RgSfYZ76cFuh44UK//8yDZJytzKBWNXi39EE/vZxPnboEx1E+0ZPOFgyW8bx7APnLARF+ON
RFR9kXlNqxcrSypfdwnBfyMkWBF7Bo3kngCu2Lz9EPYIkKt6DvEZfcCpuSUpCrDO3TJM5jMTEuR7
7DDM61t+feqUjjYc8JvmQWrx8pWiuFTRsSTNLLMrau7U1t+TeBlO8sO8MbFQBGT3gGTjRr46cnE4
G/rYYxOqXIphxCHPLDpAFc58zEYdO7olKo2nnMaL2stQk8zSh3qzesUKQtHLB0lt8utAAToTaK4H
OPdzAXYfUPrKy2ANjZoyw/5eFnrnzulyB/PaqYSjyj807SxRoURZ0IGvUmc3K4mXYd32yPTTCEbi
cq71L/4ZpzHdrO0oLDqpBH1zZ+NLRjTLdiB4jTd4pNZGkH79fNJpEOsB3D/oqg33I+B8QbVnPBSS
TmH0K4ddiIja8zZLa9vCQXqdMbySFXSYewp0+r1LnlLHMkRSabIQST5jrOSHew5R4GVNDmEahWG7
KRfwH6nEkNow6WlzXzoiGyCT4Vw/6J2OxR0b7+rULMJ1Zc6oAEAf22SMvqlPaP/nFyFuLudCxJYc
WiipGuWpHK1wwBV33RLuEvghHeCeTtk/1nyAi9EjFtC8Xd/c7wXSWO4pBrunhfr1bs7ZsC3Jj9rP
5PQSlHEJAD22Ll9NxtxqPdapS6W33L/Z4XtsrlwJLJZKKOBn13ExQAznvHAJHoFCyDWwdTdQp5g9
sqABeBCGXbTA4n/4lwrfFOFUe+CoMfXWM3ZQxOgmLukfP9hg2igyj6h26ZCYZLOt79QR8bmMKwkA
T22sEHAZRU88f72clG7Za5MrHQkea2bpLjwZN832cSh6otMNaW066UFax5G4YkelX09QzXqG/7b4
xS5guxdE+evDOEJUoR5nPqH+Z9wGzgxSBsLI3DbqUeB1EaVgbeRoAg2sTMfOP+M1Smc9l18+2qIw
+VZMnQmBm9Xp/jGwusbZKI3Vf1tklnx2LosHumwcgv2zx5Ff9bCqlwXpECQttbh9rRcFhqOcxQYL
mFLuYnntDnHLE50tDs7h8T1h+Ucs0V3vNSRrkEc9QXjfmGH0Pf5j9Hdbc0Jd+TxJaB8rcc8MC5MH
MncbORqStPQxpG3rj8TyaSkx1DrqB6dqAyz2GQhmTASp7Y5K9qutXRqxzPe5KK4ZHZM4y/YIP6jS
0uAqRWCCHSCUe6EE3qkgqvpamuDV1nkT/lDPZDH+o33UU4XEWulAi533l6R3hDtI/DqGGKcOkQrZ
IiQYl/0OwVud2N7k9WYGyoAYcyWfeuz8aIe5OHYYJ1hUWGhiKpGIgUhsRxPiAuj5G+IS4Wb5HGFk
FxdEpeYEtgrGB2acNZ9os8bHAdnfmoRu1Aqs6wC6Lx/qWqOw0z8nfiSyyHYRXoxL/FPd2lvXIbbv
rF1d+dWLzXE4n7Kn2omMVtyuZg6ASe7QGlljStx8EQwAPM+IweoWC1iuSGTpw/0eugdBYpgNrb6r
vtVS6M/2pkyGkwJ1U04bMESf2N1+elUL0X7CJ+5Ulv2FA94FosiWzO6y3aG2f57PH05h4GV2zRXQ
YaVxlQxD/rfcFRWMZ/kEpuI3Yr2eH/Fa7W7O+S5HNJwsqGBp/AsuZB0N6rmLIrEYG+eEQKWABiD+
8UHXjHIneAXEdwAtM3zbIu9T5+HyANmx5V8rYL1+/mN729JT+pV/Gbn7SbltUCpwa+90QyN3SH8h
SqR4vYKdA513DfR91dYhgxJ7JaewF5+SpOTIvbI9NqNakcG7qF5NWx4A3rdNq19cEoYoi+3sL2RF
2eshDC2ermKAIh190SAq4TlEId7kbFALsLmjOZNQ4wQTdhgE3w5y+uul/66nYCqSy9BeppjnkIWV
YI6WHdb6SzWhLeMf20VDpTziDQHC6WzDzHS+z3woLnzIbQyxozWLKFRr1psboP2BJ7k3RwlQ3u8l
Arx7ops/fV7FzAdKdnTxo5wEQx87JREu97GFdBK0UcS9adkzABTDNd6G6D5+kQC+Cj6fhUhBpLBo
EQroP3zcyoszelyQcGh+7ywPJzem+ly31bc6y0Wz7XhHUc+HhVaRXHN/4SUE41Sl6hH5nFdQNedO
F1He/nsAGaeJo9SLwL/eOeOD1X4eviRQCLzKU7jKO4y4mOCPemwoxYIOrVOcRiWY6f+B86pMHxdO
X5yhUoEajAnEzGlOo0RkndrmqIYfj+9VcNc9HB6cvKAdFWA+LSTDI+haOlmqf9JZWcSR9WlWKeb6
h+01UA/7nmxwDT5Arf+aBNFTG8B1y97KceWLXq6ELxPGUml+zEfIoeTKvxXNmYF1nHBM9W26lYKQ
aO9VPx2vdwCapWRHvE2uSy/HD8OVgu7mzT2lupAH7uiQVzrZosv9lAmC8mVWMcj1lgmeZgFTf6oT
HP79pzjOtR81h51K/U5co6WixlBg1JimfMcSQFQkltFJTG7iNd1BkA0Fgt/hLTnhJ11rxn3VS6Ot
Ho9KAbpnjjMOiJmv9s7ZhzSfVrHIPtEcMH/73X4+zkatRgcvK3yFO3DzixAdc5IscoMWc+cdiGy5
0IevAGdFb+kpLDqU1sqjPkU+GfDOXNZPJQ3XdnfLPytJgqulYtEkF9DxTopvrG12Blxha+b5mrIw
8WXdWowqXbuNxmFb6wrBpi/rXpWEMqnaGwQyAlL1nQAaTaOw8cVppQuYmNy4G3gnMqzZzKQIjrzG
KAqnfEv46Z7mmlnL5BHhZtSL+qKKx8628dyxTADmZaVegT2ksTf2wwOHQKMzC3Ui+RujsXY5Pa+r
93OmfL9q0BkYDowUiKWJ3hl3P5xYju3MpJHQ4IhL1NLbQr5k4t4C0lPjvZ7IFBQ1ae2Wk75wF54z
OHFTu1DksvMXRRAEUtYFLodpFqKhxzZFTLB85a5VYjLv7g1Ev1xmy5ff/lRN2sVPtQhnWEUUV3Fa
N8dk/a0hdeOX58DqdNIvaoLa++q24bS8jRDbUdTi5Sf6DgBHYuCR3tG5NMXyC1n6Fdz3mS5tTTa6
1gX0Cy5vA0+BMeewhGClTzlVW5Wy42bjuavcoL2HV8IxOvg9KPzpJGzHhfV78+mSJYN8OQk7BZNI
9d5v69KWOOK+3Xc2UC38iM1RwwD39Od7YDUb6JpcUKz0yafwHOphoLFmk/ZwiPPoqcNu4+X2fJMo
9bPolr6pgbzazi8qiHDDIjKxxiBSGDCmLfyvXx3/O7Kji56ZkCnSe+1I2t5b+WWxcpjdlJRxZ5I9
UGvUmEA5kdKZhOa+8vFI2qisa+dmN11iqgxyBdJDzOu7nDbzY16w2vDCnpiO7EqZyNxBmDSTd2ru
TVUsc++uWk+o0zk4Hzp1k9jP50xo+R13pkR03hlDKLxraDx66CF0t+38kzg6tEUIbGKSJncjvDho
u2a5AoW1QolEQWEk5FK82dN3Zz15tGYwNjyS21ZUbdsBTcot3V7dv1rDszeNbomMCFXOw7U4mzwC
RnzhkL0fmWntuOOffnL+4S949nLRFozoNOj3WBdp/pp9xW4trJ/K6Y/NGpO6IUqteq8YS3K/HdBi
DPidWpmfU/kQ0KmGB5+wB98DVFE1NkrDYkuXsHGjaBcfoNMiKxODD6fs5kzL27Ij6ZhBC6u69rn+
MVmlhQh6B6haBQ8ZOp+3ql1H55bXA/k0pHBRhoMnZxGlnadmjV74unHPNSTaAhZLAAGhi/hNvij4
1R4TXKXkWd/n6QBl9tR0EYzYLzAZeKroceij8nDJvYQACprm+/vx/EATvjWMHphoGlAhloo3XueW
OJUyUG5KXYmUr9wv9YbeX87ffTpnNDkoZQNVGLR46muXhxqDJIISlCCViG/q1ZcykK+EipT+cvmg
4gJjGTTeL4uRRfq4Lh4S8HeAoJp+i8mxMQ2+Ve3WnNOQg/fX7WImpTf2PXUZixoZrKph2djeEJqj
nPxaq5jE0qHiu7HFPYN7M4S6ajrjGJAPU9B7f3mS4WjPdEAEOEoyXHQZhSz3bzZH/ydK4Ebk+6uz
cNdG/nc9YWjFzaxnWPVzJ8Ckvvi5F45fJoGxolL/UTc9fjdAWu7+KJefhW9IjBLidWcmDrpkNviz
hhKnfRwi/3dw63K6pIERifLDrRyRWWeLLzhKCidESaaGYQ04gAyCcWAAj0x7X3ijg6cdR4jEbvip
naQV6MrMR6bEWsHDpXFcZvcDF+bI7LImHaNnBaJDVY3KebeoEpoH+bQVeRW6iR7raFJEDeGtZSHJ
w4hhqqW2Ik4RcREosc8rS2meX9gQWLSVcS5BCfG1VHqRJKzogbbxgj/RE7h9IA4QK0eW+XKZm1af
Gn7e4D1tGBe1CSwZNie2KcdLrLGJCdOqbIkcXax7bHvmNNk9BOuA3wk2iOefsfAxVaVHTpbv2wcO
+wHQlk1gEPGLxmPiPKbD7a/Zbb/OcDcDNxuY8UQwGy8CHs518v7MaTTh+CHhUAxbsEoppPIIdqGb
IoBXszVK6XMHrWWEYdCC97+S/+150C0OacobskYbtjCFzTp/Cl/zdwEgnY9DAvRheotY8R/swqir
gGpRsmlcgttb+pj+rQoYY8sFlxGW5eap1tE4tyD6bKKEZB54uhb/X7te3Wynnx+Nk3olYwqXSdj2
zlMK6rZUdn96in1NafAlwg3kbEtXdIWfGCxgkgQAFxCGZdFq/K3aPirTJCSTdsBgsKl4GLq11Gy8
6HHuBv/GGRE5EwYCv+st0aFYq+1T6uZJGmZPrk9P3f7eGvT1gyWZT9tWIldtPInl8NQDBJeQZF8F
tQh4R02iWV/drXODjZSq8i9UJVAfCcfeM1WaQGw+CFNxu25ddiOFdTfoPpY88agX8/hfKGN6Djo/
x150YgVrkTSbDRnKlu84pt5hDKr1gvwlZwUiVgvlwnV+VYhCjsrt2dhk3s3wGvSUaVlprREUAl9z
Jo9g9l8uWFBgG+zUe1yyJl9oRCqPhdNjbyVTkWCfmakHweBLKAhLtNh8TiVyc8GnfzT09kh118wj
vLkK0fM9tZc6dVoGfL0Yqh7PPiicIXeEf15svjB5uxP2ZKpsUo/VaFJbESHRxtjPFLIS5Vgop5Lr
NjvDimscpMBu/eGE1hr8zIWikI1BlIdpsuoYoXVQFUZ0Y57VzPvsU6WkcjUwuHqkDIvfMFtoQ4cF
DD2yaWLtqH46+0epeuH+BEqezgjtalVxxXssornxxlklPqQd7wZe4z0yS5UcDg4jsym8xCfhDSyq
st7HOangJ9exh/vtkvkn5ylWQ0CRp/Ridpd/ITYVAnKlA8PGtKqD57rFNsu/CWKLy2LNWoDhTAM3
Sz4frji3phrJFLPCDABc7nTi0M5KLDdrVwLkWOz9HeRfjOMsbfwzhz4PXMUmz88oDjp68+fPwpOo
Gr2qpkPYqncVR4QlUIMr8b4JODD3sVfc3y0VXOev2xrqRNZRFCoEkJESUsPPpeNeXqYS1kbCJH0e
S8/jCTyjFqIoLvRITcf9vREoHvdsymgbvVBm/Tt6cKR++8hDxkyGXSTMton6FnNgFMjv16qN7tT5
Uv0JJjEo53rKr9R+vOpmk3khck+nEHyqIBZhEwv5pdBGgdSSXPIaF05EK1M/x3hkxveApWkUC4CA
auew259DwNQwpX+TOlThsaTbCI9qXKuyIMrgNFpudg7yY1Eq09kp24RbSpqnAlPdzmXHd3Fsnsys
fXj5nU0wFP8SlLwujgrn7XpzmVsUrRLqKBZHD7wwxTczorPHbsWF6DsIwgPsmOsJwCc0kXuZpGzo
IOwrTT5MOYaymLc++ENNuX4rzFbfwOKkkO4Qt3vyBynPKpgXB5L2XGmxtXSK/mo1Hf8pKZbI3RiS
DWQ7dL1X2B8i5PbS+GNmb9HOZoq2g0cakwpNMJ/XNlq6g1JHinzq6RKqaRo+nLJ0+LaMO6F6vgG6
4ev6FQo8jaXGJR2Ul/dmZMTrf2O2gpCA0PJkTc4FiOCtCe/vE0+cCq0ZD/7WafUGFI1rLShoAJap
kwjSPB75wjoi2zBGhpCJmQ+ZKerIZDLaAg1plhtUyqKx4dEigIVL86rMMs+6WnkoRrT06Rsx31IS
A1kPQDoH/yRQl0S8V0LXDhzCYr20WBaQskULOf7yVu07F2a0gR6Y8u77sxh9Drsjhtvc6FiRVlrv
TX8x8GZs3e9pxEEoHmBLOKu5Q2AQJiRiWSTSpzW4Ee2pSe3CwX2gGIhFQa0DyuLOcZCYyDP+5xCH
Uzm7SfqfvNoDaEjRs7oxRKwLXAIT1Z5/6jmEe3TLAQHw3bmje99hV0fAEiYloBesUuF6nq3m5eWQ
8VSiqwJez3HZ3+EhKWkNLh9d05VY/BpkLADaUjalsDpVJ3XlsqGvwWTRtDM4nCfPKpTbKTevRt4O
xSTHQh/sUnpsdRpMBp8CEzREZhmwXHno1qqpIJzhUWKvjyxhq3kJxNgAGDEJ7Ish1SkVyDFcCZN9
SyXg6ZCtNtNrg8ItjNwWc1rULGN7Yovk1Lo/shhzS5Qw/D2s9EdmReTuPwA5GXXl5hV+4R004h8C
3Lrfaj26zaYcBC/xHcsNqH1oRHLqQRdU/yIP9BYfpKq/HStN+fsNbc3zMGN376aPkt/C8ZT+AP3E
K7GHpTFrQBFxyykeBQ+7Qrf17oX2pJp7DYRq7g3NnhzIboCLcciqkL+sUSpC0CeMF2KW3OqGY3+2
/TNH2WsWrZsOYqjoVDytVgVOA8pr9mSj/yZ3SkhO3iOFtXpmApjtGR0EVVICvt1zdX0YObRDPxxL
+tQZWYfDXkrvMcTlbmcr58x6U6WYJlVMmsJ8h3R6pXDxrQNNJxioPkDNDWyudQdsEp7AMr3DWr0g
TABrg54aoKBvLV2+5lO/z9nxQsBqs2Oylo9j32NgUDbJTfy9YUsbQi7Nyft+XT2DjsBQnFC91BCV
V0PwRvPLUJ7kIz0WcNo/frv3mY6i3HcR8iES11DFqwWfP2jhr7VLyAxhVJt+BV9UN0QVoaJSA51d
nQaxiUEANriVGIHH6iiFni+z4Gh8wVquBIx+M2uuSqta0FkyrjRNAL6kUnx84Y3il+4mQLOMvHAh
GhC7PrwCWJRZ9R9f+xUeiIqTWgkyDW3LkiGOedifcwaVkty9i5GxTNOw0xis+ymRSIriNmm8+yZR
hUrym2MpeadNt+Wkwh24Cov3bDHb1Rh4qV27jVAx/LG9r1ZRIrVnUg6c9nKppMIWIxHQnSFQmdJn
wYSZftMoTg8qynt/k2GY3JS1FnOvHLiRw0b3A3lPE8vKmNqrWsIVfrTij+LRavCGN3HhmQaQD0h2
ztqiAzALKHK7KCYOoJRTT4QdAFU7pfmx06J48njB0SZEw7Jq8UV7yRz/obY/Fr/C5LrDb1zDeRyy
MgAn6hslX3gmU/qINeoyNMwcW+A1V9g2WhXVuj5I2lXRfBcusk5L2IfhgrfEwtcGGpaychjAqVYf
up3Rb7iMFUIUNCrotq3U3ehzqtlTXOP8qmrfg7NL5dpIYR1vvTfkE751WfAinxEAoUS3Who7UqhK
/pVcXcLhbuDObaiYWtRMA0wXhhZf+vs4e/0fLNVUoWXU6XeBbMwfyxochDalz3sLVgH6qb0M76i2
H3f51NkJA+YjM/UXjiMg+WVUBGYynwoo57y2C+77OuTKhwvChFpnY+U8C4Ckttm6NbCGLFCzYDON
xxgKuwaZhRuS6hlAIZ4+ySImOB1dYyZA15M7aRzJhDUEBMzhiLGAEcn6z+kc0fy9TNL03eEpcFpB
UVZ6PAtx2hwhGVITVqOL8+S20k6Yb2Ke4p3R4XUq3qBgM/uKEOp9U02CIClg3ZXfVRPLd10SAlHT
TaufJ5p3yuSJnVUFapR1eeTK2bE3sUFCijPqJGbhBZh7OV+ayUzo8HBQ4HUI1TQrSMSdXwms206R
qJu6I/mTE7WM+9o2c+5bJGbx7tEXvtaBh+8DB6QGHcJodTh7rB8agEJEzDPsu3XZtTn4vTNF8dXa
kklGAz5/v0viQXjpE+tj65JDWU8zRSyJpqFSPnHdtfB6nXGBCdyykBo5IGegm5HSNdD5UFmxNk7n
gSWMR3ukDPcTDMna4XlmlCG6ogJpmR5RVMoiD3OHFu/myMEUYoWiGNta5IafzPB9/pEGk85PbQFn
pWC0LNp3vgJ04f11iTFyW6SHE+ot/sB0nHpvC6yx/O3M7NyuTTNb5MKNkMmIVVOD5/osWCWxSC0h
y6glOPIiGI1H1UHkJGMGGpr6mMX5WuZDgU0V++4jYRDFriJaw6vKLAzMSbDOUJq/UGrxFlCdHEk8
NwzxW5XTi4XtHaShVic2V3LiX3dxtQhJgKZgRkBNqXfR6bGl29jENMavmS3TEIC3QiDuWCaVh/Rh
cYg/J5yfwfblBg5rU7vDNs7KnU+qWXEQYx/owxE9bEu5U2TruGdrXF8BlxEKyVwGtafBNbk0tWdB
QcN1QXr0TNNN/o8kQszPJh06Sz/0jzpqaVniZkLKeAzLtqfau8xStnUP5PQMf9LM74kG8pSDxM6u
59Kvwuxqrm29V6NZHSVKwguQyBE7bcJMTDTrmTIrJ7o45vl42HNu6WUS2H+GPzX8LuBFyNauEf6N
a91WBMsNoNP0QaaInPWDkilxwZQGHY89ROORSfVHYRcI9BiJwqwrSUiSKfrV74FYn47BuOBZa9bj
1MhFQJILPTSTvMjKsladZOcOibCn7N5jbT2ylE11HvtfuYmTS716M0/3lufRZk9BXNP29nCW0Aro
hX1wXbRMBoiyyB7Ft+HYvFbCzINpOF5RjtlnlUWlSoDZbDhe2fAZqlr2WnCRSTzZJXwcU5ex/yfV
sLFMLKs9x1pL6+pJB/Ec2cCnhTAsMhxRTuZpgCrEixl+6MPFNeV8XkGHIeun3J1jx9Wm4YI9G1/V
kWcWC7aI2v7ocTHstBUgiovu8yGqxFSg07LzkesHJMo2mhgQP8qE/mZ9Hl6FSrjXMGwgh/rHXM/W
9w3RucdwQnD+btWMQcXEQDJccccRkW5ckmm0zUgn5mUi6nFu4P/dKeCCpx3LCziAtOH3vYi7hvGb
x+KURlo1R4gEVytkemEtFVCcnyKZccL82qM89ZsN7Ptx2eyJcMGmh96t++j4m3XyB7dFV2kYwmUM
/P+bUz1CSgXbLGSCeYR5bZRrG4StykdXnOnLjLg8KAJSbvJVnFYGit1+JvWaElLo98CIsImSDRHf
5GNk/r92XHfy0y70FA48SwUM3sqehlaCzug04TVcHC/iU3DfFz2UyA9VIg5vvb+OuGC3WQOnwIrJ
AXs5YrvGzWiozpukRoUXdz0YVkIwa7d8G+s59TNB2IcTRUCzNBT+C+61jZeviNAJYdSKAr40EDYh
g18vUeUlgxJbE5QifFrunTMW+is9/lVqdKfV4ljTq191JVml80vsxbHEHQruLoI1xLgLqy9UItLd
F+LLyRAV87E/pGEb5mIIEYoEQWe8TAF9m8R4bPL0LmwhDIr0HDbgDGZuo+xnZSX0Yev1TULD0vtA
B/oDhw48Wr9/XEklud8lrMdfeK2ue3Yqjg1hfQJq+LGZk4rmRVNRnShvStrDC0uS7iwQlqgABS4V
m59U79d2AQngJPxA6MjUhwmqRLx8ggk0o1CqD6zWYhKzxI2pDwcP3/7MyHFwaSiLyfyqaDVGr2kt
W4oEkn7do14z72SCtt2UKmoaCYS2jdIV7p4HA2eD5aEX7w2vyM0TFv2pQjp3U8Qi6MmUeGUSl+OL
GWnv2TJRKp/Y/C1V55FgMq3kLkENeQxfY/A3WXJkOSVZWUHGZpTTAOngECvN03JbpZ/HLwEsUx3J
3UKua4/ylPVC1JvaS+z7J98k70SBs9H9PVCOpAt8eoCDHOdfH14TrO8stEbLtrqxHvo5vrqYo+dY
sZNbxkvWLs1CNf5kn8UN6dJvCw6vPqjJ9MtXEzbcGVC8x8IMA+x70gqDQuCQOD9MYPsMb+DMBG3w
vEMdMcS+A4XeBlOpl3KgkXtosSiyAMZ0bVihiaKUN3yZYlm2hGVd4xlvQuL/mEgUmnLbfSRunqFk
wEHxpyGTjHQvr0zI7J2bD6cTLm2sRU+GbRmb6Jx8kZTHhSN0N1mrHJMB8GPjepL/lQXpEXXajNha
T1iVhI47dj/RQnvuj4s7CyXMZQLdWncGTmDeJpNQI3d4T03q1FQB3z1//8Bm/I/HqZRkLCX1Iy55
CCFlluuPwLpUI55hWNsLW7QPpZyilHGqdxlCJ5aJVwiKbGD1ru7+cMVpbwDtbYz4fRYHHQLPP5wa
KCMa4B3gfPDF/YKzQTk23YpM2Dkae4MYI2pT62AM4HIWTPSCLkU9kWOkEaQCKoJSKK4+1oI1/9lQ
rVZlatM1jJRdWu1jinNvpqw9jy5TJ3CwsT+U0LntjKsm1MfHnlILpVX0BDpOJfd7+aH3I937739r
V432stRT9DAzaoEn8ifWtzlVfIqwkj4LZQjv59R3daFIgyHuBVG65JkVbL8BdIsP9eI19rkJFieW
VTj4Ub4iWoJLP60hygkWIZf95WA3Li6AQKdo8FYg2CnkjSoGy1PwH/cxegpOg/A2gtI5Kebsq2um
ryvlJWgsuo1Dg/x1V0xJjBBvmcHWFgE5An8jIm/giECf/7ia/9iGHVegHC7hsgxJcyrl6umTTvf9
n0eCMhGz+cI/aeL6tTd3FYqK8XjAj0f3QFI15qL4om7Cs7EDD59V9dzHUUUWxTN9/4m6VLB0E7pm
YMv134yI/G1o0QmVB8jxDPspy0i561YGUTl/+/QEHjbDber81AF0n4oIRGK751gjcTOH32rAvEZA
/K9U3DfL3Uy4cMu0wiFzCe0OQi32jIhlITCCknXFZ1e2JHMuDnxpq8qX9DDz+DvFIcIHrmyvjqHq
I4igW3c78ZK7Ig6/TrtHWeZC0MAgmSQd8R4RDQSNUXC00cPn+TMlnAtfPuG8eYzZ/+0Eu9HvNzaH
W+o3t5xn0yO+fmpc7Bl65hh3td4x8V4nEDt4ts8zDcKdywWuvmxX7KQcszH0dmLxqXp+T9bzD2Wr
yOramam+d81DKzFASpsnwP9L1hoR8w26mH6W0I/0ycG7FIkyLOsSMr81+O2//1e9C0fvXdn16cgL
BesIuggIHXMipl0bcEMO9jGYVEabFYvP7OJpbDQ1nAE5gPK9za9xZ+54YWQ9gtAPXyrmG0aJh14d
i9PVmKwBumTXPAT6NGotvubKbOIozlZgthQaD1NADjnoqd2GKdYBADclJoTA/dpdmxpfFu/rAR3w
QblEjPY5TAXsNWpQVDnpfjw/L3kwnXqybfSzqM1AccNwRER5Ob49WFSflCPqUHGIg5BO3WGPyOap
K2HEUBQnsrzUttckNZj00OdXp/czYsRP+tqku/KqubFVMstYaClSXmIvQmhpjsVAEvEhWi4aW/Eg
ACpJR9Z5ZeibgBuI4Dn+JVf7O9gQcCyWSMaXhq7Accb3k8HwX1BzJ+aeRDRH0AFzqOB5592qa5m2
umojL5ELrf7i87vPcD1PK3VJ25bLF2+th8iv9GHaay+CoTQzRKidNuyiNmFjx240M9jtH7i4ojkD
1SGs3FbwnE5PMlf0ROAYk9TKhJ1/Go7ib/JxGapKobk4YW2FK/DZeYgwfCykfp0+nlgo+Rf3hLFg
tzCMnKuIWtN5suWWhAvVWQdDK2lyXBHdGNZ0Oz2PCPni5l1P886ksA8Hi8ti6i/NtGH+W+UUwe0S
uVvM7qIoUzh7snecWG59pKW+YvEw0cNPEVwmaxgI/Aw3vtcPhyZPN4rH/H4jRAQDb0c8H6Sro6gu
ifPjqqjXtIssYMVp3+FVt41HbmwFz9XhxV2TEDwDhIWrwF8C0CyBvR3ymUzCcANkdgnxEsYAq43E
e77+dVnHUZDaxwyDGJIzvNzICT5VLRIy0c4rNtjtSeZ9yYp6aiesJbRqAcb6fCEOTgSF6DCJV0sZ
PQ1kNzuEIA21IhGtrC1QzYrWWiAuvoGBy3/7r/KrK9o90oLauntsdn9gj31NhTHVZx4Y/Na6Dk+u
FEHPRrGdy1f+uvjblAq0wmPH+qaNlYpVpUMmVHpwhWyGXKKKW5Fbry1INuq6bw7paCQSJqXkMJYl
sbe2IJBhY42kGev7x5reECmB7Jq7bW5H1J7fGu+XKGduFhRlwzfe39pt6wsABYjWC5VZXQ5bgA7S
Ceh4YbX8ZJe9c+4Y8kF0zxQ7ra0beyTLcj4U7EY4c6nRfMUSHFf9zluOnnBtZk5mLEP9dOoZtgev
Hk+Pi0zCvSe+7QSruknUTjqATBupdN5aBCLVO3cfnZvgJ7RB3H8yO72br2dQnPENvv9QocLwqX7j
SzP9yMRfQm0ghuDiLcsCrBfjlPozSqYCt7bQuQZt0VYHG1WiJ+5TG+fp6OfRXT0JxiECZreL4Obv
kLvhnUIyGrFAVWxb/ApMifnnVod1cWQLTsEQVlhSJS1M18XTHSdWCZyZDoCbQD2qrIb2BULf8eUW
0/X3VcHEuu0kcZY/HtKc8grMGLQx7qoowJqDzFKuH6sxLVkm/oSV7pzLkwAX0G3bpSLvt38yEiBS
nneNHRkiDP4J3qi39NZCfAbElp47LKtbArdzCLFaDVFgtlYarP7GqVM7PWTG6s9rQePqSCUd3eqW
FXx4hLwk8Nqgh/nmDbk/b5MWo0SkmvBl/s8qIM8uBtpPH23dRfCrRaJ/dm0O5PYESec8RgQUuING
u/SmtnfPN6adYL2ThYCV+XBfnJma8CHFuJW8/Nu93RWIcRCl/TpPlfUjupzlGfozqlU7NI7tkGfP
ruWnDcCMTVaphjGZgaL+rfqIcg0M0ScAsvIH4exnxAKRYPTqeUmJgQ3FTGfvZ0vS2ZEqoFPNxSJg
RLCl3c0qAHYK0lOgDjPkD9maYqhCsTB/rz2gKilVSPZXmOA6LCMUuf8zXawcOoX0rc+z1yeywDxI
Tt7fZ/MWbReexkGdyGqw6pu+Hr0My1VW1PBXJ0jO5zXerDL/SwI72yoPMZSKXTlnmkNTYCGm7YdY
qrEYk3efDpy7cR+J0gPf1/e7urI8W5DZSryny32BwLFyY+s+d6p0Py6bdqwz3tjHtAFBOh4VEHQ1
B+Sp/MmzepG/wMynlU0IFglga8DmH2TPNBC0y65tuVqP9hItzI0DB1zn7k7AaD/LxhHnr99GDaug
vQMzdoIuOz3d8Ii7WCMo39tOUXBwNWTDq+Yur7L1fs+vy1dWjwI0a3rMOL3k/PeIkbcXcegK+sRP
FRnrCNWOm1uiDsQyrstHATkQIYPTVWZyhmkCW+NGNJro5itcHviItlN9q46WIxdJ+4IiDpds5Ukv
EG1dZpLr0GvpsgdjjsKjdDWrZtWBhrBJB2Isb7Ka8n7QWQrOPL616jnC0gbc4YfkaMlAV/nIwWz9
xifdzSAZeWEJTQKqE5daeqsXGkq98+wTN7BLobOSz5bDmB+kXc11k1D88ngQxpg0ZQn6U9FVbgoR
EFWXPoXqy/5vjjvzWT2jPzhn7kR/cKg8qolADT3dm+uWp6VFC7lStYPoKYyA51lptjuarAWnnCEw
7SpEj4bNVVwhTb80xMPO6deh4E1OByYYPrfgPQg7nrEMmAPMEG7D3LLLDOEJpcsmODmZhh3XmR9j
VsuqQAqs/zoqXqFlthVj9lMyPIW5jjqfIaTlj9Jy06nDr/G10jqRiQypKz+9MC9TiRNrqcmDWvPz
b8pu8KWrZ8aYdzkJHkzuKeFWxuBRYs8CMKff6tsUW1Nms7bI4uiF5/0VZQDHU+LBUpSxAubKGllD
m7t5OnfuodWA/UDJ3NB9ZRIA8d9Pe7ZzyGNJwzFrdoQ0e06RJ2VB4bZM+ApEFiySYGZk0EVpsX1l
UJGeZz7et1X/Qan9sW7d/WguhcTLegbXRlcjphyYcbnbKNQ96CiykX6lrgC1DdD1g70m2HroEPdI
wnzVBcVJZSim6R0tdmZzLo0wP6g2qQh7AXMcuWmfL2jM43fd5K7hse/MnKCupxyoW1XV1RAKDVky
2Lf4cILdnB9pDwaPHF1V3Zz4orBRmJH+bMyG50se/k+LiLqx3R4V38l3AjCQovfbG5fVwGqztl39
ouy6CZm6vUvwBsTtoL9nGhB7pmIF9ig5CpYfpnJ3wCUbCLXd5MTKcB856OdUB35RnP9ACDCNulao
teJkfDjEJ+TeLsZtwI+mocDaAvE6iC+T6pZdN214bKXzzZVo7MQttcblSpk0BckbFvU2GEzZ1yov
j+tY9FmThIsZQ+2GLviW96e2Gmi2ynNur+6Xi5GzGd5G/bxbk7ncrJdvAFLyPtCbjb+p3GPf+KNX
fVK42rEmf6DNWRGcOvUE9k2+jB9PQm/1l6+n/434YuRN8Wg56LbtBEQDMrS4704qxB4raP3Iwftg
+/aUrHAByDk+/8a0Zx819pf5767eRWqSno6TtK72gG030SOQ1gqApTk1xX6dImE4hhywPz2ybRg+
JDwcFxE4SEkBC9tvcmS3gS8x7CKY46vgf2757zHHKfbHophuF6OP63CkT+BSxJvBSFnziBpnu/3q
NPh5IV0R7Do2YRs7q8w2tVG3ZyuluFTL/daHD13EiJumMDAF5Cgm3Lf95Vl4ijQhRtQKtqUYEMeI
u8hVPA6y7MIySGclsJ1BzFnZ5fSgRLryqOuXP8YUMAGb6fk9lleYfEFtuE6HJcEtQa6P6iKNYeE0
51wAq0iIbjipv1Lop4OzIGeavAiK43tgrATPJNAMhmUQt/xZRGdVZzZDMjUgYhFqWTC7aJCxfKO/
2977LEBltolyDQv4V6U4ZG5sllPHRASkmPEAHwL4JYkOzWriEFWDDhXSJGXAmIJ99+X0D2m8xJzZ
XcfQILqTsnfhw6mhF7zZ2c/D06fEEjT65Nv62O9CusxQZMwDFdhxpJMwpHBfMKUDnOq0Mj8LUUS+
I7fpe05rd0GsVaGiDxOvCASW75ShpFZur22GnABp5DtuXsN4cED5b6vNfGTwtoSIGFZesH09pgqw
we/IzK1pD7cr68/vR6M5jljSPMS9ibndcHBZv5HT/DZiODtEHQxj9JiuYidb+Ag3oAu6kFmablkE
Ob21oZD7hj++YpGFMzEg/ji7Ch5cQioLMyaezmK98HPBTy3+1ryaUo881RzWdJNIl8XNFxspuqU1
uqKsJX1hCzhtrJHzslvqHFvPJ/HOMv/brTSBZCpZYiSOhEnZuudIbOFRPIpvcZ9x5HXzoV5mB8/9
kH6/W9D88G7ZSX1PXif89jEdUo2WGEk7uJNhHJ3EQstyLMo2njmygcDHbVbI87HqZzZph2f063Ju
jVnDiEHCfJq1DJ47WgF/brJDJR6zW+yS2qHkQHgFveXJagocsIZ4ovBF8ujNslWE3wJLQ+KZenFs
8SPfXP0hWUtYubAi5CgPNhgltS4EJ/cmpKxNDHyTNTfjbOMHucG+83ocAmTgUabq2fI73PyNAOEw
FSKxUKJYZusgepTRmuWO4Fvs0asdiBR8DuHE9LPCA4IM7+d0iDd8WIBSThcMI8pYbR3FSiZJimEx
/jA+NLKpjD4aNLeWq7qw1YY/pjwmJX6bfxmGNp/z2bkiD1wUErezod2YMxnoGum7KzZQXLlIcp+H
6KpE/cxph5I3q3flvymgO9/k9mXO2C8wtycCr/N5Qfe/52EriQpTEHFrRaAuswzoT1KN1hKQfSS/
P9xVai1uRlQZsqUVW6JxHzWoPiN9iLpnHUBPe9XNON/SuFY5RP8jz2youQGh4ZHGNuvGlydWz58s
0pO3N/JCdz4zN6BctioUTbWIyi1a4rI4vOfBgex49oW3e8jMIx7b0WXwmMZkmFvGrjzX0x4bnyvx
Q6VZKeKXMtugnzAjDvlzDghVxHDZ2n1Qnjq80HxOJRiUJGVTS6sXtoTJ1mtyrYUx+kpamS0aEvvz
Da9mkPivffvmZnd8W8Tum7q+xUnoY9O0QqkwwVKxUkgMmwCuJ2hnmZf8FeAdgAPFq3uoP9NGtMbh
uEMmcltyTgGdkG9owFQftWwI6dF5dCB0KnWtydIsEC9+9SMlMDlrmvqz1k2Fr1zteo9gUtq5Q8/Q
Q6zRi3qL9YMOpruuMu+qrGDEH7EnbSU1CL7EmkgqAgSlXHBaiu97hKeW3ezPXBMpPZMTqoNVy8sf
ypDQoO9W99JL43uE//TqyP3iM8cH3QJRXPSHgg3O8rvsKCyBn8RaVACrqNQJzBNr7ah90ge3dNTW
m2h2L76n/0lGKrhcmdAMwoPyF+oqsnG6icSmIwlPvsDnq7Mcon0dymLSYZ5KuwhcGmWBnk5ljtD5
y+6YkETzrs+wmIKrx471ORxpbIb9dlR/lYnKBxFq7FEcwCSgyy1eVGbEfJQf4xZrpCHSvmq9kuDs
mTCGT4UzDWzUEEju1kDAFSFUnoo5V2E/3ZEok3DED6I/ypukLXEYAg5GgVHwFvJK7qep4Uww1rf4
QT9cvZxVknYZ1yh3i/9UrRAeTYOiTQ1i1PLMiw2VnsJKWtxOAMfC++y/9toafShwxG2TdU/66DbC
N8fgv8FhrotZQ792gSvk1CEr6vjNSavxhE4Mr7HGcb4N1cLfE1FtDXsa/PrjaLWDr9iOHa62uig6
ETZWYW9hunDZbYJK8reOZKK8reI7khxSc00qXWVAY9cXRMMpo32qnxQaHRTECN7z0InFS4BK3rDQ
xrT9KuyQknuSqdHV7O8Q/BT81TkyF1gzvjk9aGZqajFVngi51BBCu1AxvMJyhRRe5abDyyCZyImq
QE/axDDysI1sCFdlq67rIfFbJy6eUdcEozkt1RN3V721UafZMnREcX9H/fEGfU4UUr/DFOCuX3QS
mGT9fdsMGsUzdf/Qu0hJf7BTor66Pf9m2fHAa2FfgxZQnKtAA60O3NmSbIODQw2OBA+LoG4tl6W8
9rM/QT+6VILBsw57sedGO03l30RtbwuTN1QW4DXlfZ/C955hR+1EbrGQWUaQzvDt+aA2gJPDEoPD
FfkmAuEJ41GVEsMKPqILl++lQATdvjZ9M2aj8135W0F5tdxxoobUSmYYvIBmuiPjohfsCDM+cegi
Ip5pPSR5NJXeGiPvPNBtxuCiYFmzLH3qH8aX4/xqxheMT0kcn6iT57P1ujutr02uCLsR0lHdDhi3
wPv5/XrDF7mZqCEsyR3AnyiYTByZGWGxzaYd8OIzAVyJVm7aX/Y+EmA8dCNaej/W60jrTRdlPncV
9z/X2bwI6RS52Og53VNX8xoyWLxrQaJutoWt4w6pfDf4MipvCwRer2/wHNpOQbwf48B1lxjEsEo6
C8wkOlSbBYwmlzjIEENeIjEauiPXKhGuMnFkaVNvVv+lL2GcRkl+nz0a9h3UJqapmY8edJ08QBA7
orV/vPn5NQ3KOUxi8YX/WAEg3BXVXvsnSjOk5iEOKoca7lqFKEvEZC2+ySMX1S0xbTXenM+aNXwl
avXAJ6HFzq3UFCW947eIySN2qdmhTC7twSSHTEHeLUNycqOuSz12eZbAjMaw+x/eTWfvQRUjvHfM
daCMCtXgYFn6G7AJME5L7E8tRJxShZh8QFxoeEu2CMEZaDcNDepby5oNjqArXLPYagQtihWmJh6N
BtgcpGzBKBvb7Li7U/1jk+s83QRIqiJK614cNvTYj9TP6uMsx9aBMGggfJcjO0Nm20Bl70izVeC7
gEfdlcDp4siH3SOxD41aesdi++/QM8FW8zCldu+QZzogCSKvI0wXAifFOsOmOlgBRVK3v8AYG9r3
MAQHAgCO2sUz8555sXIfUzMI9HejOu/3cBYo5UN2zYxljvZP0o8alRQX8yA3R2T6fveHDG7VufkC
ClMDlo8v1YKXw5Rap5J8bYhDV5Z3pPrFhu82O5KcRDhO0wexiziByAbLFHz0oyCG5kDr69oyXEtf
gRVYqpiFi8rJpIAj/pCoflD6CnPpObJl1vjyj6h0kCAZfTihrZW+/T02NBzk0PsYSzkgEjaYg8Pt
g+kvXVRusLZS0uytdUzNWWoV4LlnTQOcitRuDVMl+MgEWlZe3Y07cjSs1kdaxLmwiTDDZX6eynvw
xzurr1/Fqasxz6v8h8hmdQ4UyXTtGAg1qiBygknfH/vpBC7qUWE7osiZsgrmQYboepX6VkA6gWc1
Shfqz0UnkG4DzHMcxGzTrYaXHuggQjqDNV07EmQYSAYu5cbA22ZGxUcbZaGAHIr9P1Xw1OjFBHX8
yr7OO3AyTkh20sHXvHymTPynuRjlncABsQrnij27DVvJ2MAq4fpKZXxg8aaCQduW1xBtWsgqC75C
xaxIZxEGvvKVvaK1/gaFqe5Fg4XYuu8KcdoiSoy+RBohA9I560LXP4VXfHUHTI7v1pKbUDaiLEgz
jB9NkwQnFhL5Hrd/ZBSfCYl0Vg87wJYi+3MNQYVMsOTF7kYnedIPQH5FQRBvVZv6NGwF1BjBgYa7
g4R3DS+5rvz/W+c8ntskZNy+hoSnEa3gWK4HcYa4vmJ+0HnfYUYTl8C/GoXG+B1Z8YQScqVcFjUW
UWhXDBj0mbkcD3Yk5ZkpsN4+t0kS2CyldGUNhhzBkfx7Gsi0QzZVv9MrafMc4EAqFVTIhambfWDF
W447OC8NOnJC4Qt9gazqc9Gri8ct8XvM1+yRTF80tcwrXxbGJ+rfzG6pIz6NsIyEhtIFbsj3yq7x
CLH4tRaHxW3wKmu1V4Uw0RYtURU3wlpgfyrgovusmzr1PFfuOp+XyCg44ykdRcgyJxv/fivIS7jm
eulGmTxpaHhLkfAVaDF6PfqoaVJVPk11s9k9E8E1fMAhLzpIQiMBLjI3sX9Fq0QOaGnzy4yK3F+S
fQ00aZ01+PYNomrQohGi1yqtM6MYPDpycvis/d42oVQslUL7hCBOlC37Qxa1S+4y5jWH1+yRPRsz
iOnHajKa2c7faC4+zVaq4h7NIm/ju8u1MWuQDaPbsIo+8Wd1afefzjkcP1a0ac1d11o9ME7bcF1z
zbWGigFyp8jh5DSJ4lPvX/MS+X5uhujOhXbmAsFhrIpVd6b4dzb0wenM4QriGShkM63O84XZdI5U
03Fm3Qvvn0slydkCD70MKIYTlwe14qenPC3iKJh4Qw+Dvm0123Iq+UBEqY1cwO+qHrRaHoYblwrG
jaNfAXzlgphevCPJWf/4NJOCebgSz9/OEdXKHs92VpU7TSnXE+ekLpFxu7dkWe6RJhtb0DlIz5+S
GmLLRGN5DskCoG/pUYERZxN7UwDuyFb+sPXLAtrsJr5ARRJf45ZSxQXIswjjP7hiTGJGLQ38N9xO
vZhGj/zgcrhHkv8Rdvh+2gb18tMwcmgC7HjYezsm3fUFZ5hz1spgk5f0UtX/i9MctNDwkWtFW64w
cIeoVTypUGg0oh9oLSB+4/tj/cUi+aX1j96Jcr/8pRb4tnJ4X0OU3DHLIvWBoCGOU/Isnjnkavcn
1hU1nw1M26hSK0WD8YXSr0cb6zruaJVdXWXjmVs/gsY7FUQynw2anjsBF+XWM41ekE1UeSlaXdUs
TagFc5PiYOCNkLf+W/uEHP3v8k5ViQh7grUL9UHe5d0UE7+WC5vxRHaAyLOB+qNkE9e9wPSjfiW6
9u/GXvebvKKVyB1FKS7I3QcDRt6+og3RMSQ/3t16cHNgEh+bTQAAjzbVi4goNaIKd6l6yEEzTCUQ
ZcR0pMj9dRY+WLZuEDnnLbtZwPcW1CraiGDYtKbkc6FtU2GDpTNMqfTbnKhd016yJ8rs6vRMjKte
qX5I5c2yZ6M7Gg775WpPUQHA8VVmxt49vhwlA46J/+ZH7ZDc7Auh0j881Zkm0kff1O33E0SnM8uG
jUONTQZR1F3b5knyG2dBP3TV+rH7oRVqa8X24o75/dFQZfOUUZaWjxFVBi3tMKS0JazR2J1xOmWt
BCEuUSHQVJLVwJmFnZ5NMLbzernzfxt2C+jUKIHBUwcAxl/WQz3hK4GBLBMpmaaz0YwfQDAhaSTH
QKchLYfIVlBehrki54s9IePM0hqkVLC3RUkoobMUx12hS+VW0Y+iOG40ejHOcSHSUOQWCGLUxeiT
g5ZfApwMF7lm2sDKRD8zKWEUZ2RNuc7NAAsutC57E5as/dmk5XaBTPPuxueIPSBiA5ay8ALPIOAV
RG19OleJzEfRXmMThC5nd5hoTKMsJtr6xKgmBJIDYB44dp70D+rXvyRLdBMdaJYFrj2hkDpXcT+m
iZPVZu6JlZXAoaN7Hq2mB4q6DqeKEdYC+jOCghX3zpdw8YgIx2v1HN5XeAz4d/vY07i18KWZyxAX
EJKpj9D+ymhwy3eGaghjQg7TcSQXu4T5BrLTkeh43wwCRBBV70Qyz0Sz0zVKzD5n/mhs3Ddr1h9J
1BHXaoLgtFgYOv3qNoYKTUcbhELotP3RM/PDlcNt+9jpHfKH8uVcCyVi3y0hzMsw4gMsy+iPKaW8
s8lF5dyK7dyaV2E2nnwoe3r1CwzqC+dlX3U94HzCSt28u3G01a9IsQHR8DQrXF58xpsbVNrWehGx
F8XEiY35kYx0pYNdyAK3eJv91Xs4Tmk0ThFMNjKEXCghNJ36jZsrU0xa4bL+NaHygVog5cGoQWr1
40qgu+KIEFfMJn9p96qJVwASVKirnG0KNJLUNrNVt/irA5OeTgBdHIGIDYgv0ej9RyGfWjMKwRuh
lxSFrg623PLvHpLXzkZNuiqszBlRPAEZuR8bD7H8Xyhwoemiov6afTSNWveBhip9KVD3fvRut25M
C+718GQu8USDmNYbGA1G3iRvPZJ9t7in5JjXRK7QeBDvA1+UgU3d+qEk98DHsS5EeyzB2+0WTqJw
xWK2NzmZqbtB6LQ67BfqDwJpw9/n+QI2TXwbzItA+OaIfPG/u2nRldIfYX8TwxTRHUL4VFpIlAA7
EHKTWAB54Jokov7NhfVW6NhbFlBBglnaTmtOQ6YlZg78XytEF9dM/LL4JZOM/+84G0zLaMv6PBZM
LPJ10xvclFbYnrKRVMW5QA6+ewCYSgeToR4ssNt35x8y5XtfP5j2LbgAz2jtipNH533dYyamloyh
wW4gylelkd32PsTxwqr6cMHS0LhLfgpHCrFo+zriUBM9x5CkKpe2XPD/LT4MC5WDc9ud5RKid5tO
jLXkEjHZyqj894F31MKCC2J1VmZ92QaTKHdxE6aOiez2yjFrldTiq+QegtuGEysVExOqJ219AUXk
xhiftzKrkebkdaGTP8s+KyE0cfOn0YsA4TtcYob1GsWDVDIGVjet4HXflOfIXE+EvUs7SIIGpOV0
8XVW1Jhw+6jgH/kDw0IYTLWGQHnyE0qwVejg6D/c7JJD0kQswNNW4wOlG4nqJt6ZRCFmKytbqN4F
DjD5AyFSP7qLvO8QP4pOZPixOt8jCdG7yprrbKpX0PgJQbQMHNmc2OeMEgRtgukfs3o6kr9jRLhy
u/hr/N9hm05HCJe8LatwWwZpHCtHd+dUK+XlKWKz61ADg++4yyiKJHvIXnrKgLGhpIa1Gi7RaLZg
Wgh0RGwcsBIv7KtuEfMuN2dUJJz0ChVcx5S9QDkU2X+ftQYspWkiE9rfPKZsqAdRTfwa3kjkSj+F
wksnni3fCRtR7y5M+JvM0hMiBzW9//bWqIqmKZXpt5uE6o6fMeNP6rf+4TVXDq7Fmy9gbF2x8nQV
/93xoDMlTG6FqvmQm29kPbuIHSY/0zAVmip22kij7CbYGiRpV14Be24tyge1GNRpdC/8j8a5ebJB
3gHf+F10sa8oNouXnfTWjZp228i2Im5lmxtUPMDX2JpC4y4IhO5pcAtek6b3/6zKC6FPs1govSNn
8NSkYl16jheTOuPg8MEKdF4F8h9adh0odhEuZ8mUkaORowtJyAzasWvREgzf2OUcXD+PtZnSYezW
EFhAXsUtwRSGsi8xfBBOE+MOm74EOYwEw/mRZAoQvlf0NFEkweTLqaPbphAcY4fpqOT/LoVOMERK
MM2dGw7+UmfIHJmAB9JKiNlICU7OV6Gk7kXnuJED8SSa4rW+wY5Au58evwDVrkTRflsb4JxfdDL3
BjYWO05F7TcyBKJhKylxXD6caZ0+vk/QUXuGzXDeltEvVDuF50ZAOYqeyvrG3ojZIGxjs04Iidyg
TyMZ2QHLDCQqCUn5/qErW9o/bSNSYYSssLPeAAw/0voSPiM1ts3lcwxGAvERYDHooBDyO6xb6O9/
wKi4BDQ9a3T+OlvNufuTskwun0Ccyu7h2d9N+YYoJCZiJRAp05Fb+pcx1IfTbk2A0wlHu5XVNN7z
48GPi6MK+hFUx0MUEV4OH33CaugyTav0TFH3zNlos5qI/trYUQzjx575oH7yIveGgfYaOIvBNcH5
ibBTHg7SmT9uuE813rpbQrg+XLPgZGgFS39SctEVu+GG5+dR2LIXHBv4uQkHDg7UclqiZVEHgQ0d
teOdZ1ReJDPB2mxIFL6y1peBjJaadE70+V/H8fdqnlrsQUUMEF3HBcKLlJJBBcJNjOeFyRUEWtxG
0V0vusBZd7wqA2pboAKMExRSm2cuxduzrHT7sO4teGVBFMnbJqatzEc3OPnbjsmYsWMx2shL9alS
nf0jSxtSNhiy1B8Ikc+q0HQji5yt+6UDlSL56QlxiPmHBUgYXmwpppPNDY39cUOzuv2vWkqyahYS
BK0EMivW0jN2I6x4w9UYa2O3R/DNTleKhvAbN9PH/gQjMgXKUm9cLPDBE7DTvlZDAZt1ljTsj/Px
9pvEV4iwqDLSEtHhH7ExHbHcZhxRBax/2+d4FzwULlSFbaHjdhEvj+HUf7kPdLLU+52U74eM5n6X
ZgufI2ugFi7E8f6xgKKrAJ/N9FWyB7CGWqvpPz/BTwGQyOC1D6ZWhJy084WUUakA98TFYDUCSooc
W+0+n4kJXgX3rHBajpoy3WFcQrCU3788d2btBAvfl2Tui5qlhQL8FB3jjlrcfQzPwnyXUyQBYpCD
PhrGUHnoThn9tgrtOAaEMzy+QToVZo9vVTIOpgG/eohNjDPHRWk3Rz4a5YhxBxOOgXzXC2aMy/JS
8gWk3gMRkfMZOHPTb3IvwN2PJ+6pVsI5ffrt526zybeJgYi43cR6Mav598tlCyBT4Ul4FURbElim
tAFD30VWjwTNksmheQWiCvMwn3eBJKMMDAYtL4LO8Uv4uMublWFqasOSWL1ol2ai8mCeWhB+aRhv
vRtQUDHqGwOwzFgpoGG14Yf9mk4E5M6BopNRQ35LOC3z9cw6eGaXTkDF3aNi5eRdZu3hkoJ7ICXC
MjxM5mbE4ZPXOWqidDFJmKCRhutVkiEWOhKQd5YcalAsxVluvNHQXPsU2PpjGgDmtRT8BPBo/mDH
VDwoUL8EtXQQhnKqXPc0NFV1/pkMymOi8pQhMSZcYMHkVPcCXozLWYRQy657Z+5OKWUYnRaMToHE
b0nGKpwGGTmfK0eBQMuUm/ageQSyEKQhZ/3IIN5rRD638i46X9X7Z7RMJTgc9Ydr9dOFoUYuXAhv
Qcr/LtTY8Fm0QRerHTSkGUJJaxMWBnnWjPQ+mQ6jTYIaC0s36p7OXpFoqu64vebSmM6/zZJsw1VM
p2QSaCFvwDh/7me3rzh5zUJA4osq/1Wjd8ijyhfyepjMTIk+RrvGvlyFW8/cdwzT6y4VRgCTXl56
34hXGYdOyxWDMx3sTspaL/OosXf7H8HoBTf8ahY9dxaAthxpmn1ktIX84rg6iUDYZD7AkDnE/oMD
RRpiXjVtn9FDtl2UCTKl33Pp42QkcuRCoefpjUHV8C5U1AwjMGR7yUMKUOI2WTfswzBiOAMQhx7p
dbJF3h4m0E/J37i4UVnEfug3T0j4t4Lb+T1TDNxbjXv2YPhksFBqzGzJsmVx4A/KsEhFN70raoXk
yt8x7AWDocyOkxoGQhoJSe9MB30DBMybpxpHgHeAH+AKFptx5TmvHmZW4hTy9wrd1BJ7lOKJ4FTS
M1ONQ9GhD8wK7ItSjF21Hb3ZhOcxiN4Zt0EiImrVU2m5Il7EbrQsHMBOmYB1vfhoRL16KGjlKzub
bjFgkdZQArw8usiniYbBmLh/HJdx1sSC/8bTPxKsMGP0SkKNhEd6p5dgwKN5X0/xwpkbV/ud/KYN
dJYw36xQ/0mBO0IwuvZ6t5iymB/YNt38bv+4KF1VMCHdNMQXC3RAYuru4pkdjPFoUpCd6Mt0nLkd
5/PZ2kVuvxcFGG8FKOOHXFtIEZsE9owQtWgsaAinTUAU806uxricaIVKbxf92+1ulU2JC9MaYEWG
3T8ulf4JEFkfKuzQ1Cfm8DgBhUdceXX6sRRwMZdLLE+L6ZPw1LqSmjPs9izWNVATeyvyJYnk1Zsz
rMfLZCrMtAE6O90zc3vJUCubC99uuAhP6E/wRsNN3bLzuWGpQWsbtsgJi3hwUrdKW58iAnkgprSc
a4RiOFNCr412eA7qcVi6yuIWb8lspKD1bdQuWNiG1ATPtYmLgjLfKls/R+pUMOZ2Xo9IfpgmOD8j
HG/QM2w/965tJgGOFbmO3O/Ip9f6GO0ns1MrPZVHjJq9CFCtyOAuMpBKoZP5ahGm1HLQgsh5wAS6
H1NZKtuwuo9Fu7dbS33PvxxCzgZ5D1Xj0vpDVQ2+YOXR/LI2I/dCTTccPqGkT56NlLwK05neZFg4
wElN2K5fGKarZ5SZX+8Gdh5eBSNBE830825MziA+5f0XyFDGKij1YttbIjdhUoVYwkom0/6bpOpA
SuZuCWWVwKC8g1d0lLnvrjpwtzr1bPxFaFPcZb4WdsrVxKQpe/mpT5/WAejD+I3557XU7KIAJBtZ
uhL4jMeQrHH7iII8JnN42rsZ0pqa9Q5CRChhgoTvHdEQ8EtE4uNfpf2Se5w4oCR+FvAVO/A5jdfP
8iKWFZyhjdFSO+L+o8d4BT2BtwhBGtswA/pUIoDemEFgrq2HYiIBagZ4S84bd2a1Fiy58fCLMvL8
B/W4ky9PXGE9mY7TwoRAHfLSncHAIHgWcC1ow3AqcpPmKoQbaMbaIIXHzKcCopqPYt3O9gqYZhhf
HasCKJR4BX9tt7psgDyxP4WnNDvIE1Sz4UALRKuagiQlRDT8SEamKphDJ1Sk3oH9y3lH5nO0SW+W
nAz9FKLHlDVHMBl/HxcTB3p58UH3TtGnZBKvJolDa1EJhOKJg6lwY4aDGy3kxtKcZo71YjS6mxpT
NHJ37GdgS6/qOHi2H0g+1dwkmU8F6BDKKMfTamv2D9QDZv8HsDxT43sRZyd7GdSbDZDYVRW4lQSz
x825pRCyhjpJ+3DqMjDjffv7Oi9Y1zShvVt/sa7y8x2A5Uvi8vKih2S/55f5pGNh/sIyGoqSeIwu
1BqcM6CeDT3g4BZoOdQdJX06eQy68WBS7pEOag8fYA5CrlmK11boaQcrP+lSkbTrSXeBrf0YGE8s
lWTtaJZ0oqopgIQK16u3r7ljcHOdslNCn7FY/6qDldizAiMyLV+vef1TKwPWz9mGjs8fQS7S6L/0
vd0N1mUptj6rDknjju64CGoKNFh4bNLBInbZbcpVcARglb01SwlE13ITCTPGbf8CwlWkFUiS6lKZ
pgE2htmYF3coSaA6OpsiQ4keBT1t9BH4DhPoy8DZopV7T2BXiBeasM75lQvBMH0g9OFofZndycAh
xAxMfqF1+7OGzlHfCcTzinog4yGAQ6Hj7kWXJuwTCOysw4EwN3In5DaSkjV2Oj4EakIrRE3o0FlW
Re6gDcxZErLYJpvo/eLhPn7LbSJ902NP/2wTSc9O1O4IUAxbJ3kQ893q1hq7jzZCg2WL/MnGDLBz
KQRpBlTBmg2gr/je6RZHpBLSLFvxzE2590fB8LDFWRPIDqe0V8Zt0giMIkU4CFk7Yi5JrmKtUDPJ
BD0uZFE+P5R+W946OfxwcOYmq+HUtMKyr+cs/kDw1DmP3ZdRV4oDUyVoRDKIukzRT2M77i0/lmFG
jyEZVrAWQ9uF+UrS9gi1uC8YsLTqfR1gxwnrfLSbVRsksLe+DROLwQxXUr9UC1oNaM19srepEK7l
UCXDD4OEUcmAsPa9KyayfUhAVEulyYn+vKLWdO8rfq9y1QFeXEvEnGGwKuvHh5s8bWYEF1lfbdb+
3xc1XKGh2Nz+/oY7/heEhQ53ppKHyBcmHvJuqqOzupoJt4nH23o+a0xyKs+3trDSZYVL9uNbY2zO
cbrH6RtDO9chUDX4DP8EA/7rqFSGPe878oHPTO/zzhhq7syKgbK6f8OynRrNePXlKU3b4pH6TPG1
h0BMG8L/IIUc/0Q1Y9UuQ3Shw+52Cmxwhann41PsQDbNKUtDeF54AYQ/Q/ybP1wdxKepi0TcSi4S
ZxiYh7x6Wvd2Tg+HMS5HINqex27HH8U/pfyg4d73IhbxYLdyv4rrZeeBMKMR42mau5VGQc44s84k
eNJIV01BtRl+n3a38wwPLfEb0K5IFxPfF8MU6Z42lOZb9Kc3y0XCQoVe/GpvxMxx0P+26kM58cA8
Iezvpbh1Yr9RwBJAwK9LUr6IvS5SSS4D0Ijx5zi5Bk4ZD9BSwXbHK+o20lE97Q+949PDnpQtnGgb
cvlprKZ8Qm3XIXZYPA3sHLjCYoxeXlWw757Wz8WNvRSZXhqMjKqSa/FyDS2UV66q+p+EDgMRFcnM
XyDRwev1Cs6flBhJ2BS2HQ9I/VXlbmCXb2GXD1Wl1OMNCW6pBy/f1VXl6qic55RaMDGvuvRUGj2J
tYxXywdTl3mjBWMrwxkaScE+M9Y7YyQxlo4D2YioOECU5XXjmbIZD9fR3wjJ3pOjhgjCkT8tj9ku
X62QkhK5lbNd+zq10lTTM5DpXu7zjh6Wv5iEfB9iFfU7srHmN9XwaU1rzz4IewqLRcgVasKKyyuv
L48CkJVc929Sfi3asoJtUHV8LbmyRVW9MRXVHNbiQO0geQxvHPiKKRJJ3oDuwlv/Ruz+NP6qSkoR
W3ySgVuKpmRc0iXZdUCB7Zc0MgMjR4Xv4zpdIrCNKa3c1ons40AnVLc7BX5x/GlH5jDXWtUDb7Gy
KxBzYt/uYaZvaL4A8wQr+3tai9mjrGU8IqdOAkBsjTi56gEI7vpbBYYd42rdQ9uszEJZ4O2kuUHD
oxWJYGmqGHfu9TL63qGSGEhANDItvZgV/ncOXKLzIMqChCaepozmGcZ7d3vw7I/xy40+43GKAoQ8
qNv00MJIlkH489cJKIRyY3CTt78nNJ6NPjM95AT0SkXEMyMlbiHdmJ3xeBf39b5/wFn1m2MR2x1f
bYrePGV+dzqya7RAO1ERCFMZa3IFYef6hc5uP+H6OU6yaNfmB4Ijnck4XVxY5QitoLYqeIz8jT7f
8q55W32FS5RKEIgY/L2HaYswVMkrUi7+VQYbjWVcdFZ2o5ElawzwuoCqn90jJKWutitXxdqS/ORg
KYsDlqquLMzKAi/sTNNXQ/NqZ4aRfdZHTJ/GZyg5cF08177XTTbrDB1suARjGCVU1Z2OrTSWJhVr
GPK0XslKw0q8CHkg6Kl8h2UMkJ5WCl/mWkMqIxMWVH/OeE591lYfUKaUbZk3XIlT0sUbOgrh4aHw
dWAac3XulMmezqIMyfgujI0gdqHwjiz80yauckYdSKywHPSIJdpyDgQ3C9ipz5Z6/9K+nJ7vS53w
GDvgu+2ys61DSnixUchz+ivMzYUV/etOPCYOMFMhWviaIyvoiVkERbJneHP66uPf38ona0grCGJ9
VcxAxjS4c75YH6Z2TuAZlW1gMejnQpMl2/alavml8ofqKmKn7/Yuux1Z8R3aOgFpOCUFQvC4y25A
/yV56PiG3xGy8jY3LswqaEGY9VQQjilt65o4vbjuahGVlwzzeKxYTFXeCqitQSzT5wYx0itYvPCp
i5C4YspkkrQNL9JLM8/X+a33upPK1GQMUz7JAtjNuhUM+B+IUG1BGkFDfsRRbeU+D3gQ6DOnCCeg
YClDFnH167GR0B0BKSZg3fkIB889XHPcZHL1M/dLYgaLHIrPPT5VNFvzrsm+rDilE6ZpfPhDPjQo
avnFh51HUC8WsoIiQszzbTuIQAxa003ZZ4QY8VnaSrU6juo1p/9/XMkAuNTLCxeBk5lpOCIbaicM
yZFu4c6UYnTa4N1f8rJTVxWPhnY9MBTpOU8P4VrYxUfqR6m6GpNF1Lf6JCkRutrSPu0KMox+DaM/
SKR976NJdGYTUhVaLDW/koC2PNWHYH8F5rJ3pGdQN1h5poRrDuc6Ll8DfHtc6UL/Moebbwezcugk
kDoMOo0kXvliQ2pnsKIH54Zg9rZ6NOkzt/VQjjsHGlFwCDlOhT2UYuo1iQ2Vb5EFCw/EUOCUKSj7
3/f7qVwbzsd3O/Z/YDxo2AXb+P56fS+Z4g3XPrk5VP4MHsrlj2KvFgrV/eZbFW1mUXDuqPoiO4/6
WqvnnGNNh1mq4535mCuNz0BTi6OCq9uJOjs1FsXlL3mHvzUY+0r2rWTbF09DBMdSHYJBXD+1bitl
/4ITm13fTGl8XLlsMBoZrHqXzdhIybyzpM8rYFxfuJAX7t0O8Tp024VPEu2L54aH35KpRzQGzuuy
1TshylE0PdEMD0WQns5XjD8rJ0pnRYssvswSfyjdu7MTqxN9oKPTBYuGXEzpnzZSqymwBBxuybrD
8KGTOx3LvoahAldbuKVzpmNaJh1085K/6yY5TIE+I7oeidrje3QQ+Xm6aigB0Dxm92gYo9Ks/TNY
bIFMelImraVByUv7dprtdfO3c7fgq/0sGoFyNBScnVv/Y2Bz65XNJ7vUhw6QJmSQZJrMdot1ySbp
iKXaRbe32B9VdLg16Ud0JK7wdqdA283uBab6IM/uRgDljx2x6uQywfdph+Hi8xb/tbwEwoPT+8VM
XuDomn+nxXSjumv1kY7Y8VEUl2DuWAkq8UNY28vdU4iofxJoDXge89y0OKVGbXluxiX82Q3EK0Ue
4/oL2JSLzQ/lPI1QmBsvryClFoj1qrXW6aZqyWiNjaZUBj/LuvSekvUxtkfXJm7lj1/IhinZOXCE
Q1HXz1SWySvii+HzUA8jr7PbwV9EIsq5lgRBkUDw5/C2ZV5vvN0sBlqpXvV/qWQfXMbuyrDkDKyk
QV6ad5aDxo9EMQifcNP4yEK+nDFaqdbT38V0e53qhQsTK+GNfTeBfxvh3Eh3dVaT7257vdrgrWDR
X8BpjA9dGrjC80N1hcAZPUOIf5N/mIxE17K1VQiV0TEyxZ+WPZLwBa6ZxGSVnDQFfC8aGQjgWA34
zvwYAfISMBPe7uxdQpw0g/F2RB1S4R+t95q8Mwg22lnlbitTzcfldk9LrtN9/xv5AWX/q0UHjWy3
2ni6j8ilv734eXs3bvEYBW4LsGG0NnSbxYC28JMmLgEajpjaVgftacm5QGD7uvCIrUT5zd/I7DGW
XHUeX/S2CXQf344MOfBR1SrE4oI40NI0QrTqrQmg7u4qrly5NthM7k7jzaTLMAR7ezxuzIfcqOjK
AZjQiiAl6kFcwXLYmF2+2GKy6CilFSKERK6W3Ahrpg0y+BNec8oRmq/4soUcM7XfOwRkHVzGy+XO
wT7EnFMsjpeBaauk8gtoboqzr3lC2U34Mla6Vepdaq7PQH4KvmzfV1Bw4Yvn5ZFUQpEZ3bKxiszX
aW/A7mXl1OzapNYAkpZ45PNm13Y1MQMJrPHOtDgNQ5UhW8kBknCo5CcDcx2oL2ZkDrWZLL+VNKJe
2ptH2bXeKCS836juBBZ3ePea8JMtAPI4kuJphFLfHdANZGs7cvJ924dIIfg3/oqrb+oSZC/GJlC/
h/qubVNSLCZvfTRrSTainQocKNf4EN4suQHuZlCuymWKuoZziJYxXqcPdSJ7IFTU146LdAAzT/8r
IwwmiT/ScssvXYUPL8AvbUxKbQpraNVvFwcbAMcwsXh1o+1Hta8cJ8AmN+mDhbQNpKZxq4UsJGlL
55Kbtff+fq2xV86slTHlJJyer56OBI8SrsXvF+6cpQHXZBHo5yru9uAj32kvgXKhZYJggHCWiKG3
ukn6t7Jf7pMyxRwehW9KIf1Dcz2RCvHo9Gd9YHtmtQQx/qqEg3MTJZO9fa0gyEnUqCbZSHaw/3LF
C65UCfbvccfJX0TUa5nJS4+rPQV+q6JZhex9OmfgnW637jRG95HpWN4bjEKeDdQ8gOqlQa7llUs1
AOS9KI6EIyX8FjUWDoOzKmP53QX1dApBkfPXUYWM0tcG6Nq8dJpfbq9BnVJi8XO7f/VHgtyKpeWT
gp7RIQEsjVQoPQQWrtIBshC9ZcWPiik+GyoCFqkxz3Fw33ds3EC8Tj+/LnL6StI8U6q3X1ITYNUT
eCGyiyF6Hdhf2pErNGi60aHY30xYM16Ov+IBcswMpR6VUvhQV+IYkZwkIbE0OTyEYfaFtYAQH0P+
68d3+UnVSAHlk3+/IJj7JR48ojVL8i3Jqm/KwDSdpJTNjQT3a/KZ6RmK3QFHarcXOxHoIXp071Lj
zl7kj5x1jxndTNKgHJklBov7dDN8QfNfuVaoJc5kHdoSROJojFphpaIOdbRQZgH8SdFDo9Yt0MQn
sZKCTqqS2K03HZkZver3XL3twVfwL11YOjJX4vJpa4yXwieagsIPKRoAFcGxJ4Qr8hhd1R2tNbt9
a7SfBsCoNGnx2xVyJxMLhAXl8Ex6Ew61w97UTMRoQnz6JnCKun+iMxL5Fo+49C9wmVMhNqGNodnQ
FaPaQ2otk/EZqLdfYij+XnPnie7Q7aMT+A1mP+8gBIiKkTJAXP0r9RJi5WW9sy8LLIyMMaz2ynXk
6D0Fddrfugk/SRwcGTjLGrj3mxCLhg7uP30KyMHtG+noxwanxcS8MSnpwBeUIAM5xZSwyd4vL6gL
F19ezrMRkR1wNq6ediiiuxLJLU4ZWgFfg9XbH0g98kU7ZYtBPVkMp6py/1A4ZWM6VjO614rNB1qF
Ytx2atlJAsvTiK2sl8NKnIH0dOYQnvRA6K8KYFk33wXEeZeT+DE30BKMbKanH6oH0InsDX1BsokF
cqDP2ZMhcSN/sHYPfcoCIvEnYfFm6M0v+A9MiuAU4riR92tkC+S/3nARHgNTj9EbyqqQO/+CXqpl
bLIKUcFM60jgHEOpLZniRyOYVjRR7w+odvBXqZxWVABd15Ubcqj/6hZo8OraWiMHgqU1ft0CbhAj
Sx6WhRrgfCteaIxvVY4f3XouHNKK5jTKygCTKdjkX7096GYCvImXeqWyoLzlpNHYJLn7Md2h//2o
CbpHDBLGMaoWbprMhe3vBMzY+6vciWlcH8ZzFNviCIwfgdc/fH00xhBwBJYX0kL+He8K7DJ126ds
4Pf0GIfTvkXZ21p6RmcFlcE+H+CHHjrfqGaiiS/2ufyigH8eMt0hWe6NcPK4D1bT+XQDqQjm/UAU
xLETv8ERhm2KhHzJWWRrp52qIv4WoMcM7JpCXQWtYMg0jq9gvEjFQLY7E6HlHbq7J74XYorugyuM
5tOHzvsaxan09crUktFA6N00gEFAjuc33Th2DsH897JjND7Q0At+GKjmewvZXJX8Lhtfvcxc2Wyh
+Wgn9hHR2jl7dlG3ogFTifByCs+todTegnqPTZySZrjyaaS8JjaIRNwEk3yzI+QwbeoAUBH8jsxr
mtGjwwTnWmzzywqrojSTXdMuMbjqrt1Ngs1Ucg6DZLt3VbNmnDTpXC98MXnwxuMW31TUkdlE+fd9
FHH5w6rXBSctk98de75S0+JvPUFPYdy/4XgoLYjZu7A7Kbd4jbHifUHqWjyCxc9XNSrWHrxVwCCk
QgFvdrV+aWiHe0c1VJ6cSTfcbHbhuQak9M743gp5Eu/B5M/MI333LpnvWuQjfC9IBdHUB0PZBy5e
eHVCSaYKAYCKOa+lepLJ5a1+MUdYnw2C8QWIma4tcl22v+ivTAqvcTbTore09a8u7iT1JDi2Ch3u
e0TjhbdeiWaiPyCDBoOhWbq/WU2qLfwVfWBnymNIHCOxVEWCpDTHftT6WwVmKPYynbhUVm5CrwF8
gcNzSARQ7ZFam6Wqlu+PY8qi7M2mT96uaF7PRWepHBGMtfTUm6W8+CPZXlD+jLaS5BIOFRgjrDvZ
ppf61Jpg81luaASZscm4stSdheFPWfXT2ZJrwV8cYHiygAuNyeVDzLZYJ9SQFc6Y2LZyZCkTr76U
Tslm3xhPFkFx5FNFvBUA0QkRmrVnJ8/0SQeT9i1HYzI3J/+afLLrOyUNQy/g/JCBV5oQF5CBQ2Ie
9J0Ju8DACtyXaLZM0AIB9e+XnknFAnLTmU7w548upSINLPpkmoEBe0zgsY7pzo+itMxhuXoAwUbW
WJWcbmLKUG9HkeknZ6rCouvE7gXYwdjZEKbBVg9O++odYT1rLC9PtSB91AXB3Eqzgcyeay+pRwhS
Nx85JngMUHy8TU7r1ntoh21FIlxN3tkrDWArqvzpiEv09nCjD6E2n43LdTqOaqUf+EL5m5GOHZDF
nebDlNUd6KpsSGWYNkE/PFTr/9DB1XkyrUeWx/wBN51RkyFTI+kDTRS6u4ui49fzvcrwy45a+Ib5
LBo7gSLZuJ2NpkHhhUTEZ0O3Nl/pD6eaKyEarBNEGCmdCjH6IHZ4AHIJwpaOqj1RFeIJig12K6qS
LIydbmZGsoSIX9NFSrzK5AEssVAKbD5LmiAfNUq9iBtqaBwiiI34rtF+EhqcQeMIhOAF7ISHX6VS
LL93qea4m44nllagZAbRFATMsAvu0H9NV5w8XG6aY9U/zpcuMfeuwoJ9umDYHSBj1es3AkRjYAC0
HitPMEInTPsMkMxqleeqj9OdWS8IV0hUGYPXPnKNLNfU98W/xhr46Avj7+WFEei7cO6ifP0F5USs
lNQZ7uMAD8M1MtFpsaRRbKC8l9W5B1tc9J4g/3qOhq1ds8JSab5ZTmvFHNmelYa4mHE4QhqMWjyY
GIvV29+6P+T3JN0eEN5nEA4o/GCfSjUEihqS3j7UihtKMbReQ/kvNJiDvLyOyLnMMr/ewJbp747h
jRG7zJJa78A2LBp1/Ii4S3eDSlLDF++AZ02esCt/He530ZPhrIVbFsH010kP9jJJnSYbwo+tHvDg
nH+z06ZCENbMT5wlCXPra9t5JfAD/lz4qtm4i8sbRlQIKAXj5tuAK2A7MV3/cphXez2EAyJ7pee6
DumHI2fJjSwpo4odZQQwGShohFjLnboyQ8MSRTdS92WkLWlj/ydBNK6eMTpLRjLOrbT1Fo2KixZ+
b08gSfgBQ9HGy7a9GonDtEUK/sTLbMVR3fdbAuVn+VwdduXLILODgy4GnCghAhZnCSpX0WpWQFFU
p9kk3fQ3hdrMWeDjVDgnDsqBGm/ThLd5WRbTzj5F47JpE4GRZ86N0vxYxV7p3WNIav6tkGKomz46
0TDxC8WsGfsu5G/PaCnJThD/ekJCOa+cN1OBjQW6B29PVsJmeChTVsnHKcj3G9utcNiKLum29Mkj
me6p9F9CotkZGVkWO5ODm/5d4oj7KxolhG3kN0FYhNZ1pMiW4jNOhHQ8oDaFF9J2OOqtIGXdWwvc
h7oSA2Xhb+Z0jtLCqgiLHnAiZ49jFbY/QhG+FYJ5ypuw/lIc9diR0JF+d1+VN53uKGsx1mabqvHK
eVJZkJFgr7br9nrh+qHeHsmAkJluHvH7LxL7yiJ/m5+ebDhb+omxjDTZgHYQWajUdtbTuS6l4Zwu
60ObMc7iOrw0j8gyJWsBmiOsfMIOUW+af5u3ZiEEFPhjL7FTupa4yroaAU5cF8ZdPRfzfk/FEBfw
BQEJGJJmHJ+K6ykzhLuOdwS+T9KNGDe2GQNrJstJjAnmq+N5vSaf1M+/KMKbfgH5nU5w6/UJ1mdM
PRyiDB6J8OZKJSYTaI4uc5KexLYWA6RQpwhP2G3G+r9UaqDpvmYmscueOzeWUE5FxwsdXSPgKiZa
pL7Yng8+Q9DBBw+UUJ8NhRE8YAoMn2VMq5wuQ6IFyq8ilUmWHYbqEYEtSQY1YG58j1xpT3SBAyg7
OqHqTAhYu3eqmUKRMH+iNAD31Tnd2Y0ZmGASRvzbIzr9/KPjXPyNA0YVTq1No1O5NJOjgn6HCbzE
Lt5M/2hPKxr2Tu7/3UjNsquPtaxU1XZriYGQXzRPezdthMMNq4Wls8EbVq/82/ohi2Yrs83pxQBs
mThsYrsLMUFowp/u9bUoO4KWXyfno+9JxyFavcIYOvrlTOn+atJq2ZJ90nMc5j1motyd1Ypl8/Az
/WGUOyU4F/wJVqU+Z7FUrJhhr1vjFiWN6eMge/MnMdrdtdg9iId0WKlFID20XeQxRnZGpnk2Iqk2
oIfB4XSvYOe6V6/mxmv1KzZUs14wkwD1Yrny+J6izIwXpXTu0VrhNuPGi69BglV7ORPI8dVWLIIc
TU6xNraNNRb1Z6aWP+ZLGIJyIpggiKN7HASOl6qpmuPJMAboLgQAwaoVdCZHcinP7NDYj9F8Qe9V
Mxfy6Izw21eE7SaTspvp+7j9586N9gn1RB8SaFVueYIpkLB18HUB10Lg8LxKZcWOxPDmUWKAg05M
YLAQYTDwU7VYX8rOD/SSMZz2dtb1khqqIB9hcLtPqRWnsIol2wOPpEajPKg2g93EhwFYmpR3V1XH
E6q8XKI8wCPD5pfkylqc/Qu/IhDtRVJj491MO69VHor7bnooHgVLn7rGlH8RovunJVPfJ7Fpocgm
dxDiZR4sPwGVKJ0vhOS0WSfsW7p/OAEOY1M5y389ot+y7YJH9P/AwdBE/InCLfwe9F0M8Kvxcaoe
Q/ydA4UwWO4PcLMd96Pas18CMSWEMwzRIGXXJyAaou1U+U9SXPrwXi2XPrH1AU159HJtf8+XwneH
qzhub3WuEUZyFrxcBlRf7lpqD3ZjWO8tHSCo5BiKCZhx4ybiM70hg8lybGSBzycUPqrFUc/BMdtA
fvoAvy0fXtEFtJiX6F+lSaCYi6BLbxwkbRNmiDPdKJLW2rBeNJciWOY+XiMQJXBYy7W92dF5XLX5
qRgbdjJcdIfgauiiHVDi1a1ggu8JFz3jTJ2FtNCCOx4nBFbXK7TDiGmNHGdCm1OCE+MAhDwUrskG
4PXNo2qOG3iTOK2lnvlO4hc/rJcVv96+CddaddPmtIEp+urzvjWdSnNjKJVwiKV4WnZpJX8GF45k
m4YjUrPy6FXQqxTfpM3LlSOLhHNuVXyDiToEiOCwC7VMeSwWUF7568+Qy1tUoJCTD1iAqKhBy0Za
vqIPk4bkoLIJK241VrH/YQb26eGLcLu8fFAv26OXxc/76ICxHtZ9XHwEaDNV+LcTF87Z4AoQQFcy
85YdVjL4cIXv9YfuB+e5JWdGYBw0j6j6KzBwKet7PhZvMMlmUVvnFhx8D1I6yjkzjCcQ03s87J2h
8TUH48k/ylL0vtKZ5+d1j//fCKnCrC2tWX/mmBYNItQF/EMxVv+NsWpLRQ00RDU6Y34/H38b/Wph
lgkakqfMYihjNn7CruT1C7wADnVavZNLB5Di8MosfZJN5wmFKz7akSpn275veswBXFPUNcJ5E8bK
xtZde8IhYn4nNB9HFh54p4SFbQkkw/jWNTuzbOb8emLeTdNoPf1phsTwmu+ZbRXy6+zLoWXhOHag
ocbSVXemxWXax/7ym7uUzUpMFhQ9uQNS/zJWOD060ZqgIptl/rIkbu/uQORiZ8aoeYk+EUhyCWXm
yLr0cOKVpDqlhuzuqQx5tHjpcr+v7SveOaqXic/SiDY2KsmsXzvQAXuRRG/4ogJ8kpHAxSAhD2z0
e6s+/je5RilipaCGon3VuPfcnbgcUBint6SQ4vRgalUrg5uQeDaaffjEvNRHt2C+22zZjoFd2gmz
RsEoVa8C2wOnQovmKbDp95ttNNJvDJUR1+JdcGE+uauphkEi4bPTFdozaTJ+zZd7UKSGN4BN6Nd1
e/2MGaXuPZeivFHjU4g+C8m2DYou1o++5hOtdl/QFnjNUSBwz7d5fTXOArazjALcshefmOaR0IOo
SofLAjqBdxzoaW2A8HNuZJ9YQOfrVC6QxNr9RAuy+dHnmKUh+7ijSawg46tQ+rYqhWO0kouaP/y/
UjIHcsFcfy9lwlAyYphtxnkPIEmcYYs4WXKJ/mUOMCfJDb15YN4lhse7uCqUMyiGAl7+ufQtxa62
OvlL6Tr0T+tULWp5BWrGSUfHGCWA4X0pcXH+9UgMYtCJkEeCjZs+2ooE+TGDSNrSgeyHZ+CZWdSE
uigrWMhrv52zgNZPdpqZT4O7cQ3nx9ZhxNpRyr5vRaskMXtqbBftFE9899ByN9isgjEwBxj5y4r/
AyEU9b4wlyqjNHcdzgwIMAZjS5jFoRiDD3mugVF7ZPjgNQ6WutvphML45jOdITm3NrpUEOAEeOd6
qFKyExL+2M2H2sDfSl6/kNszsHMZ33sB9nhSZscdYf3/uopeUu//mwd4fLKLIcX2v2uOvc64B9Kt
q0YUBtshFVyIxTs73y3wIl2SUHrlfyywdOBaWxWRzFa1WpihdnTLmRVNw3+ZukNPsuM04341UkdL
E/eU0iER6m0ESMsKvvp2SmYS6bkAXumVsskw2Gj7qaoXBLngN07np6B79E9sRu8ix0bQWV8neAyo
CaaMSYcx0q7SZNxK/J6lg9u4Pc7y5q0FVTP0Cd2+K44cHCP8p7kY1MyUcS9Lj0rGDqwom89r6pnW
lB0ibOWgKajAyqCV5bm8TaS3UnFgFxF7soiIpihWGEw5LKRaV+gkOAjn4nUwmOAAJ5CbQ+/VLH09
Ti3X4KkQmcykM48sE3msgNrrCUVsUe+lH4NeEkC9j/RwYRgWzX9iWqRGGSFviOpSTCIliKaPCfFj
M9cenBv5p3kdMN4SaeDFQxQ3/OujsxL00Yg5K6y23ur54ZxmaOxBO/tjjD7P1nrnweWQZmJLEp9q
sFElzhR00DbD1v85N5MfSCLd5lkE3QHgPy4NO/mumFpalJiPXo4coMskLzYqRje5YFXV6f+0bLKa
2ST4jdapz4JVt3aFfzYdOvavsR9y2ObrdCJsz39PKoX/dhZrquVY+Lp5VKD16+dulJffqTeCSQoh
flOYT25/G/q2JrG5VOr5toPRB744s4K+hRxuplvGAlN7/tkYPRMQ6w24VllVZ2zTyyaf2s/iJTCW
WBLE4vGU2qzWDO8D9Nktg87z7o8torSw4oJgg8aSnRq/tXFsEqngffdkTQGMpM8UyqHw4GajBV5M
/xQZE66I5vZ790CYyX5IMYVa6SKx8WgRYE3B/sfqq410Tjsk5VVcxB51SKQaC8iNyjXuRVH9KkiH
iQld3piRkcDY0TEOiAhW/qX5OPfFB0EirWynhThjrwYgiY2+3P9sz+zY159z9YklBKUr/GrH7NVW
lCswzU/NPPYwlSFXoXdqEimYzREFFqvTxYWTeeLiommq96fAkBGGCSYGDDsMnSOBKYSVVWP8KnlU
XFYEnLhPQnWD7UqY4I4Yh3KtxwCSPGAuFpBk5Hx4YhTZ2rD2ET+CBIrSImKu8gUElGAbvusTadLR
iKRkHwnSfp5GpLB0FFCaibYMkDm4tV+rwdz9jNzS4c2KswyKf8g10YKMyljFf2VGIhKx34m0lpjy
4g5wabYgxzOX1u+e7XEFP0Q/qHTc/9Mb/z+1drxRY8qfrUjwGmYI+IuqitgXxpmDVj2EmwEJkb8c
Ij3y5V0s6FUk85GnTAEhYJRwb4RQ//Qnmg3EjamDdjCYPnmT+W0E5uclutlPXEVnsLfhJ149AHW1
/yhwJs4DaPqX3kR1XydSSEIHvkGoZl/QACxfiwGcu21WjslFoELYVtR5OruzTMV8m3pjHXVZc83X
sDwROOQ+BhW31QFVBYgp3M1Y9UXJpUbVlU7jzcUd7cQIgfiGQJwUmvTmDHdkR8lldS9Jwc4dwWHf
ALdZ8rKd7A+WUyoKy9CKTYwsNVC7XZkHGl0BGeUJIChd07DMiCly22bDVrKJqkYjNAq4yQXExUB3
D/JY5e0ebJaHlkmeTcaDfvpjWe2PiU3UvzdwCTkD1DwPj0kiBB0LDiuk/k//e7h6TcaaYurY1Vw5
wEKnIMH8EzwJ3jR6xv9IbXwV6E36zI7xpnnFj1vvn+IGS6tTtRSZrw4g8XF/0ragNr3lVxpFcs5x
vZVRV4DvMrB2Oiazr3yCqoX0ULaX5Ip0XJV4K5kV3MlgL80D6QpoG/6sTR9zY8YdxsOObETymlup
1sQif1NO+Uksh55weyzT1jThYijxh9LTboxFhGM5CAgwvQzfnh9AA6aR8eoL2CeEaz/sDXxdoIfG
wqk6sjlNJC4KyVW1WAoI+Ws+yBNSZL96azWDmJzOVcFdLofXAolJiYr0547oB9+LbPW24d/5rWh8
snnhr2o71QwJR4j62L+Y9kWALtqfgb+j1C26YwUkBFqezn7MJyLEp5/fByhkMSyrjmsEB3bxm+CA
E8hBzUjzjXlY4vWUf5p42rgukEn/Oo/TuWAWYPUeTX1qNurghGPu1cvexd98LVdzjkShab8btbce
qc1Vp4134sf1RbJS3erP4d0iQQkya93J645qLrZfVb8OzcalKMSnLVpP3Zwm07GhSEB0Bjr2E18V
9ljpcvk1jkoL7plSDQ9TXQTQIed0YieKt/fZsuzy8cq/Dh9eUU6RO+f/Xweij4rb6WpToH0wYnJS
IzOH83SQxXvbZEllNmMlaNR7DCHav56xMC8DH5B8N0UlwOymXxFRdPcT8De1j8ma0D1xNTfQcaNv
rcEUvqju2J2WxlGtTMepMS+VyZwRiIdIYCJliyZReh8Awjx02AfuNty959g1bucmXnWIqTAeKcII
ZH2Lha1ng2yz2Q4fYhkcbb7UJb3K910DRo8i1c6z9Xn3EQEmm2qx+tmyOqQUkkgXgKX+sv9LZXah
DcKIxRhcPuqv9zi65H34QdOk8IvS8BrBuRvf7v4LjTdIkTIbE0qpOpEDv3tOApDwjYiwNEYfvKZ/
GKjGzj7WhUeBOX+kZ8+ypJsb/QQfk/SoyPqqeZL1ihkGuInKiASTnKWaGCYvE6XizCNWHBzDD63W
Rq1tBGj5AkC3573XUHA+ppf+plXbbAR0yj12xisgBpktQ/KQX6EtmuX97Xas36/7X9gwBLGJ8cL2
shZmtyRGPKYKyOPigbrrk9DemK6nQr4JeP8ZuSr5wI0WKmpY8FDwFjn2kDDNJXpeVHtrekNrqCrd
elqyCvwmsvfwim3CtvpswMDjAAE35IkQR9qNd6jkgGhbu4Ki4S1HeiwLGGP2TcREAnE/QrVjATQR
ArfebIICANFeqOdH5a5JbZa3Y/sAMtrbNefv0aO7agvVWU6dmFoMwlu7XTKE6i52H80rZluJciIQ
PqxyMybbkZ4MEY2vWOzOSrKl/EU2gMk/q6oBdEQG3YCHM99E1/NgynU5Sh/2uPTQTszh9MuKh5MV
Dk20dPIBBpH9KPMP1fMwtLXNOux8qfbvH0CPeoh7IKM6e6d7ZV9dRiiOL2GY+QQ0mw4x6Myqi2xK
bKYa40dhtiH54/7ebJKKPHflPgSQqXu0cw+yoi7ZS1Mzh4mjJGbD2e+9cXnJNM+ATA4xmOwVe9pn
esRGWxoLF+SBqXIleiFVks8n1BNes57GH/47nxglri3o2URHiNzi3Kd0o12YSrhzRQkEwLBIRBrS
rUuGHICgakElHoiNNZyBMm7qdcvXmLO5/w71MFYunBTXX76DJ8w1OBat4XBLI5u1Sdgkf9U1TpOm
BzhOy1E3MCOitG0m4txxIo7CGvZwmKuDrZCvCdb4m5/iysX1qkkuzPFtlx8Daw2vt9H0GrsCK//O
UMZRHy32zx0gdojwMKWEoJULJwnow2tmM7xpnIdiFF+CUfwmZnDHmUw15t+MlxCKj8XM+QxKTurn
QE6Aj391PItIHYMPAPBox+j8hDb14zrLHgqnSuII+QvxOed9XoS5l8S/cLVnwe9PNmnB5LTPvXU4
KFbqEIJ9OD5ROVd+ckrhaYmSB074bXu9uBC9eDPGniQ+d9EAgWjDDLtmnycCNSzZ8c1uBCU2/82X
nDQmp5eE+0hAIBJ7z3hgBIgo3OZYrxqKDaa8DVvMpkKrp46x1jdHsqLBAFomURTyxpeplWX8W7cQ
TMxGlSYHiFtkSBseeX9WebqFyhlBhwyNTzCKJfzQ4Bd71/tRo2pRwtPIjqsnX7uwkBukQlOdunF6
pAgArVqufZPOgmtjw6iMEIHggkyTCWbZ7Y2Jal7vKzRcDU81yMkAWEox9spfAdZEE4REraonCJxB
qzptCE28Bipqq8YQr+ehYzQuFI253RXPKZHKVhkfHmkPXX8Mvu/zHgGFqM0yUcl9PaCF10s/uEOT
aBwnF52gFSixHLEc/LI6NneoH2/TjM4BI52efnTd9rcmdTpUDwZhNDLoOynd+vxrVbyCM9upuv93
NxnfGV+0JgTwlCHMoO62dK1zxvixRESOxgTOcT7pE8kQf4BG1b7dYthQtAWIwTyVUrEPnRPNz/fq
umRH6DY1nrAukbq6PfzbD1gklfK3HA9NZUH48Puf/VJmkIi5zOcBgCZUNNi6fZcQQSBM72XrghTC
v5LHRYJsvXSAJG+BN8KIbVJmnk5z9iN99Ijj8eOJRHIa5EiuL8Cm8I2ok4McBbn/uiWu9UnqQ1kB
rDOECwfZol/g83A3z9C6n8UpGEmrkXP74leRuU4eHDsBW1eK41jb7N61rWBepgGmRnp8vQ7jRpuM
MujsDlis7t+Zgfcvh2v24zR9kkgv0vZeTPmLgDuGXqy9/Od5/cuKNyDsk4exMjpbOx9knjY/yrZs
/fl3t93zjmwky09T0ocLQuW7XF+M59/3JEkg5s/jPz3RlFEohm0SfCRkrg8U+r5im+63kx2H2zvD
Bio0W0+UAeYQ0yw5bk6P36dXCxFWDGySzSqQvxXBayqAhLOTrgu2K/5SXNvSjSJx3pYA/KOtn7Ld
WrnGwQViJQwi1XJWCkCMaQuCjhFhPvri6HSA1XAArigOXeke9jBex9MyJMLy9ezin1c4/LHpzziz
CG+oBItp3MFiUM78+qYJbq33qHDssJ1emmCnuRuWPuHMopFkCZhdDkZ7RUVjTD5B4p8NdTCNMxX7
d7JN/EYNqoXkDn3ZneyekAkVSr9Ch/PllaR79/+fNl8JYKWKuK7uTZdYbaRHlQziXcqh7rEDzcSF
w3XlobuoeF0gXiw6y8Z+3rQbUW7g5SlnYsJlqNu8AJXt7fIxblYoCDajPgNu1sNq8z3Zk4mI4a/2
+bznOZJslMbErwEq57IHq0vctPoIaq/ZAOnN8sKjNwD5SzzOshLJkXlQlbMbk4Zh1RXnVdWKOZCF
ZmGGn8sdDbDw/eEYsZ9XNd1rKl0RZubt82D/0r63F9EkRkKDnX7R/f181xCqpeT7bBJ7pOUxsoCW
E6sWD/Gk/ay+kTqBKU/uaAy4BP0vBcmhUrTaGEQRWAyPBLSIrKayENGZfpx7H78zAQ3bDEZxX/3U
EyO5WmZcslFV1zMNbqa0yoRG2HEk6CZTm0u1SV0DckLnSY7gTUlaMuAsMuH6UpYi3bD4DqoltLcM
2UM4T014OCfHWuVwZ5Nlp3duQMQqpvh2fS1w/YToxb0nDA4lluOglYHRSlv1siOIp0QNK+NTKXjW
XnBwqf21h/hG+VuzT+N3DimuExmuBVROqQNLcPlHMLKy6qD1qdx08bnLi7Zge97rltj29M3fJs/b
oJ5u2k/Uvkl1SUKganCe6pr38DSIfIrn4QAMdhbx3eSjq+F2rbBAYMwvdSp2nRm03C6UwcSRZaVQ
EOzq+hgi7fr3f5KsRL5hvY8bD3/9/34UmZdrVlp4w6AjV0EDEgvayDxoCVHMkWjZk9wkDIx/7rYU
zKny6bOTgHTg5Utu4Sk77xKgmTX6qWZxKop7dln6fCdKUn/agC0imJdr546LwpKBEGL18lWV0MLf
3Nb+rS+5dSJvvvDm6mKFBdsM25UlGHC9dsNJfVmi/gRTwvt7/+FRvAByxUK14pewk4DOv/g6NGo5
KbYtbeOwOFtsCI7AHkBcr8i4yWClhuVmRzenOy4AnNhfqxj5k9OGsHIl+NPi9Wi91BgymGhaMC3N
tlIBbpX+BKnZ2xBE0mP2cBCoS3BAdKLYEvWGAyanzVbvLIFVa1oKrXZqQZYwt08HPtewxHmG4FYs
1aTKOtHU3WBSwftUXLz2gvoCuWVk3+tqYOO/7jagm6LyULMl7nAZw2Q72kPO3hEH/Bun/OS9SdrR
8IQx3WH1Nq3fyuigdUY0Niv8wUewd7L08xSzjG47WNIWZEbZficC2bOfnv8XMoFmgi29HbN4B4zM
jduABh7DLy7+7XB8S8inJm8uL7Oe/8r/nxBz7LZ8CIs0VmDR6pELTenDdiN/ojUr1spaa72pvcVp
tZEoHjcxCToyn8dSWeg6OwCyEaUXHa+ErDXt33c/qmrSPGW0ZhavpMRt0qfSOBWTlcV+6iJqFgHv
A9AAybfBXNgV1ulLFC+1mlE5l/W7Gk1I26AR9L6kbCkkFxbxFhYNEKAeZsh4VeszLM6IYzhoBTRg
sIuCC+Bf3CVKjWqDbLx+hRMVVlXnbWXq2lXPjzF1pPd/JFVw5arVwbqpmBucIKIB0EwKm2zhS9nS
ZQxRPL/rcvqvFb6qUZ2nVGdVClvzhGT/tqrZpkTS1ZXngYJGLE/aYL8UAF84jswgrlCcFJ1HLlGS
fcBhvxflOe0KQ4+jl2sun0xwIvaHx05bj37j8s7R0mKOw918FOVzwrO/xR/KkPnzu6+1gIER9Py2
WPScMCX97VYYNkpDA6aZ3w46qosCuUVeisCJMdcHuCKAc2JTl0ndFW486RgRLhhdUvIMj+ZuzC7V
LYxfAQp9jX78eWvUDmNKkJzxmEn7ZUmwNsSoD7ip0xM1HI2zYbbB4scXU5lFK7bGT4+Rt77iEWJ4
rlVvsH60dmm19+9XnCa4QEinstjEb+Mn5p5e29KXGyQPOulyfvfsjf9C+WwgbNRS229x4IbnRh6x
QQAuPoowLNUlJTPDCoXX007k7NbCGxEiLxeO1oy+KfAjT2AlX+qhk56ZL61sFtWePHIG3arIBn3P
Q/jwK6nNS61QRxSE1N3IWa2GJGSlPH5EehfF1cxRNIFWc/cpx1MEhVWbr5oMfyNm2jsAOUAnnHyY
KJVS9mpBcUxj89xShmZJnzCtEaaoqoSVp1BtzuC3Ub4mYmRvcNrlvCcwZwnOT+8Pgi39BvqJnUn0
0aPhpnZaGEXJwIYWWLLnN/Bq5Qg1OiUDbtwNn4EgqMyVi0wYjQkOHpr/jHekbJCaVBdC2KZVTfLw
jM0wTx70awIoPoSRi9rD8FEM9bn9ZRPktVrneIvVqOw/z7o9ZpFM3C3qjUnTx9babgloR7bouu4K
X5N0xTibyf0lIRB1Wp28seevMvvBiypYuEpblY+qZKUse9MH6fXphs5sCY+lzNqMzySipE6xQjws
ThXQ2Xeqh2czl5oyOrHVq2B9d4gI2D4zN2bC1bxbr2NnYZyejk8jZVp8LmEPvOOWYgBNkRnpm3RO
/c9KAlqJ0889vGmHSPqCBcHc5fpdnpUiBPkXut4H2zpImeC3Y3P3khicw1PQhqld/Gq16J8frggV
m3p692Mw9gjgx/GIuCCICgzzGpUjLb1tlPy+Mzrhy2vNSo5gDlC2Ewj3cV0c/n405X4R3aqgy8Aw
bAE+lamWFOBeXuyeME9oLvSz6H0uJOYMQcmBrPRLrBXx81xxtBZsUE5dfA2wK9s0ZhmBRpgkApBn
iNDUzq79jYd9+UtwPF6S6XpW8UjJYtVRFxAx4Z4bdYOhDaVovYN8Uo1dPQeSMf5dilhk4p/5hF6E
eXaLbiCat29SWqN5XN0HHW04KLDdMfWSjkZa+gn7zGZE3ZPV0/C2o4uGOCqDJYJiSGrUme0obtyP
owLIbQcVuVWt2JrRE+x4JSsXxlTafGx7yKo/3NOooqhLjt8VjZYkx76gj8eohEdLjW/lMdFHrCh2
bSBYhcX8Zhq9ppUOx+v2vFRkp4EkW/V+7l0pqVkezJE7wVUKuseL6UYr66G/Ip5Eatquiu0bLfJB
KWZn4j6R1VV42pIY1kwuG81v5MDLZVT7JKByTTxeDPUlMsKVmd/jw2DDvju4hlAafgV5pUuuULaM
SmgdioTjGKEEoqBvtHgq9eE4IHkCA1Az7/Shn8uyTVYfYbzpKHMb/GaGUIuy+dNEWekCslF4dCiv
aLEN41ztZxn69YS+9Cpe1fLcG/1w+sDn9HjuwsikWTw3xb076WG3KdUmpnlJGjG/EVViD2ustdgi
RdEaffHfF2aCNlrmBJYdEwvfZWgitX9gCg2U0CS7Fx9S7bM6wSe09ZrILO5u8ZfYJUDV4awuM/Il
Ghgqarhvam48wx3dlVLk5XMlDK92Q+4TcWgj+Sk+teOp5NMG6wx5uJnKba/3O+5r1uqYtPe9WhtJ
EJ2hfIqnwJLt08LDYYo9XIVZmrep9kBRY/Q7GslnlKxX8rpBL6TWul1oelb8yDr4gyhGdZM2KkMU
W54qsjFsB6YhrFTsfzD/AkVK9Ypd2hbNNzKlZgZBFbz0g8Qt8ZQjrPKBDIUn59G6pwchQ87MXWxa
itn9BpdZyGyBYf/1Wih6YicmFJAT5sPinbNk/+YvE70HU0UbQ4A2oce9Hu1enVk3/mWUcoKkZrUm
Iq+Olu4UNz/CymZWraNStxcepgJm8GvKHPaND5/skJ7XbuRvk3wfJBlUO9XPigYVWtBb48t5fR0o
A+nVaSImk0SLw/1LByiDLLFV1NY2A5QHM/kAbsUiRLDgYaGN50FopTvhtvwVOGyQMjRs4n2OPhXb
4uTX58O4gy7WhWPO/mJXoBG/lV9bnLuKlLdfRG337yfAAbnxRKjorL+Hd2jIayzaD1xtZEaM4TaN
6h8koYpRhesXu1LfhGqckSqAQadoBjUBTU806eqiUVsi+oQRf0T6v1EsYR613/kxyeCf474f+hBZ
38CAU39vBDG9H/IPKqp2isGDdWQ/UzjVzhQiGVDxdRHjB6KB7mIJ8dwS9R7P/tMtwiW/vRZ/TXhJ
gg9hXPNloSFWTgtLK76aV57oOulobLhZodvaSZ0oX+lZPkKw707xTyYTvGWnas5aJjF4SCY9pE5l
7tU0j1D3R2LPhGsdNtlKgYJrJQdclC8yDA0wPsyK3/ymXTz4bz2exhjEGxa29KFqTvuUsR7uOQCK
qDveBPi9UyAuq33TMZoZYp7NIvhkJroGPD58/TqGwxIVQ24Bkg3XoBnkKzM8AqRBnEXgUqt329xV
wKnGe90Icbfh8XWy0ZfZlP7DmjX8XrHSz7VrUs6wM4AFkR4zerZf2hBMw0OZ0mxLLKjCZdv2EVNY
qQ5oPMjE2JA351ELFf04vlSesKtu7cedra5nHp0XvfgtwAkxtasjqeQcxdCTSW/ScN1kcYoTvUbl
bhri/RzOBtohGO3lPNr+FPVSf9jij/o0DpdRrSRxAOOeXVcjEu7CuMzMQ3EYqSy8LcoLL1MZe7RZ
BMb2Wps6ZGx1DbjDXKpsrJ8oljPAn8qFnNhs3qQUC1mc79kw9AtHSjpSAckrfbs4Ympot1lE/kMP
olO/xAJT84THsmAZenZPLnAazPAIYverVmrgm9gjk5cukQ+7YHHuZ+I5TyUQt5VSmOZBdM9wrGib
Wp2ZJ7m8l7QSU4KqiKgMlXFlzvUsJf+wLHsWMCQzzvOH+a3CwIKQl8xhn/+Oo3Cq59yTnrEME+Io
/7PHtUIWMYD8txWrG2SGccmb3bkHnsZgb7I3ezYGHESfH6fJVb9d9JtXc89R2WU0nUziv9GfE1j3
zMDM4gc17bI5OIQyiuuqHqs2MHwx5PieCd6Gy7AG3MJYRlHLJMwu4hMJUdKK9MtwzyYTiBc0D/f9
dj5TDL9lRVB1+HTxBcj/0y5yVOnw6iNcg30Wgem1XlOfcd5mrYwxnycOH+oOmG5vyOgQrd5fC5t9
o0Oe4eqzrYnsgRaggeLHzW5WibiC9zH5E8iPA8aSf6lG5A1Scez7LKnTy+n6A9lQnD8d2U31DbPy
caa8txt2SmAacp3gG8pa10FJwhRdwKBcRYIG3PgcQyIBjjgAPzMDJNe5uaAHZZVFqnDE/GYBbtTW
Lvz/xd1R2nQrwlBmOP/uDdh1f2kWMKMGpJXKAc0J1ItapilsoXb3epG7rYQdakBnJFOS93w39BqU
ZCGa8xtGPF7MXP+j4k1/WdtTyz8C/tB47WCnFF2YHYnZARmpZf2C5wiMLy+MYMFhqlVYdqmQoSg9
6uaMkXVYU+PPlVOPkn2YosEhuoiG+4spN8hKNwV7Qt4hOQF18h+DazqwMw5JoQEvTIF2zlsD5e5v
++dqB4FdxbEDgCiEa9mhDQTMTpCvoMyL238A8CybOhaBYT0GUlHaXiWUhTHXOXGdn0z5ibG1OsMu
6J+9FqHuGXZm9bcvHD30zpsTJqB3CQyUc4ZE8zvJmDK3qv13opvyyrgkEUd5WhWjtAVrBOtr1BaV
nnqFdTV5NzIAtXC6CkyRshL18RgDnoiYw4DCOOrOFHBITpZL2Cy8zoa3bFj197riLarJsy5mcpuF
0tpf257QOJcjVT1czpw6HIMHzHbwoJb2cMy4tDcsBZ7ifc9qNzQ59eczhfUmSqVwnaqA6QcU7/yD
yPtzlInIXUv0TRWX8MLXY/uz2hzTe1QDRIp4uD2RjhWQ0bkA1kS9fSAm3wrxAB63DVQvwKrYeYsk
M+5V9jCtFfkDw1hngKdBSpoFo0PYQbo7tm3e5iaWk8hIFTD598B6zcvkeImBWovKk+95Zium8mUl
RFG/0h4MFdqrB1+nan4bo+yylIjc4nmc27sdy7Me1VtXrlfDyjgZ9z0aoQ5tfepR+wgxvXGJzJK4
1epy9gsGa1d1l/rU/6qzHYrs9pQjkPJSwbwUFanGL3sp+8Z2zSS9mTsi4ZklmjNmXwkfqCYP2PYO
FQSgLgDFB8G4U6HDVQKqxM4BQocMUQdDKhVUGOd8QU387KXqCtjkSDbKP+aHfM0S1qusbuOjxuf1
YzZQ8UhSZ4wpldbF8zNrh5xi7bAq3esFW3vapaksPkd8g0wF2jEOSOkt/iGj6OeMHt0vvUpgC54q
QbGL6FZqx+XgFo87rzGuDYjc2BtW23v/B4+kfwYxCeVDFnJboJjgLDq+EBaccaup29gKvabmYrj+
CIvrxwBx9reWwH8CX5qGyIbQLyaNsmA2aIpW4Drz6GGu56yeUYUgDCvET8rosOKkNcQDO16tCfcB
7GCZl0XStjzgvUGRI+pX1363FxzIDs/KttqwkT/Eny13MMgALZu51nGwNvzoGvZDYpQm0kKmabXE
9X4WhHtIiJv2jA7zcR3FTWvlF4j6ZD8hMclOOfPP8uvL3PHYRF4DenFkab01C0egfBhnDwJXilyk
6ud7OneW30yVJ+FktbDlKdZVQy13Q5tZi5XT6qdzMrPI9AmPMJc9tfgQOtU7qAmlczrX+7JGLA+m
3Duqgi989wNihaoCIjLUfe++3IX8izOIR1kutQhozxpmNn/WeKBhnisupw8Uv2pNfR6e3lVILSRu
U02v0xdqtWXm8TqW2OtWa7s4ywDh/b6UjF0ZiwZZvrBHM2PKg7+9BrfHgMXZZPDPVxybUHYV3IB4
2b7fPApfMgZ1jkBElpQFsq83IrSWTIobwqM3kNarAuGH11ldEGR6maMgqY0z5vu9gy2RPAWx3P0B
EJyxg5LFHy28PBIWey/dCi5hznGZ40wR5e99jU/7O4fDgqVTIIpj2AzOELnG62QbsqYBvLtjq3tK
yAfqStrrCiSjFYgQ2oJebgJJ9wkfhhh3V/GZXi58b/SYHWls8F4J56EIxMlqHuRGNT+PhEB42iU5
WG5C0O3fe+Tj8aMxJVKNpkIoNNqG9L3o9DWV4OTzWBNV5zuBGyFsOHQko9DtfU+1jLG34D1ZExKo
5ZuZx+i9Or6ZGgYeVoD9PzqARCfoog3xWzpIqQ03DZ62LUeKriyIaJyrSWxAwBb2K1HDLpvPYrco
21AbeqGAMA5yNbIJ9N5NDVtVLJwi+SIUbA1qnbEUNLVtyoPDBXkP8VSd5bQMQhbT1oAU4koZ+ZJl
qeFJDG5Uvw4ENDkwXjYPLz9imbvob1KySWbFA9LT8qDLTkf16nJzePnAxLUXnnSmvCRylXx7qH7r
tS7uLOxLJcfI3L0rbImmk+BqcMV97hfpz7qGZROiNi5UbSwnhVuEHFCeDemAAg30YcjNHR06b5sf
YlhHUjmIdY35eHGc0z7KXoONbFzMv2QcMRmSkS+YI9z/DRpjtlLUYshPOpLDXXKxF/CHxKnlUuac
UfozO0S2SbHFhkwNQYwG/9u2i4ln70iAZ26nMpou+3HOPgpFQPInWgc+csTaW/FwPt7EGIlugbCl
vLQNYFtLmrzmj9JHd7V0l/S8Wh91r93EzT9tMpk940dHX1VJphGM3U+hzpD5aQyqxewhFbKM0XmR
tlCc6NJUb2vPwjnbl+bx/ZD5VO3PcMG20fNhozEr+ASarpv5FlkI/nSlLZSF566D0xPxIDDQQXoD
LNCfHaveBrxbxYWyYgHX7rgIShjBLGa5ONGN96x2nOga238xiltgZ5TppoLSQiMGxwEMbAZHcoEK
ztGvRIYYo7I8tNqcTgN5cSAD5l5UyRSfDkQN1TBZFqAj2wptqit4xDhhknQ4a/yBGRo24XRy1+sv
nZ1/GFM1kaUnXpHmfoAtEUKxqxpTsHRgPDxkSqXjnueM5aAJMaICNR741EcC3DxPXsOHL2c2Ht1W
2UNONINxizABlRpWLyWMWqTG1Cl7t5x1f0gp0IdWCZFUINJwA5r5LVVPC7yk/gp5Fn4boT3lA1/2
0dH58UhoHrvHs47RvZPxQ6f6SXQJLXXZ0NPCvGiSlGDv0D13IAP2KWetknwFDfAwnb+IJCxVeXvK
9MNTmr+/VJuzJZTkBvXccDqs3xHXJYI17mmAMHhUchMXSX+z6BPEzvNktmuQlAN1FIpQpMt5z88+
bAvJ3sgNlIBtXmVuHT11Sflr+fODXMtUMX3J6dxDj/+PYbqmS8Qpce2Y36Q6FAQ0vRQlms3yBEYu
wCH2zoa0XPrZtknNnlHfjwBl2n8tNU6lFVPj/rt/X3vCBcn0ZBbcIHW4LTegArlyf0H1YeqiAH5e
cAWARdSS9OgGzcILgmCEXlYfBncCAFPxvD+Sj7V6E4PWxrwwsSPmzC3dSENdjM6fD8DqlKtAPaqT
2b0COjJPiPKK4ZG1EzHuFgv1ArhIAj85DXBBEZAdXxKyQgTFoL25yJ1sTGNOdJ4LTWgv3Efi5daP
9Ky7222MlApH1/MO+qDspdZz543R4p2gZUDo/5mg2ZfCHMTGe0WOidrW4CZ1gNMgWFQ4DEa3d2E6
dlnl/vlnbq/snxehHvonFH8XF3I7KQIDOtMif5DKEH6eVEkOToHJfSOkCBMTwkiZp8v8shd+b4fy
q3MXEMlxqoNL0CHQkTYckA5ic9NgmT7zG7JXN4yLg397EfL7Kchs4DgEdC1RD+3MIIqr9rQrWYpc
FBUQK0uYyAV7pA88ZVyCodncpzfUe9FvOdu8JnVe315tMIQwBTkE3VtUY426oT/ZfHC56iAFWhKN
juhX9riILh5fvkfUAfXmkPTCOZJHsTCPfgpI5wS+j5A9X39qD+TZifyb4q5UJQ/NAlmRcTGF3fXu
PX+sQtf8TscxmutdTai1zDtYgBBGvtuGjiqUpIFvPIBVaXZrLDHV++mk7XtBg1StNcVT+QLpVu8Z
58pjFfZX40yzJEo9mozh4mTnSAjlN127ZHo9ss1gDVI5M+hlmVb1unVO+n8nbsDHd5HRkM1FbZpX
N2UC+umzjui37JF0HM93dWWdsYDujDmEI4qQeqCS2Z9iDDdm0ykCpaKY3+8V9slDoWYm/hpqiWhF
bYUlDWSph3Nb75IStIu0mOZ5zDAp2vGEkBFXtC0RnrRImuS/1QOQOT50vUe0c6Y3Vu/9OuXl34GE
BNzSbskEdE/F3oXBd1nnzGTn4pVbNTJujaKcbeHOnd8aVbxlYki2vQeFMIJM0lIUMXDRPnKTnzNS
tuXMopmmOE3JB8VajXPRSxDZQV96S3vQkZnd1JHcY+9IBeSymbsMlwluWVLHScSklhF2UMwCfpyH
ZJUFVt9EWoLPX1QAWW+lD8/NwjjyQ56LB4n3oem9oE9a6v5PccY15+MmCB2FycS9sq7OSFBAt/3l
5cbqfZ586OOzEOaEItnItpi+cn7SUOfIUKs1M2/DupsUUYQPghwVjs6wOeAhbTGQfJFEOev1lL0s
wFcbUZWJGcgXdcf4zWGPy2cJR69SBfuzqWaNnRZbGol8IisIx2h88c8KPnegV8RAGqgTYKH2pQXX
3B9FLheWLhRbI4QVz0ypvnUfUuW4D7n4yjNgs1XBanXVEeigb2fYdmKrjwKqfucJSfWp+AdnRLgi
kupmz6AKmOHm/Bg2Nv9O/tbkfIELpV+Exa0O+j+2lTSci38DjmyzrQS0jDqOpunopuDF+ulclgVL
bXj9wpPq97wfOmArwkfeRSRNVH3Hwfj0UCsaq8SGiuXuQxaTMZF0Po13PHy1RdfzYt0z2ox8GQye
WYFLMOUEDzEsDeIquJsAM8SYA9FwrJ+hFN1dIvGz7RhNU43/Yxz0/76MTmJCnRfyE3glBghXkfFG
YZdtqgecKmYoH7aVBZHooTL0qjYw8RbjF3C/NtnOpHV/8NORhAl30bCmlhiW6/6W4XTIIgSvUhPZ
8SzZ74qWl09/RuHjSySWQpFH/dFv1Eu/remfetmA1SphGECPJAbAK8L0hx2jt7nOQAQJkJYfYet6
Q+XPEK9AWmlPTFOsaTSrJbpmXPzPqzqF2nUstKRRxjESomMsBwGTSCXns79Zyj0h/SrnnbBUw19L
HImwZiExH/Cml7wc+tVZHaYLKsJxqMDLe7YTlwVUKafnKefLt/fPNea+qQhxa1S6Y00PhYbOdL7A
f/487KPPKRJ9cxNJ7DDHltN2kPIzXQw90B+amAjm0LqsYbOvQb3SCNouRcqlxdG/+B1mPT1x2CID
r4lRAx8Kez+yWktjoprLq6Gax7mYlVs4I8fnS3QwszK7sMl6Atar6+qKPR1jhDl5EUSzaghOrIyY
uYcw090Lu7TXSBV87uYXP8GBqK5RuYNrvxMhotwn/SZNXJc9qZvExTXa1IXM+BU8hhXQd0VJsP3L
7WXFfS6cw58sXnlKa+ib7lqDJpBa0V66nqBx6UKFmJLQcpDA11AZO1Az8GnOueHdLddIk8yMK5Jj
F7yRSGUEQvAKQCHmu2t7feq0HoTNGzpdPxc5aS5qwouhKr34NZAE6X1+UBivB0MTCTCkt6ENssh+
N/hxa0be53OHGcSz4jJe6GzcOr/yqIHBz/2dtLqoxcV1CXCg2+IPLAPCtB9P1eGaNhpi6UkliHTO
dEw9oN1+I79dbpKZGo4YZkjEdCiwwoNm1rk0HcyB+uEQRuwDNtIRRlSPK4MIDVNSO1tdr5/g2t/C
qp8fJQHzzbn8qb/A190EzWIvE3yVEbnq2QOBu/Y+tmwwwYFit/j/W8NQb53fW7iSg0m5LBQGj0k4
xrmIfyw3n7aQ+zG8FFYeIhobJ+b0oaHUgUY1GridxfG0hefR4nxSAJzxx9dgIfpfuDBMNB5yhyGY
w6OKghQC9fg/T+BubmtAhEdBV9pdYzeS3YZ11YYbPkGRk25VAAv9l7J8MQN+B7vLMZfFRBmu+kaw
DAj9VsVnAjWua18p4tbfFaBaOiBesh5ABpemZriPc6Pbk1ZRcuLEXokPWZR/AbhMjHfOQsdMTO9v
NK0Cc3mMM9PCIevqop4cVlWudSm2lE++NjiV2Ejx56NRhGV4IWYKLK5aU9XGYhnqbVk4U1q3LpiU
tbe/y+KczzF1ctEJ+WrYG5t96P3YYqDS0dkcO1Df3H5c5pSWKWDZsvjFoYz5XsCind45gDQAURqy
XLTHy1GGZvYVgG8CeFupe8LUZ6FAk4uh8H0Z0WFaPVCZA6HW2BTiZdHjIfyQKaYWC2Xq7GqdmphD
Q+OtQw3GmAxE2oGTxnSm5uA8AuW5Ii2cKiEonl7rfAyWz4khOQMwdFAA7dEgCi3lFTmJ8vWHDSrq
IYYeIsmQgYYdoDDHd1RX6tiCCR7I1u9C7PjvcDei9Y/zZN4hNBWyeFW3p6anxZ/8kgcS3TFeEGN2
Lp5R5Z4R35yqsu5/RuawSCJViT4b5bSYoZzwOHQaroHRTjaJQoKDVJdjCCW0exkGG+HFoCtP2xLO
hoProA7L1Fo1cGhz6ZC6jSeIuihRWYltaZRwqj6yAEWu2aukQOzeRuXZi+cvFmSs3Wv223qQBKg6
rMc9fkHoqnN/BGBo0p8kZIEKyp+M4mu6eV4o30cnW4Lj8LZ41YqE3vLC1lPKcpsqC9XGoNeVFjWl
5TwyYHf748FPrsszc14XKkWKcwtKyp02o8s3Sd8NY0xJtI53MazHZ7hpGaWSwBt4plNpesL4S/CK
6BgLOjmCQPDfaizFCnsTn8vR2/+1S5sy+ncUR6xJWdC7wOoNBOMn5OzBo3oBXY0PRG1QQ91vyDc+
ERXNuzbLYvc0j2+ZUv/ZOwBlUAgvwJWNlI6P/xDsPiVm0EIzsy0R/lsyhe4Pr2m2IVcSOoYcf0j8
HNKxYlv/FrqqUybQofZHOv+oLKRokyEi81riMlQNIptvdV4XDSmSOoSAOWFIAgQ4N0g9O4ugOLcp
xFWY64eFgPhuY23UT7nwrpknMUorPonjLvnvE3TvSj7yli95z/i0nGtzoFfrHThkwz4C9rZBfKC6
yHSfoqzX4V/mTV0VMgb7VPNJ8+ILOpas9NbuminkDcsWay7Qg1jiSjAjOPEh1szKhdF7UaRT6PXL
lgaaxmRC8hXyZo8Tp3s7/LZ0pM56L0p8daMGqA79XkvVvYddph55rlmFeTErZQn4RuASqIobMBxN
HuUkZa5bgF026+SOMiM25GQ47kJgMkgc1dNWRr/FmfS9NLHmdowCb2gxXWSn5sbzuDqqD/A7VlDt
fgC6VzRFWFlFwua+D5AfplRSFDeAr2ZtiS8IGlNwSlrkx/x3YvNLQX2H4J/aNlmEZA5twiTYY4KN
yf4HhD38eoumBwa+q9ZeP7sc68jY9WDE/DRcp/XkJ53Ai8CaLDAR9MY63/5F4P3B2b656AwG/W8s
/rKateWfBtoO5ns4GlxfzwjD8+wYV8YmtZ9xpYhn76krs1f75ApGvSpWdrI9k69i6vo6OBKPKeb/
Cv/WP1mZ8EkLsTHVqQ93nzFAFJjPH6hDFb7LBG285ELysksv+rBaztjfoYLEgSqM+IgEGogMy4Ci
lnbPJNECGxrSArIowwH2C1XLj4GxCAEWHciXObSzxnL4GpLeky1XJBek4PcOquVsNorram6AhsEw
70Pjuz5UEKsm3VyZ/LDruEhINu14PxJz9c7gO3UGcXgocEa8QC0sknoBhRdcqoCyfo2rib9r3Oy7
cVsvVCvIokxmxHWNDZs/VYucGTeQtJrdjU8ENyoiZpNmj4JXjtGM2F4rbHsdOOszm9/5mq5OAiof
B8q8TsxPOswt9idRHnfnLcj9V5F681PwZBQtki7CUnP5kFE/xA9gsHTWQA/paMSaHyo2FfeFwIHB
e0MBA63eofS/TSJ18givwvEcD/6IX5HB7kyR/AHuMEOQZBojVkYOvqTydVYkoDPMcKHTpQVvd92P
Ch8SnHubrdSZAn79UlSEC0KgBtaO8RVWQFs1jH3av/rupt+dfKV2/KRuSpsZmzYv4h//WsNN43qu
QexBE+LOlr3BUIJuP9MFRtjYj2Zi8WzLeqeKeRcPfekep45iZKdFpD9E146D5YomRTsMzKdcxx4b
NzVflnEvqgnCdQ8J2YVBBce8ng+vAhdgGqpoF2hSRFOaCvbBvGTbGiVoZ0lrUejLyTl2Nazws94m
eLzkWpRUhDTyQYe1iSu/BIEHc96g8oZHVmurCj2EW4tVZK/v7bnrv9hhJiRz785vQ6k1pq1I50at
k2Kx7fHll1J6CecABawAEj06WvB0U7Kdd5M2Y8APsBJHuovCtLcE7gUAbrl4tPwpk83zMFBNQQ6Z
A2jA9aLuUCiPP5saC+nY2fCvJfTh5Id3R2WdzNHNAXNhtX20znfpLOgpnILDq8jeICdrkSzBTjg8
txtxfOvznPKv2Mznr5K054AnoW23sZc8x/BiqCLnnTox3/nEH39wo/wfHUznLuPxC3di8HNW/aMY
vHyS46dunHqcVPyPsdzb6sTrvmNh7G7EKP2gXJvUQ50IkAghN1NJna2roesSyO2HSCr9DHmSEkfQ
FUJ6vzETc+RIzeoTB0G3u0rOGxl70CNa7rHz2GCE9MW/wJBE01QJYe5WmgW0gMUYRmzjlqeDEtO4
3Rztj86c3qtIB7YvKPGjA9ubiksPZVRtSDs/qLa4pm2TkF7dOrY2Mo0WxfYue1GSWBx4U1Iq2nbB
Lz/wK8pjju6CvIwMb2fepuSdvnhcd1fEor9rTKEmMhOMwbcs2c8J8BkXuEhPmyDaXxVKm2A1f6by
yQOkD73Xjes86t5jTcG1FlROzR3ttSDmVODtTVdwgAz3FbSYPPZkQo3ItiGyno0XUafIUmgR70TG
HTy8GsA7xtcV6zDhlonFUvYRDnhHxPDPixwNhTJaA82yZ6ImQQIw9Q61otJZa5zQ1Mm4SrQb6ok6
+qC4EMhvTWVeRDP4ytJXGyiIF71n3A28PAl3yOZx5M7XU8dxRMWFZErVlJ6y1yDvqCZzzT7ipwwB
kcxgNkdIIef/V5cUdq51hrAPgxEUhVaU1PKGnU7lDu7RSg06d7ckmNi2qtecHddQ3IF6VnzHkPqX
ftc+7HYbN+5TjNtNzEHWqy43+MclhKSVQ1KeaMyf5+Ith/DAl/3y4ruT9G8uWLjVZZN10lFlEE36
XEiGkgslr7AKZTMRA5ujR6DZ0JEl6pNijdqKUPuL5hu22eaIf7aXlQEmgP1CL1vo0cMvozA4px4u
ETrxgy5cGl6I+MGhtCQADco+i8kxQG49CDL3qC6T/a+HzR2OrVwpOnd8ftqs+Av6QIKkjeiESs8+
eiujGs7IGNNo4VXKe281Db7uYAdILLcGtW83/QgSfxDgqrze9M6K84KyeGXnv+Cg40wGzkEo3XcG
X6MMmkkmwpdgsJ7PsKbsYqlQAkYyWqIB2dCN8m9i04l0k/X3PNFl7qXP22ESm37VKQMLQnaN3wSO
FhqsGL69YO34iZf15zYefhvd0CNNxx04ENqcDWbOxLOofjcphNaEkhrNMLvzfmqtnIcxhaQhYFDV
6N9IWY9rjA43sX6QtHnZeNMl2VqaGR/jccTeLuQ/5RoqjbffM2J0TXBwljMcYY8+PYk24O5JbVb0
rlhmxBko2t1AKQJPhukjRjx/e1Yhmm//w7fYb+xM6HYbjBvIyu0zCFS5pQV4JTtPAcCegQcZ3AiH
JUa1iGDm2khN+kd+L6g1XpbgH89u1o2suEr0O0d5+3zJL5r1QutvQmjypoQEuWcI492O3xFAtdAA
ANFQ19927/AOSYhF8EVCnyRFnYZFpes2W4R7gOuHUgtIceRfGnN+JAbUdFnXGBj8wS20O/hw6hJN
UkvJ+InlBH9WBXeqrT364qU0Bcio7a1NnhabcpymieCPYU/jwp/cs+K9GPjDiL0z5cwuFft2EdEP
CuM6lwh+CMEVvSJDFG1kuo6XHB569AtBf1c02GMIq8eSe1ubncYvB4AKgbvS37vxydStEGZwrpTt
F9FlOaheVJK4fx3DuKOYS2ay0hyGgVAtJj9hHuCuFP8DoFwJVuQXNdr+ta1jlfZRM644TcYZKa3q
dLr8eEgKrFlup8f/TJT7P6vZ7IcsGr0At011jHYqVpbvGEJxxaoJMjSEmEuFhwby5ZqHHrxlkqOR
2bxHgHAkMG50mpAECyG0CspNvxUUI1PIOhVNWKdnELdlOg18uLGVuP6XrWDlSuMrG2+ZL0Vcjiax
WIrkMHiqVEPwMfjPNgIgwlhXEh8LJsv52zdvOjPPbNHKkdilhUk7dEzvHik+XjvZw/d6aujJzT7n
yK/0VPHpIhsXWHeU34uorLCMCsdu2DsCMlV1oqN+51zCfGJ4cZ7Pf3RGhnMlqddBdsOxo5e2KkPf
nnIIXM+Vb5V1KMv3f7KPkJsXiqY+pQdaHK8ZzTuJEpXCd+Es+KCJx73K+eyz4a6rYC4NGxUW2C7r
jYMt6FSAzS6cZoUSAE/0WoRNOGs9QpAG0lpDLt1cuap2o9hGB520wS8rWIBb3BiVbQt0F0VAD9Jd
x6m/DN4CwTK7BKe7xUIYHD8ekOnNU6qttWe1SfwQLJIsbok4MnigwmEiuBoc3w/i33nAgxvsTiwo
wRDDKuNFh2TfwJLWaKhhbGWEkPHd9ESdc6wp1haMXHXx5AmtCobcQU8NTzz9FzWsX2oRT6MeuxiL
+Cz5f38EmGMQFDlnUw9PN/KKesU80n0hK+mT47HU+Kkl7qnd+ndBUbnMSysYJocM7OMIqK9OkCE3
qbP1ArCmuclYBcg7THWrgkVghiZWTFX2K5hC3Eub9q831FOtEN/9SpGT0r8burhVFLbsX2yeHEH6
jgeY3o1jXwFub88xpb/6y/CsuOmMGFfT5+MTQuvMQogoyK1h4ZLYDyUtUy5ESonMrELmBIJamz28
EPNU0Hs1jzm7q4OlijCUHYMHzOcHfA7f1f3d6ca8fGxLstcRWtTS9GHCC7bq2Pi9Y2p/qgJ0ZsQt
omPuhdOddCTYH1vfGb6Mj/t2Ov4p69Q1KvXGMtT/0kY0Rig4mBMndqVY2bBN4PvjWK+at3ZYaWBY
Moyd6B31AQ1/LNbc6Jll8Jj2AHKJhqoEtAokVw6+KlJjgV8BkE5PXlQA0/hpWui7r0i4aeUPvKdO
RD7ie7GXBxhTQDcUrke/pnZtWBVHOd2MrMhmjmKU/CzjuiSo9pb/FUu3lbL+HvZhHuatrVfaTDQ5
9xB+T2iLUfetge0wvkDEMT0Ke2cRzl9iT6F+joay1xNBoDrcGmrvoOdbQiH+1IW+slRIzAKegq+h
fdu+j5pWRD+XrEH4T8aCV6LEM8VF8xG0xDaic0NSMJBXbhP98GWZwM2tUspPHxtwaBqSIxviD1cV
QxUmLGn/NUTew6KPR6IFVir653RCcd6CK/WgY0hyQBc0mIMXq0juSOjw3nHMlej2fL+TQ0JwB8D0
amYml3e0pbOHdlqypn84yrwov+Cug0rbFVjBoq6NEd5LmhNWm1xhmiBVxLVabbeNeuyyqvHcyGxL
jzs1+KDzApNEpQ/droEvLKJQVWToCuBS6C6afD4q1QCWFPa965MTttzLLeZdLyN6UDK94HXT4WoJ
fNOoz/zNaIVPjQ5vNEGHYIl6d5uY/sm4GpG2W+Whe3nobBCTB8dD0RVWiYyE/nwVekMffPsOArDE
uxbRi6XYKyPP/PNaDb6cwqRdOZhSXSHKQoKcjZDFGJJxC0RToQoR+Xy98ofRnO8StKQVW9ZMZ5sU
DMGQqUfjylHI9WwE6NbH3ly/mdZ/dplZIL1oJx082q71/e0Q9yHDd2VHpOWFvkZwzAv0VQaIsvKG
xwDHNfHhkZswShKrl/GCMrLl3LT8+Wn0E+8nLsWkrss6fna41ttRsEfpGxgaXv8gNxTpqgYrz4Y8
LLdeWpaZFN/cQQLZGF8pN0CJp/ikaQEE0iu51z5MR0Evm3eXdG8cPEL4Rd8QpRaCREhNfOAOMCe+
8TaHg3p8fpaNKd9/hCfcTD9K2WpITCOPJjp4IhBPpCboDjyVeZULoyu4UMKiyMpmqQyjQSoAwtty
D8EwW4vtftWjQdGyK+8tlMHTnE8JpiTaz33TRlVDwUUN2xd7BnyPb61Hpt2tS42UKS55jgnK6YsK
NayKuxYT/UKhAbdWZ4djUSrmRLzz4nqQICFdQi0kzVBESMsa1fA42k0yUnBO5buGJpmWPtZOQTqY
2erO8nLfTBmX8kb2O1r009BuH/y+KUHWdKWIaJW85xocS3Db1k/nSUKI1VQtbZsVFy5iJWEoGV10
txBC5W0OyW89t2+vj4lOJouSCSSmjdll38LlLqSgUzj+MW91dnTcraVipcb1SWMsBumnDpmIGdUd
SJYS+yVqTd8ETPSpaM4wrY2s1xS+OPdR0OZDUFKF+Gc/fkwvG1RUsGEL/HBeRdWklFNd3lqK2s+r
0LyoIke5NkB6KklqNzzlNIb2ah860xX9SyEof8WzpPdDdUMYePGNRWV8LZXGphuiK3QcGf2z+nu/
wpzgFep50kcGAkn+vQrSLDhBtI5TUJ7yK0QG7IdwdUILzmMdiePlpQXaX67m70MXd4oXe+5kAeL4
voN0/LkeFGQcUOLNBT0eJRHq+89JJkZxz4rHuYPXg2X0ZQbE7XuRxUTWYrX1VpNwOiSubwvSXeul
VCsTUd6Gh1RPy4pEfWBIlwGo9rrjnl015FpMg7eMOoRqWQan9yvhd1coBqG5p2PzwM1rb+/4/V4m
308tRBY2H95YNoc/cVAFCSw7seTO8cqO8thoDTIQiE9deP7KopVeFzCoD7iNX4FdbIE2pGo5JPiO
vLeT5VYnz8EhdZHrCaAcAS+1+P0ZDnlcl2Bua8a+d3em9HBGBMd3xkEjRBA6goTydpP5dx79UK1x
5EPy5hgDBYnRaCGaFduVU1lC2bpstJFeDzJ/SaTl/sFFPOusJBkrLLRXQdTg+ik4aIotIpU1NgAY
tg9gYYy8zW3B2ZgL5HReOO+dH8trAgOps/MClqOKvJ9py1efyEu4NNDLEUjGpBiSXslBsR6iQIxT
0o4wkdpcG5r9N+RoB+NagZ8i43nB8fKxK9zbxT1/C6TRsTdbjjlQpPgITuJtVf7g3povKHOnfzhs
IhRO+nMpdGmAFF3gPyaMY68JI5rZRhBFpelFulLpwuQ3pIHS5Hhr6Q00dNWr3XyeEBsZZhMPb7yc
R/OEwUKixuF70gcTJjOk51e6IE4PUdNnUZXQ9WF537kYV8vucKLFR/01yDyiHTueacrxSBTDkkAT
fLNRiFodp/Yq990HTYbnMI4ls4Q+tRIKlCob35I9+awIU7HUEXVGsZZVM71w5tpaO3z4al3PkNBx
Il/tpg78ZTtySh3gF5vGS1ulKUWKR8niF4o39Jb2yGFU8pgIQpXMO78Y7k+wB48cXSBY/xekHbW+
QMi79RW0IlJ8upMGU65ZzT4XWRetvwjYnqbbEmWyd4PJXMpXYQv8xzis9Lrs6dRuibgtqPrOhVcC
FL4B/VogaA2oPZU0M9FP29RQwS8DW5UH6GrOrFPapl+t7J8yzhMn6wbdlWzUsHGEeEplqx/oXVE6
CoLsUEypFutxXA+vwKZmGnLI93NPGSsA9iCtYeG9BylV5m8LcFk3+vf7OzGitkji7I4V63ZjGxnr
DJDmPJ8mT4dg8ZCotUCI+DiFa6m9n0H5iMKWu8p3qN1dvUtny5rontJiKttJzPbdrhfXOg4+ZVZK
v8zWn2guQ6APJ8hFaXDShQyDlErhfCSn+az7eYedPynEW1EF6SPnbTHjOR5J0jZ1CQFqZuU7pE2B
STRaXRFY9y7yV4wsSAxO7zqJPXVoqpg4T2ZiLAZPF10FKBiJJx2TCYX81HiqxQgxC0TVXO/p/Si0
g2CULFm+kRShdEndYuBfwVR/kvayGbGm9fVJbaPBLlVutbp+qFo9WgWrjSHyuD3EMwuUXS6IaDdT
guLI7wzzVj2GGQwth3Xga/oCQwY6tRK3iFSeaE6wrrNoJxExJGmKog0QDc0+mq/54jo3vfEKkYR/
DKmUpLJOwtXnKqa7AdkBnOV6iCzF8anpAdLTdxig8ovEylFR1ddipxNZaR3pt3VD3Fwe+4xVmiUq
m+++AzanRiTbA9363tLVP3UqG8EblgKzRu3bdburlniQCbBc9goA4/M2Dg2Fey5eTriIb7m6x+Rl
R9RSMglNItpbd0m2yv4Va7PR+IFxcqWOVfPYCBmarVXhqK7ijMsHO2X/FR4cq7UvXYMTZe/JLqFl
ELXS7/iwk2DozdCHBXjTXqSUtVRXZn7pkfnaMnrWhfzEJEnyY89VH+leX5tdIvLA28yVNhZdJ4WQ
BRVB3XkWX653Dbkc5CdkvgaWeK22tV4K+WDkHVCEXks8iynH81IlA+o9sthAFgOHqpQWElKajXxp
rbwm7O7qb/T3uHGLdYPQQsvNabvGkU7xVlG6K+OXzUWPa7gdyTACitzpGne2KnFsbmBZr/F3GY5O
YyYbsG3YaGI+tfcJjgpqm9/ejzv4nqwU3tfqNDxl2mdT2uNfSaB3pBAjG/rTsVNw6rtHv3mw1w9U
9bXdq9aMxGSMBPfoSIgxu0HjgxSs5bETTGQCTOXJZgM3VVEy+RAeXTUkRDrQg4EVpqQ1Ht/Gb9/e
8SZ/tbBTLfkv/RiNrZ39dW0ZCgXYnCLdss0HnZfQNmxQGnl/fEUzijCgIoI5CTMjXrr3Xix1mfZd
7yg6S7gKQPycUbAL/mFh+Vz0Acj5LifzEIZcqpRTapCjFn+3WYyP498nQ+zhmccIPVZBapZhflir
gqMUkxhDMuBnUN+FRQHFLrjDST6HpndilA/FFtY1mNB4nfuWsqDMA8b6kzQmicEg8DpfAbm65y0h
qa2wKrrZ7r+xRgXql5f+ZNqCRo3Kk2uZaQb4y2a7EFms7ShRtoiaoIy2z2Hx2s4gM7yErq4ta9XN
PbDx/szICermAx5XzFOvJktASw1b3RMMFqvhmZ4O3Zs6nsw+DLGEpMLFTgUuHAqHkfDSpsWk7yR3
Gf4pyzYsfpoOb6sb8V5ZScrxZLCJjf7cI3ZHB6rSGf95s6ldx6Yg251ZQDXb/zPj1zW8kNNy+bXm
LDKGVeNQyZb+0br87QGpoPIakw+SabGrGVCNKFnFMIsyVtF3qRmVrPflhFCSOjILsJv5kPiotcJz
CG5d2jofVWgOOREuU3XODeNQ6LqBX3lElkdOul9t1XPTnzGGi8cK0YzzdP1OavcgrR/jrFQfvFqa
80Kkl5CUCdILvJaaD6nSyT48FGpTJa7nuouXYzxx5YW3PAl/GxuxsZyhSKVGlQLnR7C2K3v+atko
o8MvMc/ylpHFltBUwj3z8+P5TuanUmNIxgi2vYQ/3B3MnlV69Ni0PoQwPpJVatke2T/h7UzmAFkH
nMNqJgKKyUO7y7/94zwa8iedIDr324YAUtXSDHVcOYiz5Qhs6ZefoogyMil1OI3/yrI2Ma0lyBMJ
DKyRIw9WcfSC69KQoj3fno3DNvBCzvzctq6aZwc0Zsxp9E/qkLIsWkq5x/xu/6itgTCIzRAE7jHn
eeu9cFUdz3jXh1G62RxQqqMUblYJbE5LgP5Hgy3Y9HeHNwX5GXtXH9ZSUh5a3q6KRWPAM6OS3FOd
w8igYH5fz0ZA5fbSUttya73TI///OR4JgqaMm6k0/ffA9OJiV13qP9wRVPSu64PBGqBvRyROlU9r
rHNYMDjMHnGj90ymxbqYvjM5Zwt/x0JqpMT7qYbdUbN9hr5+c1P4tLomyJj2EtHLTY736qxc56AR
KAnZ1RAsF2eM62FEQIAq5+wOCOq1do+D4gMZ7qjGbX616VDvnRjnMsJFejE7B6oO8iRc81+ySKQ7
0NvzzYa9CF4i6vQPUUaaF+C9ERrWwcMvwx9/rnFxw1Osj9M6LQVAziKTtFPHFvsJN6dDYpae2ePM
nMMmgCRb8oZ1LurM2Qw6oSMcZRXbyj0nG7AACgJAb/ZKZNSrkB5zfHI2QJt2Y6KSO+f+EPAgn2AR
5fZYG5Hz6GhnmUZo05eHV8Yz/+I4TqtNcDY+KhNJv5eZT7uLuxilkcfvzfvbSklbUvbne+9gzDyR
6r/fv1J6RKNGvslv5ifRmKLMYX1oUU6YSyPmc6dHxol8UToXjd+NoNf9NRBSKPgoTv2vcQagtrx5
SvVJrP06MQ39VpWwjGFRipD9XAtm7p1AKrOWZfaVlp2xIimiijLuoP6iAM1Paj6SHmXxUnX3/+PK
iglVD0gJ+hIONXKGIxYfzpwPcM+177rciLbzksDQbHpZFB+WJkNulltVTAI0jnznb4zVRiC2N63Q
EZ+iSwe/cVi4Z/nJUNLjc0f+TyL6+C0w7Dheuv6ApXpWrcU9gV/Lg3vOSAEaIx2pr01tRNkg22CV
D5mLCA9+P5D091w4g0SCQxSHXz0wPc19vOLx6gkA8Pok02xRLp0wSmRSpCA4x5RG+02txEXGu8hj
ZSH+EzlcicrNWw3MsQdUrj1hbB4duStQOs5yGEi2+bewTQyjjXjeogOzwKf8xPfodUNV9MlnYPNQ
ecEp370GrMRDz1hdSmAyKrO1HRAXm3XYGxoQFg4lkXbrgmgGmp3eb+V8c2h7MV4+8SwOk9eaqI5N
9YtcXg7vWimyGGNNR4Lxm57J1SiVpJHRTOL6mM1zw64RLf6hXksnqnnW9hFc9+7kIUhSYZGIfpyh
7scBZxrufIiyf99Q6gYLO6zU2mdB1AKgNHkWYklC5zl4eaQM1GCLqVsVqwQMvc0WIpAqzOZ58tqX
KB5XRxiSx/l1HeeRIw47nlXSfYHJ4pvu7cl3OzAUrTtD+t3o5rToVDLvof6uk29csxdS+lCQr3Fk
pQ1eJGwTYKBBd1TkeSgJxsZbL1aPMwpEAc+A68mQBPIKZjSr9E/WuElN279btN+izukc1zBivydR
XWtZTjwkodWze9zfAdyhRFs4CWsbtBBxJr2P0zGPFIscXke1OhoW6cZrUERvEfp0uxvWCsDGukx4
s91n9OWLSonGzWVGEIdLf7A4og5UXi1dR2nQEtEgH7edJB56h332x4HkpMFHp8VvQgp5l5SUpypQ
BDf9tmd5L0dGuIeb2KQ7H3ebAD+UzsomtYOrxvZgGnpnY92Eh00riwcZYEXi8liE2GPxQira/uJ+
bADN66A46IVXD0OwayDwTlX0TZWiCYmd3DuUTBtDvqdnF1v7nMj1FHjw64+HPtc4ZQVv9H8vvg7X
r4jP1VOhmeAfw/EI6FXv4nRz5gvbCM28xxw7nVnfAxF5ffTcC7QgLylfYESaea0njaDso8uh2OAY
qKz4YaCX9s2/D2ZoROq7sw8VO161Q1x/x3p0kUrGyif4ImD7vpjmqXCD7HgTInGVjQHgqC5ovGVm
OuXdzJOY7VpeCYAndZXUIR0Rkd5pHXLFsXpxO3ufoe7mHFl1aWuyjkRJbOdH4yH5gXRiWTqkp0bq
0YvNmjrZ6ztH8vxXZOm7Rnj0uuqeCksM0RgpVFlI29F50PlOI64VA5LJKeZ29tQSQwvsdHecCrQN
C19pdJEO6H0YZ+kA7h9T+wxDQOWcShO6u8jxsvNS01kKTa5iTRxA4iqth2uSNWZw4YOs/L8yu1g3
JonTuGQcRWZa4JmvtFklyLLW/GEC4wZe9rnhRW7Vcha4mTyxqMF2OI/6dinx4ajaKGW2m5Q70k2D
7Yq42fX5Wv4WwaQjz9fTVT8GIyd5bF/YAF5Ht8T01jM3LvbeW2OAQvt9LgCL6s9W/YuvSGmQIwQF
9ROmaovDUfLmiRRrnW49srhCqViChp55TlqscMYSUIAf3njzqk2pLcUzakEJHGlkmIO/1ngDuGm4
Krt43esZzWkTvoQiE90RZG67M7SO2aYK2on92trmrIPTjef1lxa1xxVxcIh6ZqXqQWbBv4OhWRq3
qByX1Wli8VlR2Q7oQTYZqBMyLo2ZtKev4XQFPnqjL6i5WulQ6httq+suiBLulU8Lr79ITC0DxKwm
abkUYKK2DQe8FrVhFkvYPBwEau8SFN+qwookThnEsPVsLgbrRYzNHdr5M3e2pyhj3PpH88cFlg+N
qCnOsvDeO1bNxSpOmQ+vK2G3lHMvFlWoMii7ER4GUZ++sQT3s5uwNAw4Ag5/kUAdxa2/jAIaKLdw
sjJ9VNTwKUGHXyYmMq1mw4zcrv5xXF/rC5Gxffat73SFxQRICuqAO72DO4gAVHIZY/eZ9scM2Ah5
x2ASq+cIhNUALAxNI/F+F/MW1G+qlWWQpV8qzSw3TlPxktF665ZQjRbE735AGr1pifrAukv9dcms
WeCuh/4V2OKN44jLco02zSI8ArTvu8SeTZlxm+IW5ZBxHlG+MC4dfwaAu3mWYCjayM1e6l8WxR9I
nWsMuHu33HB7qc8N/YCg2OROkZTSTJmmOd0x80jVIMOKjQzzrS09ANQeHnxKucNyO+ncMIGl1Yqv
aC105hBwUruDGT3ZZCkt//qKbhBH9uDrYBOTTyp/y1IRLVbUPGg8ms0hjojAWxW4nNdL3dt7Mqsp
OgUjyyD7ZSkiPCKAcaMNx0hcpa2FbMSfd2aPfgLMwxAhb2S7JYnbyrNvtf2yMKEP3GXuOIuLwIrB
jEeAHEQyQy3B811AhLPTOKEGwQzF8AK0xcH3BaHoR2UHu/c6l2GwFglhhsJW15DLkFoMTJ61cVft
wZ3Afu2pvio9srYLd980cRDN4L/piKSPoJyHfPQiPhv4QtK1fF4dpD2QaixwH/kb03Zj00PTW8PE
nOKusKeNVK/AUueWAwCB7swBNSKlOnRhx4jH8j9N27kTc8cM/kc5aNEd+KQmqf0zuaT9FlbhmWGs
mMwxG1VDF7nI+asrwVoJy3UF+ldqiySPmfhqPWTYsC3Pt/rsHBkIozpjScY5USx783r1CQoflMFx
5X2MJQsL/sWWRegECxa/BvFMkw5f+ElpFH1JvaCSo48sQKLIrTr32tKmZa6yKExTJePrE+OSvjQV
VPeWE40pvRJMhDIbgLb7LbBib1MIubf0Vm0T2qctL3Zdk2voig/OLxtWnaKWk1atYFpKyNh7W5hQ
lxeEfl0VELxUe2AQudMgzPItlGCjbYp4av+dR+x3hnsjCRlF9jgW0KOmBtIonD4+tqSShQYoA9Jt
ccAuQSo5w5GpxrWvJORCHU4H0qrrrAE020XpMn9+aTBhojKp7JOoo6XB6oQ7JVwMWgKAVkPeHDBR
7V7/U7U3jtqyyeP3EpPiqjdACKa+pytXYmZ6X1vp/SvJYSmw/I71LIj1X5WsF641OqbhfICp48ok
U0LfIr1f/nLdGp5H8NVXCD2y6G2TxDZZz9WNan5gTL6V7vnla/EZBh0G7GqCObzpHSsB9fFUZ1R8
HvMJAlamSO6erB39B/m8VDOyDHSYPiO6cb8cWvtsVSQhHX7/06jZmdQuptkkjl4AnexKY4LznE6X
wfLiF3CBJzpBPKsGqye/bGiHSvwEECEtMqvqIJ3KK1Z1Ng/RYcZWvzSIyTzUiM+/kvIVV9BPxykJ
lWKRQReNuAVLY8oFIzU6OnIL/75QqgzznNMWBmwiE4qDaWl4t5Tqm91yxVB9F1ZfA+F31U1UQZQT
3oDofuGsfZ1PN4mOyY1RqxaYOptvBHxR78BakLaO/d2xWgONJWT7XP17Aj6aGbN0KafLK/VzzURS
cSqplPgLuXauMsL5GishXZ/VMiX3Ig4b6vFfoEy8BV4r4TtLRnyp7HCROtbRJEibXRWtOFJbF6jt
+8N1D6Flgl5hPZvTTbEP/l2v6oO2QIgr6UmHj7OeMUzed5oBQRceC/BAbm6uG8J1dykXDidT6WdA
/ZFW1TEn2T3Stp1nRJ3cFsOgbByD1mrzxYPT+NmGi0KetDpgOvG/VOcLliJaRtr2LPki4fPLADth
Ho1fRE+MsaPSh0nrZZ5NM8s9G5qZFNMXvKd4N8xItG3xpW5V0h7d8usPsIGDmbJ3iSpZWoLqo6kp
MXheW9QWNtKIJ09QeOCJQ7K0N4bCj2c9gY0LgkrmoNAmJZfSfk03p1PFa0MzYsCLVpPqc0K0gGSm
cu8U/vRYTow7Z7zb+OVexG/ovVfI/Qg8na5Z+9Ax7hYhUgBkxpW3uh7sxX21jxC9aY4jb2dDcNfH
tdDLxGTFszxwZ8fFn47aQpSHuM2JRHdwIPhekWjOwjJMgD21SorD0BgfvVLZgQVI4+lQj7Mq75eX
h1hszUuiO9G/fu30sZH7BmVzdEdo53ufEqRYLexYgFW34/3XcBKDrEik822UwwXeNFz9v+ipExWC
0ncW0jHGyMK3gUueJC7oIvzuinjB6VSyJrOVuiUpB8HZ8XXDsKMKEFfGiD/1sDmknIiI57LpUBzH
DyboTH0pa8pZsS5YSLiJhbQPr46VFwawVjFr1jC/OMm3b/AdM9kaZOra9+G++bviZbXrdwPXYbwV
UakS2+8Ha4kiifoOfCjCXDGUUye9h5Np8JDipBFgGRB1b0gMt0H0WvG5PGFY3TXhp+ED6ZCF5s5/
D2d4srK2CwgexMVw+URKwgMpTFptWEOb37Z7mO8fUKFUD+vmVH1MPphtpqh5YhNPMJp97xldKta3
wJBDJeTXH+oEn9Le4ObGHsbJoIvgL2Z9lu0JcW1wUSGeXMI4ovhTtRdx6ZYsIp+4gIGxSC5o016V
5d0sJRZmih4NzqZtLCuPUUOZUPcrEskLHJt9c/JtP4GQ7i06A2j+vHXYM0lVRaLNCVOEFeWxI42c
pozk443gpI45KyFiYFcC51lmH8G2bo8XJU7ZZ1JEi5ElObdpxLpJTuu23AghQjajFC1nP6E0m/tz
WrPux45xonK0zwtz2xbzPXQgDh/LPDDpUSAWjmPSx1XabVeRQZh3PH/NiC7RHIyp+p556eGzsEm8
MrtrUp7Oux0H8S8rhvGIVC+O77wHoMV9vwDYSifMCzn6Ok2g8xwQSb9tjh2o3IraZELYUSWw3O+t
c8M/OK0Tp1gk8QC/ZQTRMbSh7E5FejBqW5q0xDNp00yp+WwYNhsRf2JehBzqhICFkzktmw0Rjdbb
wm2exEHySAyIkQ/wn+gC9H+MmXg3Le/dO4R6ICawGJRsC+w3drzJf02peHJJPc/g8EqNPb1Vhy4P
z02j5V43J9hR55So9yWHzu+WC+k7Y8whITKZ/Jblp6l1izEO4DqjSu0pO/E7/9Rw+L/k2Tr5U1sH
bAyF6Gn+m4IYQgiRcFs8EXpUFNQMjq3tZLoXN8GpKP9QF3WsUQwPBk6cCz7WRbcZW/kMQwZsUMNJ
Idk5ZX5CckoHhjot2xeoRkQsOnC/Kov7buTC+fsy/FZk2oRjJYBnF2HAtyADOZhDahl0dRdgoN4y
IZ7lKICic/h3kRHjKfr/n3HdL4z0nPJOw3Z8R/Sd59AV3Z0HQxjtCbZ+MQkAWGJOE5tpd/Ir0MgZ
2YmOSWNE7H4qPNbM9GCN3cLedgifKdyh8oTLY6SHcpnl1aqHrJVeUz0NSW73k/oex7YNb3LbKAua
kGJZdynSWA7/mvEcOWBev3oClXyjW4vfAYgrp2aYnRrIBp9TGY1sc7Hw6zE18Hl/27XP1jUDfcfV
RBJldPEZqLNeCsSkOeC0vDTfGXtSgmQqY1COZrGggq8oSPiTKTAbEaK1zYYDAWfVdhSZZ3/T06dl
gzrzpkpUcELOud+fzAzxfQYhb6Uuk8MXTK/QGK4xagxIqSc74jt3WNf4vJmMzyVr09CETuz1iPpn
nBDLvAwuHJr7n4niQW99jwmLSGRe7Iahk+/b/3wWjseiieUl47sJaP1XXsuFFYh42maH19eOagIT
HvKAF+z/Jg7D+GlJevOxzG9iqSAdhMzFV/FuWV6JlMc4II4ZwuvMFJM0AyHETzvJQ0GxwacaUbfJ
Ck1caD5RiVr6L1zlvFcsfZ0kBxyMhJ8Ivbc0rBjyhl0v3ZQMWK0HxciXPEnsTve47SlMeLZGERdN
ztxHoBJ7ZRhooozVTc5Ls+IaxEDwaYYVaw5RA9x49iLaqophGyNib6PVwmZ230xm4+HlNxoJ/prS
D+gKMTgmywoUWB17NSrTBi/uhp4b30RCUsa+ydNJVTeymmMie8s1ZKMtEIiyRVeWMHurjzO214Yq
ZOF89Pah5Rg3ybS+BQlq9eCJvIjCPcXEfe3tTvHFrkgx8yfpuEg5AiE6Jzq06nCwtoQ+EPM2LeEd
9Lzxsggr+ZTuRTpmA8QAnj1LuxjZY9CyyXm1dBvhqhtuiIqTx9kzm99vw8wDE8B6zVvfIo/cCbrh
jqjeSf7LTo43nn7N9Mu+dl5Xz3w0Q64j1RBc/MAnASa3fiicpifn7iWVYe/DNe3+ESzatQDAiHqR
rWOM7M5JBrndwk7naphzOrOuoWkOESVko2GAvthHd/rQsxfeYhKlmn9bKm+jZiYPkawQaC/zyIV5
lRkNoEF2rD3pUTU7LKeJYZDuyBKCASNigqj1yYWpOYqpzepPV6W7aSaSp5RqhNW1bBOKOFVxiNa1
uwnPltzAihHzCD487NlAYKwylXHzcHbbMH2BbFsoguOwc7/ijLdQSYT/i7+8rPXsuhIqUkxdQb3W
5GA6sFWuQCpcEwTnfE7TI2nLJq5/xOdJycqTWKJ0TAGStp5+E7LMaAe7NewFjn9PyEs+QQiCmNHC
ajSuE8uTwqpDdfB+N4nK+InJQzEbvDviU60qaf1FZgIiIvUm9TtxGkVFEaRJ1obbqZzhp+M55+Oy
7rwCmmCb0OwgyAvLlswQwRNzDMDGPbez9YSrmGma4LZVbRlnQ4qphTEnjK91P475G6Wg76y/2nTX
YH5nRzWq3znokFE4dzzkFhcfSV3BfDvfo0IV+t5w5DbvUDdf7VCP6394itoFoI5a6Vg4Y0eODNWX
rw8+FgUJG/Pv1XSErgxMTY6V0llGWD689+XqiGnanRMfnjxzmFhh7pUmK4hbV4g5ZU039jP0/eK8
wb6Wr8czqXy1ZpM+qtEoPCO50lwst5r5dV3HxgWksZqG02Q33Rr721xIulQ3660l07ZEOHjSpz1H
r8Koz9FiSkwUs7p827eStL3Ni4OzRDHbFkA+HSI/VxDmuepcVrdFpP6ggolOjzPVLT7haxg31N6P
9heUrVEqen4kNSyW2v/hBsAd9Jxe98d0gtlWRhCyVuP4Uvc2mScZjWJdsBA2ijodaIV95qDBfKH2
NudM9ewkUIZNIadNRy45eL4oRo16FbGFrTT/oVfTJTwF1T2cIcQyqJ7de5j7VKmuU3JTvD8+ewVq
0CpHA7R7HWL+lAcLNK3MMgM29GfjpYY+Qp6OdF6bENkelIGvOBHr42XJnOhoxzOE6BSzb2NF9Cyl
6DnKWNb8xxoYjMWHKSl0RCq2pKxaUEfzzyFh1zyUuYOF+PBc1LT3b6ZZh+GHGUwJIUvs5KwG1p+J
3KD0geMMrfJPMaXueDKUG4mAdYCIN8H9OXhkoen0FVzBdBRodYjp6cetUToW+NMdwhVOtiv8R5iy
fmEef0TXCbIMPhUp4/eeq+XyovxFXbCCtXh6hp5YDxbMwuBsXZwVzAWzms77oEX0RF0CScze6iUQ
gzNQvcp8yOnoFuKlxSIArchTX3U4Azr5CmbVqywTkR20tVecoMC4AGeurUE43SlT2vobOp+4LH9D
biiIxT/oMwIf8cpb7/ZX2kmC5MLmbzRk+rOyTG66SCpspIiqA6bS6lVAa08DGs7XbEnL4F1jMVI5
5aRBZ8Kpi+TcdXEctKUDutSl42Ob1TYQp721eUfbHK/b8MB4cCDw++pqooJqwIzbyueAgFxRJDMy
gxaoYFSNFKOiYQ9gkqYwsVBd0clituUzfJ9lnNw88wfWw1SME6yF2zX7IsqIJZ0TdLVb0oZRRw8c
YLi1O75zA1DThp7Jn8yQVAC9p4BZLg28x4M/TZBmQzoNPAfTFefttUMjH66rp41Sj5oVI1naMR9s
R1ZD6xdyvdM4JLo8Rpzk42WswFGMVa2axxvCF0Lgkr9TVeOjKJ8c0VP0OVgvLo36XjRIr5lJb7Wy
IcqOqD9zRPf1bnrxP9HXzoor6LmGBSp33iEUoY91BVKJvKJhZV7DcDwUPlMPX7etL5yu8TzD0kz0
MaXZV12zlvw4P3cXma1Q+dih4yhU9nuLGw9dwMsWeB2AuSlPN4CIRq5w1kAnxoD1wQgkqHOOYoYo
ojEB9tYNKSqgjiGWdmqwfFbIr/gfYsyKGES0r0jPSg3ghyMQHvgYiIozFVmvUIDawErJ5yjrZGmY
LSdjX8QYGve1gps1QAt2qpdXAc5S6z/YYQyfkNyx6Wg//xB/Lud1KjCBstkmrwdxOC5+AhMl5hJy
SZEooqvZQgMOm44OBVRDarZDJbE3fEyQb6pPRP3KZprqlYAC8EkSzrlruJ0NB4vyJ0aiBL0P/oaE
YxDjIjxeCjt9sszTy1uO/RRcL56An0zeL//0iqyaW45DYAwCgUMumndmcv7A16H+nxMGrD7ph0w3
GxD/wy8932x+Hj9fBQMy6IdgcnzVvlxBehOvIE4wXgbM1v+Z5F5OjIItV9PvSBioYLgliDw3yn3T
EpiOtIqBT/dcSKBYmsoEvCIpXHWcVVouc30Hg/PdJozsnsB9P5KnnL/h+dAeFxsZDAnU6B8M7k3k
YVaeJ0L6GA6OzvNw474FT+G/JY/xnhidXpSncRTwkK250/uKoU3A5nEvQohH9RXIX4C3kWu87Jx+
2CCbMV9td64H+q2QkuR4JBHIApXOlYMX6gwYyH6vD31O9Keik3nF8iUWTnbG6GDVTOOhIUMH2ZW7
5/yoUdxfsUkl0bftomyCV2DM3P7S1HLx8ILPZRYPoTvak9EMOa1TdYpIdxBzFstpwjbqIAkFL6OI
U1tjQwtYMHCQGPgtjvu85pTa23dfY31Kanp+5am2y6vJrQF+YMgsXo1AFlRo46xvY2yEf97u7V8h
BqnFnRv8qxf5cohZlbOX9qG4mfPjw7/FJVJUnpwxJY+pldHjIVgfyqBxKSQwEihyN/61L4wg69Cb
FNDKjx/x9Jumd+yqrZHzevtgkrREaVxHBbe72ZCJXZscgpDINRKkWbsFTjZef4sv+a0KGtQDX1dM
quLN0aOYyFOr7L+Q1EdXtaNGJHVCdlrAqZ6BTZ98Mg8dKWlRkTbWqjgutT2k/YWlCSOo7rAxjlW9
kbfb+VDzB2ecwydVm20i/6nnjppPJVys2D1xktM3Jh0hy3TcSf/QcrJGrDRij7zNt6qSUFQmgez3
WOAHsXI4uTVxGHwZZDt+eW0lFS8UWbnh1bThUe2+VXhtVt4Gel+qunovUmfg/fSriaZ/2pVOWjxS
1+LjkbQY5DF0F8aWelRMpH+d/nO6UVhPq9gyCCTb+rZD82fbzo29e8tJgN/xJI5hyw7/i02KMe0K
tvdtdJKC21lP7nL0k31fqCeFhbr6eb95WwGMqlm8KbAJRBpJmsVaHc59Tvo2N0mJ1IgyS53LUf6u
8rpTzeYW2bkRBJcBvlyutTtZDSy1wYUuuaYSGDqBI1jJHxwxvd/KAipmuzgAlsC25bNuoGYnrVxP
nfhRcS7qB5QU2r4ED5q+K3jqKrDYAEKBtFZHHwKhjwam/caWjR3gFDEW8+/cSihziUktOgURCXGT
NjbcTOtNbHQCctAAxrrLZx0iqRtmTxdyjvFwk4ChrG4C7A87b6fUilQiGWSRrY2GBBWhzqOHcwok
Ivr8rIlippjMHGaz1sWeWABuGZWjMMOVpn53XiNHkTc60j3PI9aw/GMFiy+OiIj7MQ799FauQsus
9wX2hvOgWGYNaJt4WomPTfX37leV/+GzwNZCcQBD1lAWp71MAsNqvFJ2bvCaJM6cbcLF9C2H0PkT
DENLkjtjmUl2oWYbeoBZ8hNw6WoNZIS651XYZZkzsiIrGWJICzzY+6vTiID8axVmTojiXBcgcFzZ
6Qp8EPWkr+ptDRcxvnhDqnr40PH3LKXYXbKMOSZ8F7cgK1pCoF9dxD1Z2V1fy8nJlCoYSKQ3SjKg
pgeUNRkY4cnXhZ3XF0/ce2Wa9iUaryXKPUxkyrCUs5UTrcWNX4FwPkLtSrFVSGdZFRq0oEfPkN25
2k2I5vEe7/UbYsGGou71/B+nSLg6Wm7/xVz3JhMcgQt2uVTq5cOs12ifEju95WU9K7SzFS2VP/WV
rxxIPdEuoyWl49F5lc9WF5YtkPRmDn7aTt1WQL2+gjDUHmlFYPBHYWqr01+ySfmNOTefsGsbAEkL
0oyr1ayokP8TEgzrcLgYNUjV8CPNG1ZFOxIwZuYYfZL8E0Sw/tON1Qeq+BYjpKeWMD/9V2jSrPIO
lkqXJHe+47WdeViYWPWb3P3HTPg4gdYhTTZEAJSspHQZPg2xkyww2ETwHTpO18Z3QC4fwDahxp6p
giGuTGkG0BEF1DQ4HWU2GvY3BTPkeCuB/1N3Dg2FDKJ1Zyq0k3xLyr00E0iZ8TpMCMxoiKQgaZAZ
epFe9YCgVYOKHoUaDCBGV4aBpsN+gTzSNdiI8Mohwx4E98oTqVc+kHOD6pwMUPMirYxQoLlY7O6X
/qNFneJFuhn2YZTVMd0Go49QZdH/7bazn8naB+vHSZPHnMDx7vXYNkAgGNEzeAR7d/ra6fydSDrQ
EdQ3K8tPXK976WplTbx+ibba4lbSILIUgIhE70gW09Jnto36tIBAlTnQ75dzJWVn2ijMgzQL6bwR
j5zJ1C/kWdsn3frC2UHgw7rEFLuz3ZKjigFWGOf8QlpsMTwMixyloSQBvq+D2p7rkiq6XKuTZHMx
FbSYA92GBqYWolCuPZxEIHM5Wka/409rS8jLq693Yt716NJur1nWIZvDdBJxPL4u3rpTZGU1jT+t
Kiwy7cWmSS4FBATRBJdUiu/0zkj8Ptn4eVuzuyf5yr8TKC/MQfE5GU6Z9cDrW4NHKW4fj4LbPouH
nou6fPMG6WX1esmY1X7A6zScBxpjmj4nGNhj+Kpvh9vnGFr3YbNoqV+BzbJaQoUP9qraP6oqbXBQ
9Ay3W63Pey5b3eMCY4EYbtBo2fWGV3mkOylo2FxynGJqYUvbCcj5dIdvf9x1f0wkmPBLgHPy8b7x
QMOzxgCxuuRX6FUu1zDjeXOREZ+RA+p052CUuzPkZTyYdMBaR7sKtTGbRq6k/NEoUQ9Zg1WYT85a
Rdp2g9XthHRRDzCBZK+YCJI9fQp0QfHFVyWaTUSDN+vY3hPch7+c0vKDHMfux93d+YRhyDwsJLFk
mD5XHsAxuRyzsyVEDN+WN5/bmIpiKFiJr79HMc8LZf9YV8uyHsXMqwuGpxmTJ/G0pkSmAcFzsGFg
FXD0aBDvMsgI48kyVLRra9OfK1k12yBFCmGr0c59wVUOZXx6jOxhx29FZ8T5r23WJV814UCyyaVo
Vab8e7L31DxB+8NfpcCigdFFJ8pYxrbOHVBUuGf5IWzVl14dUHLL7Ru2IvkdIqNzewkWe1sn+uih
4QY4TdrDknUVImSbTxacbskOGQWc7A4l6bJcRboWTcYs95c+0bG+gGeCftJte8nB3KMqP9F4TQ/S
bxUCt/6KIbwyx/Dzy8kGbgP7+Xp5UDdieh4qO5BC0+syiTi2YPnd/UwhO1Ous8DLPrx3RRt3b2qL
fNsKhh/zab6mi/IH1yHfw0A3JJtQ9lC89cwJKxHTDhtxEf1DDSh7yv2gUqpSp5+WZ1BpPgzW6xoj
slw/ixOWhISAfjLDzQyfwbYeu2Kd+jZ4EDnlhh9jNEdxLSOSi4DYtL+xWstPOo9895gGjDvh+oSt
a2EsRRDEppOrmf/apfevlvlY6GXogWG7apnDFxEj11zXXn0ndGlxfyPvyiKwWjOrwEDe7YfNtWvV
UqIIx2izh6Z4y0TQfiiFbKJkdgfIAy8ES2iyHz/z/5Gle4Vm8GrIjLmfoRSJZ6nHkBB7Ah8fHmoj
44bx+5c4vC4e7NQ8/LcKbegja2pTpWNEgqDhUHWDmgVensCmIhTqFfEaDeV4D/BDDRdnKPgG87+q
wGMuE+PD9ooefmswh/3h/zR7OZ8yQexWNPPip+F8wjwkkewCGhfo/4IVHm+P0U8NF7ipPKFNfsSn
BcvzArcoUkAO+H0NReSWAkqSVP9PArD1D3TyFCxWDXu4YFg4EYyMZOD2OvDEde3OnnRw1ImrQgaJ
xIWoe8oPt9o69mR2e2W63RdoaZk1gvFUlZjgZsWDipO9MA7WCRWkyD7VNxi57EKlD3QXHQPEdGRA
dzJlv6zzo1jKCmmp9JZl/2PiYXaCSFJFHkHc7ZorwEhkoKij/ZHQucqbg75tnkBbGzAO2npdL/cY
eVcLGMRNZiZRrYpBkmrqkhX5dKAvE3moD+WsMxwW4/7/hJOm8sQQmiMbvw4Kx8k5To92yIhqEB6x
yg8iLTNUO1qWzhEQNAYeZLz6ZAyHzC8/s3fJcu0Edd2hr5sJG3Oc6Xh5Yr6YCkbqrCUDoTOAC24z
KZZtpM0Kvz8A7BfroL5nRXk4T26W70RLu1Lopiw75nEI81w9rNunHCZbMxerLyGbDzwb6M1opri2
pzzyPR/Xq+lwWpu2cnPcOf66gbosKb1s3RXBy+c3zvuUsLDf/y4/4ab40hTDLyAR1eQqAaYOjkDe
/ps7pkxJPk/pAqq+WvOMR6TFPcUxD3MBueGJrKmeJ2ndjs5MixGIfCgz1mP8V4OtD3FYT3sG0WO3
b3n4BXDi7Ex491VHt7Va/lOXLBS+BHvA5/kQZWoAHJcqCxF6wfrit/+u2/K1vgPp5IaqB+ecO1EH
fZlot6LyrosJGZwDdeEOBy54veOhE/ZZ3+5Te+K3cdzr021jVwCnunsd/aSNfPTpDiIi1aCc4Wju
sQj9bBtxbS7UlPGhpAatXwhVt8yDhr7Y5wtQwa5XGQStHnXvH3I9Mr6oxrxN5ztqlYTdTx8x+XDV
EBUfJZALj98t3S653CGxQt9YQTrCZ7lqlwOROf9bNhx7vFocV5e1PfgDAPr1aH9FM8NjLbRAselP
A7XNlYySTQo02vRRKK190Qr5ZhtP2EJBQFXRIgmqPSDbG0Bt0RHBndWNmBOLbZl163mw+k7ANCO+
3hdF+nnIxrLwYSGTZ9+I6ih1397nu/Dpb+Sykmx5dPaBjewBgXmbfgvCVHufGncfSDP7ltkQ5lJT
FUSOHW/dM0nmHEvPr3hbW3C2J8+VUltMUQ0xrrZhfFfjb5VqE3qmn3aeoGispOWyDMFCXKhsVJh0
xG2XlROrmivKo7v/V9RSJQkjyihJZpFUGBduNX8WUPBnVHum+Q308buX6ZRbnUKm8x10tTnAN04j
L5nweMOCPmoFQPbDNldy9Rm65jhV9gBCHwdetSVCwYnXYRTH67eJse9XcOO/oO5HAcYh8Zwma2IX
jYKHfOa5qu1yT/J1mAcZHdIr75ig4u1ro0tROVOXW5Z6X9a8v1wIF38KEaUBLLU9V30awsm1Y9h9
Q8SbJLhzDwiX6misc8USK83gXz8dUP1A8w5SKhsvqF/fIBQIsAkjfTXfxT94wQ3AEU1xn6+EB9D5
rSkgRuqZ3vXnwK5/+5ZnH7zON4g+fIS/4O7tETiU2RAwdPRW5mHpzwyF6/UwtFljQDlIHa1ICvI0
WSwK16TJuzA/anQkjt6fC9B3WwvS88ixwehnH0MesmgexKkJPxn7t/KRqNa2B6SSZ+3WoERYT2jf
klwuyFK/FEcbzM8jV9dvWWJfgPi4DOMZQ4561RHemjwOD+VU0vEUru3w4rjc3SUjUr2Fdi8HYq8N
QeaZJGPhCaCpyDc2BM8lmTERzc6a+2YvHhvG8vchEix6UDKpjM/AUd8qVs8PwN6EWKKVOrXo4e2o
GTx6HVOmHasgQAjS16DlGdcjk+ea4mgE1+Gutj+h6ZZH5cNbCurOyhwirspCgu+SNUgsIgK2gWVg
kOiPeKcD8uNnBj1sGfI4nLFrVWKfw5z2oABPbV0hLWRVAp7MetcqJ6W8Kcn6raAXDUFtz3ZrSkyP
B/07R9IFMHBlFk5Wy7yVASnfO0pObit+1xSyVAzDFZqyvgwL9nqeiwk6QvpZU6ZJ8EPv2qd0NeGM
lhdwUkjoSWQKN1MnAzOnjNIaLuYUdc0db2rKhBBH7ISQiVYTgfuc3jZXHokomGqp+vJzssScJld9
ijofqclYdPJCtWQmRkol5907J0iPRnZvytAI7BAowPMCJRJg6i4nZCtYdTXpl8Nq9aW0hI3A4PSQ
Lqs5dl9/Ocwsi/T/QKCZIC4LmZuM0bhtz+W0TVtKUpJs8MjRU9LH2pd6LzzSMBgpzHiSLAdU6U0e
hp884ilbRb/ozxW/iJoKDS91inq98FQNaXw4zNy79+Vus5clSM55DRrN5qndw0VJoKlPC4hTrxM1
N1K/tpfilWuWNJx4+eL8dN85eZ0eEpSqJ43mwZahtSsKPTxT+ukp16z3lJTTL4lSebEm96tnS83Z
nfH4DLVshFkS3Ks3WhVpeC/UKUvhxNRN3Svp98X+ri/AxXntKDFAqUBXTXYjBCmES9Iz3dj95Tdi
pTjGvSpzPbnTsLFrHmHyTbdfy8Gzk3oww87WWH9s7PBnFtDZ46+XXM/v/o8aFvwg8uwjzfDQbO25
gfGd3l0JGp0AaQfOxXlvaUOYWO/0ckIFoo1pyZ6sKam0rRps+eUtVRZP0DQqmO1dDdkP4CCgxndp
r/5fhKJTewdvyemz/BJz2fV064xtIla8JfLMQ+FnQW2b2/ecMYH8qIDacCXOlS4ySv1NKS9P0Apl
jPZeaO4+lTek+jrEVXyShzLHyuGUZVmMia4fB4UcU5l+3R7e3xGW+cnEhjpsxJJkBQfotCBD/t4e
DPrviKoJ5fceUbNScISEUmEPGYdtKMYpsdP63yDrwr5lp8tyIYQ58Sh/uh5xxeUt6aCTg8rrY4j4
B9++ClwhhcnN7Z54JNhCYQYGB3xKeeJs4XIIAoBnRJoW9N75bbLnquTWMtH76nf0hoZ5bNGyrMh2
jB4ZCUjB1zr33hv0dRqoiCoPIyHsr5JIOhrDzGGzW1zI+rPO4Hwtjr9RXHK+Cie16u520MdoYFQl
sHhgrzloKN7GicJ4BJpvnYDP3MZwBw4MHe3Tz5cNjvCes+eNkLYRh9YsblksrmCX0CQk3QV1MWMA
ShoGqKYDo0uUu1d+rhtodJ5B4zL4U8m9CweAoAGX59hha/UnfodL5ox/Sus5QwGYBFi0E5C96jmH
xnBqosVJb0YbeUB3tASUvgJoyoogdGjAUW++bcb8Vj4LFdzq/cNQ7Zt4CkJI9ZAiikLBMAM8ckf5
e94VNyHpOLt78Axjj6GgTSmu4jL1G5zoA+ke8txNvLLV4wnb4yj/vyEemKYcEw7slVdVoQRoWqs3
2wytHamOGx1m2kxk5oAhFT47C1b7bXgHEjchhsTt19v1z0vyHIq6vyasx7KoIUaoFlCmBY5IhrTR
BH7K3rPSm2GguIdVJ2xz1SLREsu4HgpEaBiv2kNPj/609jDeN/OEBmu3WeK8hKgR6YzAdVpUeQdk
TcnmrrCgJi0iwS/45v7ihHkyB/K0DkDt7lBnazQFiSp6XjhXphKBncJzSjDrcghKaMD/wYGFTX0Z
3pGSNajeUuigkNLrzIwMXX88ux6i/F79SqMuctwyvnhWpmlmsICpJIAwPZl4s0hTLjAE72ZM+RES
4dku4axLbnlurzuLXp+qSd4DnzWUOuvEaQdNB4Cqzge9HlMimO3XO5cvmm9JAUHAYePaXPzYFFf1
IMk05E3EjbzQ8ZvlYtQX6yWkzR8c3MGByyyuCWFW61hIkNG6Gefbmd+jvftB43JEXNhLHrcUDIN3
Kj7jT1F2cDoVqr75Mst4FYULKx7Z2xOH+IVLLFXUJwgmktfNWeUN6texdB8EEG4/i9uhJHsuJt9M
0W4YxzuoZUQGjgoqm7DV207oB4U2ItmldFy17FEM/88IRkeZu3sy8GBN79ujpuBi/NxFni0a0oQ2
0STM9sMy5UhR/oy49Ty2+2/wm/ao3VAGw4Lfftz6QWbqb4zlt/bLqTz3CbXKa3x0AvRndACNH78v
fd/C17JxVg9+5dlRyH/fBPyeHix3JIz9eLDRaWF3ss+MG1Lc/lM1vprQKzviwuoBJZMArhn23moW
X6tSxoAJ7nLIy1jC572ejhX1BEr4OsAA4HzQ4gx37OwhKdjCRvx1/n0MVUhyM0V5P+zB9COzPhoO
OG5nsLJKA4rGfYVOEW7daY6i4lR+C6gZQdttPk4LDK5l3O6zf0r4TCisc/h9LRPyMuFKwZXQoqQu
q+V8a7E1gDvW4AZPL7L08GY21GHRMOxb5+NtSBl9OXzv3W+wYFo9/JOAdtQlhdjJe+uFv0VaEz2+
JuzP8pi3cI3txVZ2RKrXXz9PCuJzMS9INnqXUoCne6znl0DKHpQFsVxfY1jcMpX2zwJWeiavALXp
5uSwh8L4o3dSt8I2irI3Q0qlWKiE9vD5/fSG7Ddh2S5CZ1vixG0Ui4tsBnyaEc8pltpjzGCytye9
mEbrf87UsPlZzlo1cmcy7og40khuMOldaUp2okl8KATEXH0B6acz90fB6tNla3ihjofm5gpBZDhl
bSkFsY5ZDTHIwbEQA28gXX/Yk9DaztSYhmEmpivUPB94jMGURj4m/JsMCD6QkH7Bgs/ERFoUSY2/
KOzmS2zyXz2qpbu77bVNFT+Iq9WH2qVNJP6hnwLwT4TA3FFqkyAqUWrQlmeAopT9gAoDlEyfz5cg
Rr3Nizy/DDRYI0ALkFgRd+YviQWKvZksoe9tD/oJC20Vcb6tcLvLzyg4tpLkH1LEgRT3u1hFld8J
uRrnjS7p5LxdQugDOX//VXsa4Ff7jed4z8LLrVtV1TiWT+/fnPKxu/0wxLQtvkqJeLvc9/G+BOtc
WZ5POKw26Bn5re7DampbM/lzFzPREsq12JnuRMtIBcjvvs4R4aNAMQmPbXqDbCTExdfhTZtZ0chQ
ljsp3T9yY3URCSUq3zYNkVHtsMFYYVvDM/Mf6fao6uIq7e6E9eLu/XUDqu14QwblyqDS6dn4eMjX
9Kk+Q2+TKqb8yQ1aKS1Z9rEfd4owupoiEbjflHogUm0IB4Ck8yuiSLVn59BwycBDZ3v05JOA3MtK
FdW4O5szd8YrMkkykQ42YLuTVc8q3wN1L0rWUOgmKxR5dh8vCNVPbsZV1grtU/MvbyUwpOAln5D/
i/YJbiUL2I+VwPQ10oop0kBaHhE30ZA447BL+AimmoXnYMF8B9aS6NOYWy/qKkhZ+T948iC6J0jX
Gu88joIDprztRyPj41rvPAhAxHJ8d3D3C8rELj09GfxEJ5vdlmU9tNwMlB2ikp0jXK6v0KwKPpb0
P5/J4gfZO0rQyZfXE36rKRsyViun9jljeGX5APlPxziYDhQWpdc8mS6Ru1Wv6XEGg046ESqItPCN
4P+OMi+gVQk8SNUKPjSFqgOLMT6TgfiI97pamRg70o5Wveput6SVIJLG4ssX/cVKiofAXb8DQIf/
QREeXn43Em6X5ROtq76GVFud8z0aXKuo8dv5QlzezYrZ/H8nYKWm1GCpgR5wxL3+Dgo0+HL+1hvM
+0GcK2dveWNovhdNWrOuwRLRepG6shYxa6Uxnqp1hAfcmppOKfaMe0wXKjaCZ8ecO0N9JXdcBU/U
Srva+Qw7k4/kbhgjv6aAtf1cRXoqXD/6e71zQWsRChvhGYUIY3uI1cP1XvPD1KpnKKBlv+mYBuG/
8GMrsTH/SGvE3ZMZKGYuXHZ/qNxL2gSK7p+uF6SKio9SYYJHmfGG0RhCv4wIDZsd2BdWJbY6rYvy
hAWdo3I1h7TeUfLz4uFtQYzYzEoAf3u7tMxoUqt7t1MbR2pyibaGLoqfKapIKKVr8bslbxUy1WRY
MFPgQjUSY2pUxIyHzRk6uRgIiaUvCFkf2heo1+2BID3uUQwY+HMkGqo+j5LI6bA8OTqInwDo9XkI
FYW9av2SlXsXXd4SdEQsIsxI9XHiYc1lzy4dyOap+fLHMRZgazJhvYynFXQaZ4wEG63j9LFgx5yH
N285S01RktC0k1iSTV5s7eyTxh0wyvrfVnYr1Lqb8OcXxHj/UC1pYwyNHJFLtSoqy3COPKPATkvb
XqFAUlHk4FInyX7WUl+pJMfSk3vvoF4Q3jZpjPa17Luvcxl7G4sSOJ1rptn2rfMpFVStjSIuu/Mj
4k21QFJBza2JlhGWj3v3ucdl+uEUB6DttnBw43b3uXeB7IJ50i13gpOWXmARi+BZ6IAfHYXifpcA
Ui1aSWOkljt0vZPTMF5hLyFbSNDkb7FXVLQF/X6+T10GOA304L8z429n+MhrdHvjzo6tbQdWSgLH
t2s3INieR8/75lGs6VF+VsoG7GM0M/Y/+ywr6YxoXaDtjwOAEITCCu8EERy1BX2mFEeqv3aQxYzj
PbXUTej+ZSwy+/LqLMJclUv04I1hE4G6S9c/x1VP2sZu1h4SkqsAIaGHRitO3LhLTtoZrE5JPHsn
8ovAh4DLpTvK8VXN6LDZCkXZJ3AFxYPA0xyGf/QRip+EJjx4VpPnmSV5d/La3uB6xT63H4tgeRSK
ZCuLK3xlWFSRv7t5OsbN7qPsoPyZAAZ17deC8dGl2k1z9/R1ewzhiAS0pxpgd16YU64oKWHedLNx
rKs3Ffak2h0IdDfghPzXFrN8Z/UT/j4Jpdbgl83XFsowC/lghr+/HSNjUDqWGWZx82cy/whHiimW
LEetvnsTvcALV3RgHv0qkPkyRRFZRoXTcdW5SmBix/38ynHag0EgMEydSw35IA2PxTSLb1Mzznu/
HgH45x4JO0YjZqeiP59iDl899BKNC4BA1MxalZ3pw1DP7k698Nj+SBiLFk3JXUVv4fCAZ5K9l2rC
58uHcFfw5d+HKzRPKtjlJnJGD507JTJXWLH5Kut7LCIjpZPSxnZvkBTsjlaTg5MSMk8uRtMoI3xq
DIdTrOmWiL7A4bHKjkU91+km1EPZgLpAqT+yrP/TFN9ZTokMMJW2NynuPsBVQpzQT03q/QDm82Sp
43H9f8A/SSyfs6EuErs0iPVn2++zXN7uT5RdjZ08Jo+f7XpBLk2ajAZQSKwCglzLPeMoh0K98Clp
c1BHeJ1oAZJIsyoH5ZlfG6hpbl5y6aVXSb50Adjd5pJ8kukR/KOCoXYG/zHYamUyn8mEeK0VHtd0
JuEx+5b7ZJTxWPuMx+jBG664qgVUzXBpfhD6vHoWLhFl+y0nUkA2M3eGxLIHEX64j9AIr2XSWAKM
r0REFzzOVcgu8yDaYlF0cMN4cim+arzc2tPa/DESXd7LX3Lcr8VP/BhD9r24+iwxyn2ld0iDR5uR
0XPDxWphD060Pc9PMXhNwcXqwYEzG2la28YB8T3Zy/htem4rNS1N9M9s4e8+TSUh+VD+xx/quWGQ
FBc5erR5utmAtpT9JJ66i80BYrFk7XsPI6jGZSZzf0xnt7d4CAyyrAurPwHiN7ql9YGjhK9pFj2/
lovwKN5cQxNTlMvHsPiB5nxfSSkvZ4JmBPHC+nbqoG54UW8y3klXWlKCx+j5LZUjZebTXejaCmjI
SInbmNQyXw5gDTjWI/PkN+VN4sSV4+F2s2qV/avetTmBP5M7ELjm3Li7l2f3U/AGCMgnVIl7EbQn
837tQQW36ww24sMpPNRsWLaG16CwHL4SFfRROI51Iu1dtPZBh3yV+rXjByCdtw4KU7+kM/kY4zgW
6rtsLV1kjgIpVswNMvAqzXnQwclXAsLPNaijqOzfH09clrIh1o1WnfqEcWCiZRbvC87UaXs2FxDz
rAcPaja0u44uN+A5vm69VX/pPQ3YqCIc/O3tPAuetjJ8hyeXoF2bkcHe3De7L6a80HI3YkRl/CZt
4UZwQlydNVRZRWJeICgJ4zip0zVJIoKCDqEr/cIoP9nOWWeTCk1s4jnZrT/5dHBiKGWDcTkDy8m8
Z3gPZXKimpcvyQtUvWZbms0mubANfjcqKWAUUfugMxwyf9kG5OJNo1l1/2SxmUcTKjy4aPJPLEQH
Hn9w/VeLOu9cBQ3XUx1hHTkBr+CMEJ9FylReCf2H0KYFGJ5OZWcnoIwnfgxnuzV7SafThMmp969G
ekvy5GkcQ7AqAau6YccSBHV+weV8sXD8hic/9fMcIZQrAdUyrNyS0cKgkHV+awFYO5WgTY+iLoSB
+mhJVtrq67rJAMJXbqq2hj9GNGID1mk3O+Db2Z2BIK2cFQ23rJziQ6HnOalKWMQ3pwe+PhIlFrLG
1rZwMH/3dFYjtAFQ+Z6JD+MTjevCMDT3EUTTZkBXaAZOAShJdYrqIsgVDOOqtFo6/br7miLWTl7u
OY1omuwr2UBQ7+g3JbQ3GWPj98y3ZTxLjUk3iGzxsxG/ibcP7IzAzL3O5v3fnwCdV+0ka9H2IC1x
ZPb/6SAYac02Vgy4evCgJbgIBGcI2GNEDSbjuKYYryvZbkX5E4uzmcQ5Jf9Ts3rJS7ScbgAl/I9b
pVCxziPo2H3PIfksb2CICMviMMdPMwdcdNrc6vdNcapR0Cz9Dohajb5md28JyW8yEndnzd3E+BW5
6TklEqKKH2/vvba2fTCzUlZ2mvouHTioEOMJVelR2B891vgWqJvAOBmqocqordd0XKPMx+eMTFND
TPiHyWPDfItIjDLJp+YO/F2caN4oesFgF1GGvFmn5dMQ5ciQIvEqTex/8vS7VBGvc2qUBVMWNZ4G
b1nL+OUVQI9a8rk+7RUoL9NzDaA6tPk2jYnwOPuP2x+vH6bKpFo70zrHWyyz8NTs5fqAphnvt7+Y
/DcoatFWybXoy5nURYCStFRYA9by7evO188vy8tlDtdbBL4pn6Mjbrc6Xr5nXbN3/VtysxMHJ0mL
pXyYHPBXggzAaMQWOlmnOCZLkBKGdp6pIQ5d48hnXs0SQFyU+F/G2Vf82QBdyy7t3Ejx9HwoAIRo
iTPZNeBMGw9ocZ8MY4hra+dFG6nI+RnltThvh5Rx+6DTvTuUPPGuu/sVSyyaXuYUqND5DlORzMlv
cGEjuN4t8wzJeTrx1+nZxv21eOrJ3+0fC7tROJkvl/tUXXmoXG232AHgZ4AAgzonZlnMSQSswLYb
pfO69TsvrwcyjXKrjzJNPLJ5QDjUzgdp/Ilnl/6Dvm6rqldQ3fBaOljqhZKA855lL2hzZI0VfU/9
zwWkMxt/SQH87YyaQo9BdHauGv8ICpDXENPotlKtkTKHlIYrjgJ3mklJNL1DnsOtOuSF9aVl5dxd
qVveO272trKso6WYa3vNbtlXtP48FcUh+NRcWPvy8IyIxtd4uun7fg4dSY+NEDGsbq0JbqQvNZ17
2Wv5EL21e7W370/NbJwpO0u3tokx9nNJKKX/wX66QJJuj7rAzf8hYkamNXnUlG0n1D0gi4aVytoA
Tw6qt5S6diHd1szIzulmOcz5Cg/t/BwilQAKgMTrXBQgfkYj5Ee7maRsVJlosumhJBvPOapTfKmH
dcetjjQm7MjkjwicLFLIqEdvXRpKk45XO8c3iWiZJ2Fcljk65nh78XT+N3JrxReteW6Q3Vd1YKfg
KDgkImkTrc9EA/YrNS51oJrkJmBPzo0BUmec77epbg2DeVLUXlt0V6DBKUPV0vDOglHh+vA8OgzV
pu2ljllW7SAgw8c7vN9rC+vlDoRNGS14mRBKbydCJJBi+1Etp0OmvPzN1M+J+Bn8yq4yQrNmAlKK
qYBFTBJfdACalGmU9kjcyO7HrfXc9ukOTnOPto9pVfXm6GCTP8b2zvOtoVbZnh1DBzBBfXtiWk3y
SgQ23mbxIjB7WX65fS3VVeEg1HvquuV6kkP1xfbXGo8hw2gBv4X+lF1ISIH7wIfR9UmQLbxky5d6
ziWRU3L6VQuK5fTi6zccjEIPlaT8hU24zYCBPvr3E1ukIXxhm1C4cUW8uf9rwCva79HwlJsDvP4Y
o+6ueCMpYKm3KYG5p23XD4UmGafKUGtmsmK9WDxIPoycttBd1XPl2HFKosyvanb3gNaFlqLOPNBX
8x9YOnhpHCDaWcNPOwW+bP4yelzrfkQel+QjSu41VgPa6amgvtS2hjqog0fR8yTbFfcGF3Mm83D4
NzOnz0iBIoW8mNK7EBV8RVCvZl3gN95c57Cg1BVEPN+e5y8F79PdsXrTDofb4WaFceKpt/+/sr52
NAQkAAjz/9wdo8DVucW6fl/861DKK6ZwCoC2Nhu6UhA17kqVmybeuhCCxRJtQ42Zp/2a1ZcpeFa+
4tKVVFrWCVVspB0l/8uJld16T2WO/i8aHeNe9DOmju3BG4M7xOcIMViOMm5mHNr3VWoUELoLWQTT
TL5Ovr+MpRZwFyX15BEsBoKOuiRxR2BEi/4Qb1J/SolffZX/530nyGlTdulbAHpMl5flESL7Wdzr
z4xTA4nZORpjj8tG8/5vyOQ1Ma1jCO76gT88HltbIw+c34sZ6nmdGrBncrE2aL61s50eG/qI2Eof
xpLBv0qPNxl9zeGInIVF0e8+6Ca7SDMKUZ3wGLEZju71Bg/1/MQTs6m3K8plPsosiCQZ9Qb1tHT+
AMgj8owoP2dSeOAQDbHkdNoDyC6K5wpYMtKSuR2wM/1Bze1UNJxw1xEEK0YPGqLeeYIbm7CmcsNM
wRj2FxWg7t0lE9kGKCAdV2H7POwEXO6bjPXkMYlq6YOk0p3BQdrJ7RvDZu/bzNdoOIonwr+F4/kG
gvDeT5QouamnjvgcOlcsGjQa+Ub9HCmoh3TW5h9cqudt3Ty2GnS7ZCQqwDEMFICN83Qp05caUv5S
uTInMzq2scysgcnu6G4E+9w0GFKj8U8wCq3m6elhgdgOUA9bmugv7ICSJIH0tU3ZO8jpbXHLJO/f
iPppq7AshyWhYDRT6bjM+MERO8pawHCd0q0Yiy4l41Ls8C6MLHsNEl/nFSlDOKzcVLfvtyI0Shm1
YQR6gTxfxVImxebzG9Uk8BSWBVQsoHZ5MP9AGTz3tAwmOhH4/UQnQrYPTcVqPp0NDzFcmsE6/1Q1
Y+EDlUhVcJI0oItW6kdxNatqqjpgAxCIOJPyKom5MPkSwgFws6BYKwSw8xqZi47oBW3lcGk0qE16
BcEHM5VeO/MYYJwP/REiwHZXZUsV1aTy5YpdfhIrIidd2M6EWuvg8IiQn1MEAON5Flu7uoff1P61
ziW+GGKO4sOucLWKPbjCPSAez1B/61RPslaGgPNt0pmSXn7tyWAA9w7XZZmGwk6eGPJHqkgPJVCe
MMFIgZBJhoms/e1/iw3LPZDz6BtTrFS1ONS+VLQxorOqCslAJBI+umwbUNVJQBUQKCuoYuTgbzJD
tx13ULGADDJsBcfytiXuP/5xDzd/jda3H0FYgP1AlJLNK6YxIUMpU0rd4HAYptFXeeKGMSSHbKm/
D3x+QgGphTT9N00mk97MGxoHH3cTZns/tKiwqhZzXd4cGNhYAAbrmACcyXfZhtG41oBcMCV6Cb9M
hTHUCIfzq/GlaF75DR56XEHVwru/leOikNvEjxhctRG0PeNEUe1Gwrg3cfFQp4sg4Zbsj09yF0YE
H57FczW82KLLSdr8l5iiRjX62a6aztRSXMoZ2SCCCclwks/zPxleKqUdlDlGecT1S1UzzpHl/cQz
oVFWja6M+LsSulKSr3u/R+uwiqVzAjnNIeumPsCzXD5SVQZA1EXGnflwiaWupq9GMypYEfN4gOr+
y0OsG1abTUKQBTAtBqBOWp3RzOcqrCQhzA5zba85eQuLl9J3zutg8X1LHThNc2DS7wxfCPuHBFU2
tv3h3WQjTiWWLlu3WhMJJ6uFGUSJFaXgQ+FLt+d3O52rTQt7ukTGXY42deFVHAQts1+FqJIsolNJ
VtzOW57piWV+tNBRtQdqpImPDwVjaW2wO/ttlvWgiyNgAmQVBGrYH5x0kxlVVOSNrjgxcgSCrzUk
lZLFs5fRqL925YU3mw9dZL7NOZroY0XJQ5jK2qYWOpCJWbHjAy8o9/zvaz5gehOX3btxxKLcvsFD
wrveDzKlimlh95NIOMGdlTm7GqM5LTn0mMQPrT2AOfxkGpfIKHSYMjqjMZKu7HCy+B8dcTnf6LCk
mCISamJ71n0gshRd1tPZx6FPuTwqgBSMQi/H2cKkH48L1gQmbIh6fYRQaQiiiyvpmBtcRXYaP7Qn
VSoW0ztfs5Zhw03v3Jn7u71cpqhbUIAHz6Uhy9npjSCF5rc11WfC2NiuKd4I6puy/mioBJmYPS3D
FYgFwGHoZmOoj0ox5+qu4meRflqDzgvuuUy6bzQNytQWq0p87sSMvB26MGJ4se6ydoRHfQ0lVzdv
ITwRHNS8101swyLI/2T40F+QJMd6+dcWwJ+RXUufG2gkA11p09VM8EgPi5jBzI7Is1BZK3lGEB3c
CxUal1qrK8jtvhEyu9FcXDKJ3nOv9705sUz9T3RRDc7T83RmW+rt6xXkBmQWXIJDYjGAohXvKpgC
fY3fFA7HxsK2fFU21D63b8Ig+khBjfcUT6MCoPONvaZZVRziOsmV9IXTyYxtUo3et4//81epAT0S
wVUu2cErB4sB6gQ0A0V5EzWfHtxJFt/AammJ/ZbtOx6F2XA+zi/WHWgJ8c8WgGWy7UD7z9//hZq+
GuSydYdcNRy223ZRigjfTkMdeL5jgMaVtU0sZSMbYI2Db7ZegrmhN8vAQo9bhXCkz9dR4m03N/BJ
jWKgFX571mAQwIolffWeRdxWi7s7eToFPMXWdej5VwMoKO0dZjyi2k0vFbQzJeYE2GVh8DM9YyZs
ciG5XiY82Q41qvhLyuRmi/1AJumrINJIvbS3fKBtLwjLg1C+V5dq1ex7x/F8AE5RxbdBLo31gNPQ
w3WBWOGzIR0y4puuKaTy7ZJG/D0vtCs35IhM2mYCZsCMEJ+OQ60bglkhp2L3ysEgv9pA88hwUomk
He4PVCXsWHDngp+IaLjk9zN+YjkNYj6zY7RSJDxLGSLuNFOK35sg1slduLcf+e1eQUyBqINSXRtG
OA0/JWAQFZjvCYCY6XbP6S8tkXOQ0US1fIZbuoKiR+H91ZwMKS28JBT/Al+yJ2h9R7l17MTySly4
65ardmtjI4Qn3V2zPeO0P5B/AywbX3FHBhlzo1YRhB1H2Z9aOvnv9AH0+MYBX+GwppGOmDCnKVZe
yX4vukQO3qhGbZNDmwkfBQhGf+JKPvSc+NUaw2DfmYsWRl3aeeRw0Kbs71UyM97TWAH6a/mZWPCy
utEKPM/OQ+WAhyNTYvJkIxnYwNWuXAdNrIiLg0skpfe359bVPe+hdnrav1NKwrp7u6EmaySKWNVx
jEIp/AfxEpsiGdLFmFkh4jMG64d5pmkpcv9nddl4fAsudIEK6c5ENzfTZ1MLZZ3j9nDnUdFjfcdJ
CWZWtTLNk+TIm1z4toJq4RxwquDCIGENlj32DJyk0N/4VqA09XdBHQGqxMfe+fhw4cGg9XOv7dP8
RiipCmiDEA4hFPxGCAGYHK4CzpOP4rcNdNlO/HiRPqzTeQCWqPDjzfN/YhdgtH7LwN9UjCte/LVc
AKCVte+Uydht5Gb6Yva3N63GnxFhaVwy1mHq/FKL3y2hssUleOGMIvHX3v6SRFjG5sOinu7sUmdK
1nQqQIKu0SaWg2L3Z+gT6gHepk+JfmlkuQNAb6HerRgLDeAIg/9isEIFw0zzQhdmXdj1DCBBrpAT
xHvyEROCsa4wiGhAb4A3CMVLfx8edjznf/7slaKBDlNuivfQGE4vysJFdY0Xs1V/N3kpzfkbMl2p
61TxYuKKkcLul5tB3mNTP+MmeOe/FvK+3hr99yfRbd905ZzVhPCiosajri59zSZwh76zGMUwk8zy
17aMw1jXLJG10eW2fTg8LYGw7YsQF1WIC2WhiX8eEPx5DE3vmuPWNZjxiozvMsTH05K4aXEDjmg9
gG3tPV5/dI4hXO9tMjCz7Jql7M5nGuW4fFfAezHDNdT3n2WM4UElrkdUmBUznmFKC1T7+oB+74oB
ZjEmL96It287bRhxkSEXbZ/cDspk1QcNSI0nwwE6PsZ7Vaxy5wVXzMTWmDyuza2WjSQc1i7AEqwr
Z1ZK0xyfEOQDnOGiBXleo3aD4cyYxrc/6jqJ8NB8o3emT4C5JWKT6XEGbNk2TVZYIbq3Sn0eQ5ez
z83ngWe+nd+Zppmd1dkPXu5kmZvh0fGDoKYEwZwR+aVJhTO6PWmqKg4/U+WmjD53RwoO0eJzVlhG
Q8qwYm0qLgP5rQN5goHyOLFfDjSlxsoba4fZaaqipwf6aFwT+0kb1hotVG/r2JSfekdhFknYSsDk
gwaebrH1cDJ1tA3/aH7i55+ZyFnW+GmIeK51vBGhtRN8BkApIrEoqn771MHQFKEaIu2TRugEZ8Pk
lzr6KhQCroVlpNRvmeYPZv0wkba3kAEbNFEPW1cu9AIywHWqWBFK2rMDJ3mS0BuLcQpIGccCaizl
B+BY0Fqz92728e/JBHX9qpwSHLFIX9nPXm+FmAZsJU4h0XY30lycCr4bH0WpN4R5ccgzV5ZN3PBu
TbizIxFxOqUGbBBjhIHzMrnEeJBb7Axu0dRGS1p3aB3NgkvVxMHS8NFYrAK41SyZnG5kmwE1aAs5
UhnAWzo8XPp4ikSk/BPrkWlGhpPjoF3CvG7HnN1/w+18F00Xi1+Vn2fR3xGQBsPWD1zWE93WNImW
09p9QmGDf/naizGQhzru3MIW+kdotZd5G0K+axOpV5tbZv7lBEKXLj0B4P66IHEFuHXkZbpu6JVz
6tx/JapltmuUl3OX9pITYzhPLP/AXb6G+AgB4GbD5NyUCngJV2/SeKZvUvdAcSLW7KPHvZdR8U0N
DsvKmCAFalSNGXlP1orwULRGRjPQRyLzJ++aVi1EJ6jacJXygMVh2wwMHMhpmuZyEzJEqF1NoqkT
Zkka+tuta0WNbjzSDfyWop19YbEeKELTkjPBxc8/I5SBcq55T9sVcJwp7kKoDyTRR+RTd7yCvJfQ
0DbTsoOIwo92HD5mWPAYkf/wMz64vITmF3boJv4y5RT/2y5uPJS3kxCwXfz7cuEz+EFTZj8q6M4T
QiXRj6MqKXz/mIM6O0usUUUkCFea/D/l0M6cEr1nB8LY62jJU4jHtIkjzaf94UhDI9xI4BKslIv9
nbIgHweZMLvC0vJsgBLy2W4dcjO442nBGZIGju1PxQTsmTGQipN6H64tyh3l/PTOgAgiCJrSJVZg
VywIonUVQATxyRmZKnV8F/w1uopsc7r1txqQsZzRKmKWtjmW7+lli8s3PY/i9/RitJ42rvXKhTDK
uHAEQtcA+Mt/+Fw0jThDnu8KWta189JQH1Eo/X9y7Z5K0Xex+WwHSBEw70IakP28nIdP5qxitDFX
sDz7LfmRmvmBZcyJxF2DBU8AsfsAUFxRjhBOo79CopxS92J/S4M3FKsT+6KNxNINrTSqhn1IBwqD
2ju8iCRpiuxSjlQ96ygMmClsfrCrWyuDnoHWaJUdp2n1J83gdhJC6le8/w8PeNKJJRKH8X7dWO9Q
HSzgT4r5fXZxe8KP7SwDUmSdxb/eBbF4keVnMx3EkuCdH7l5edfcxCAPSVNZizxlz/GtLIfgk/o/
yOcxFTDwrMpEkg0FYlHZTNVJu2uCOCOH62Nu9zJerl9U4sfWjzfFR1e/WTF9ckPx+MZp2+ThqcaA
x4c3ew73bk7xRAoWtwYx7UAgLwvEOOCnlWshayU/LKdzNjdao+k6yqhWD5/g87y/CAjNijDHJZ8C
RtuQXRgcnFczCG9M2fiiyxbZ/lQwB1De0OC/zPkQAJb4kIalgyr6tcifv74ae4RZz3XR8NIyVrbn
e5KuUaEAhc02FcWJ8il5y7+YQW+62pDSknkrJe2LHwwJZhq0GCNns2+4fCR3AXPzjWKDzxfRGtZp
PK8HhJdeD+nxsL36w1VwHiE5QSNpWR+b9QJX8izBZW4p2aMwLVfaOvWHTa1W+Z77dV7lzh77xVSt
mUwR2fNAj+SYQPRgYEH7MxOOJ1UiQ5BXqL27EVXXyRplRMAXJDuF+aokTQ0wR5cNr1yzqPrfabrS
GauMIt20nU2iCwK+evvSzf4RdXlouXXCQJQkyKfXybVrG5QOr/Op4b2RAhMPl8sFbzGOzOW4wZwh
Cr1PD7+VtZdaorne1ppQYFU7PM5yW3Tsw9H8Z+/eeGm/jM6w8tuIVcdMHzF5mPJ9qhE2r8I56ZQ2
RrXe2dHXdcRAaY2AXsLgVBb8oxt6VRAQTkt27o5m7LJQjvrmOZ0j8WyOXrypAcZme/KHxm3oqXb9
ebiPLB79iXkEm/aUrEnHUAzNqsWcFKusySZmzMdMvKXUiR+kabJ0Pi80wTHT31aXEzanmCS/hM/t
cAHZpJrc9IlJ8O3Mjx2ZEIOWe4Q8xc6SmjngQELHXGbAFcgscIGmUyAyN6YO/WxGzKUouJc1wK6N
bdk2gvgqGRQhczRnGAne8JFsIyovcvURuujiVxQM/nKMzuKjHJRuyyZNnDHnL86e5XuiPUSNlJpS
2SFE6MNFjPLI6zL9yTVsa4DeSClropq8EWSaQY9atbMVrlOw/17ny0YRUTB/uMYvSSdTXQfPEhRo
QKjKDFjyUJj5hkWg1ykBS0BOfutnNBV+IiRwX8ORHtdm+rYtFsN1W9GP94yuZuoX1Q51l4WaCXZ7
lgo3bXzarVvk0LzcMTNszk/kZTHDPiNnk1y7p4xwuRlplf7X2uV6VTSwqTrI5y6N53/2dURGKV/R
P0STobGBd8yJan1Mj2tocdhRf03WIZsXLShDSsnxJNorp/GLPV5TwBBC60xdsxcEPhFquEmuGov/
MH/L8PrYZ2BCeBBKpWvqX/1pwYAGWhJNHwudrGkGu+G1if3i/HlJ0h7COwihZXkKoG6BTUApluzr
A9EWqPVa7QBLoKg90rZaOXPOD27ilw4nQ39tdBRcrsLyk/xPJH4ZjnGG/4syD5XwLtvQXaZKY1nZ
7YHZJ1ktQ6Yl2PKltrdu9Xp67CLfp9qCaIOjQ3Q4oorINV7DnMA9I5Gb9yDQxwi/MRM54TpAjtym
VIiYFptM5fcPRqyyVyC5nc4JtQFOyZJcqRAqAlOVhbyW5q9sGeEhLdN09Ff/zYW8qTQuIF03yHa+
xeicdYzyHYudpjRS48mH77MFyjpL9oDho6MwY7RP6aLUDarCbpeAx1Txnq3I1uSp9P7q+3hJAIwI
nvVuidgpgGAXuFiWte54M2ezj7quGhPmUqKScdGaCA74LhzeSNK+3QsZ1i8/mE/9prs7SubkrPWI
iQreE3MWtmnKB+b5Ioie5iPV6AwfTRV8VH7uY1LwGBgKIuaav9tuBgO19HXoGwvdb4XQIVNTjmAN
DCXpHksUgKBDYDvnQjwJHM2peMVCJPl8QCqEFyEm2CxYX4G2NMVsViHSk50xBN9LkRJ/H0t70l52
a03E5fGcqpTBCDdKIyfMEJdw6GMDMNkFRUTkqgbbjQ9s6+fTiArPZsZANVlTnyGAqgRqRj55qd4M
BCw+wNTsHtI+7bhkcA6xF2LaEUZCN/6tvLRIU4dYVf+kDeCEtqqqBmQIeVlTs9rsbelmieH6LU3v
Ri4wtzllN3NqQiv5NMTUXP9jnLr7UtT0lXkHw+ShapxL2hRzXzWv8vK4CQaOTwbvwpyEjvQEI67X
WHRctUv8Cah1YBRVnFjOjYJwNz1PYKNVCT5VzL6eimb+vwhBApNrMl0JbU5JATykFW2YuZ5vWABq
KmWvNemRbaWWKf/C4Zie52PhUaA5M27530nAG2M09awQnTmhUXC2XnYsAGQRzrO6VpRiJ7SbHux0
0aMpWimrCBK1uzWzx7XRzgaZM2CaTL3bIOKGH1WYB8ecEur0H4sFKraZeJHZrXgLvx7iWHz9RndM
48T6MAR6cTxNo3FWFKJ6AxJwQgy/jIQBEEl9oEHveMe3ijumZAIeQKHgDwn1aIYwoeWTYZgNdn8X
fzpZcYdODzFjiIgLoPkSTXiXy8J5Gm5FFqmA27cnCsxN25Zj7RS0hks9ev6vFh36Z1dabZAgSyj/
EaohK9m3nNIt6aOtD1QD0gKvXT/GKFrtmXYyrgEiIR3HmQ6fdjk2EsrlbF+7FAFOc/G0pfRGvz1J
Zwquj5xk5xNdwsQ9gLL0HIvBm+NY54U73cJRCKUUwmcb3a7NX9MN7P7NCZKxdbtbxTIVZVewc9GY
xMwVDiVPjrvlhi6WC71GKmMC2GNx4aNYjKBvzNk+C13THbmgqizJWIbn0MGFsz8X6BuzuF4XZGro
OPEq1ODtY6D/SpvQ3CjSRJ8MsUZ9RHc3GCPAIEyOVBsU+7Kes4Xl95ls6Y9WQ6CxaHnQNqFrQgzD
KEQ8gu+paEJZfCqT/f8sjkUTL6/7MRGKDBSVHo7mQRFekIIUGwg+xAsGgeLwTuwxKQnTOtYrIhOD
0qTmC6WgAgUZ2QUvHB8AHFTiNNB4CTLCGfxpirE49cHtFyl2oA/9Q/QQvMa3750VsMXAHL7oI2c1
uPukfN/Al5v/aSI4aAf262sIYKTSynOLsSKgVBriWwwz5oIxoXEthTRDlLKt9zAG7UiS107R4jQk
xVcnIplJEcTzmO/QIsFlq2AY+jKprHg0Rb6puAAcbNz4ibv1cKQh6g4xoUyKpg/Z+k3jTqBRdl9b
hJ43D8Ha8ZgaNZ1WqbKiV6eBXJ4X2/wrozqTSJ+MkVveFrqTcEDrVYjWif7WHevHOlp1p0V/vniF
eyvkvC25jU9NBm20p1YKQ1orucX4ZZ8PrF/VVKJxA2+7+fx7PWlio7DGG3GU/Z5iz43PtzlcIVR3
l9X9eUe3ih7Hn1PANoGkzDPRWzEJP1wGtpsluY74MaXvDNy5pcv+Cpzpm6ew+lQUG9TSchlSTIIf
ZAdLFuJXhn5emKSaapdyuNwTv42xWpU59JzOZ+VzFjqjobVs20wHdG2vMMPsQixE2z1aM2lQDAyg
q9rQQzbrYA4TzAQD7b1uU1sMqBbJeOIJJPAKBUvLrLCt0Ehc+IXKKMkVhpCr3uqSbiWWHX1lMrMh
0OheCP90vZiFGmNl45pXVr7hJcdQvuVl+14/euwgNM+3NvmwGRO4KUJY9MSOD+GZsvGBzTqQ5qXf
EuW/ZF9Pd537iFPQtklEUPOv0o0JX5a68WFv/cNGUWR5cBXgXxu8rtWLPsaGaQcQYO+65GQx3Z2t
uHnrWV49JY1usgdHK9YJ8DEyKRfK/a4/bp7YalAuYB4R59RRDhXSXYc6vWWXNG5dpFMysc/IN6a2
9uVUfEBf+Q8y+g0AfHXPj3Sjhu4Qr6D02sDxo1hX6MzXN+83/i0Ct81iTZN3R77q6aOV2t0tQcAI
P6SKFtArUWJdZptjfk07o6gK0sbBWpyDGeZ5m+0NQI5HCjGS4TnA4TK5r7k/af2e5PqKsE7lJz6Q
eo5Cg7nPg0+k92xQ0E28qOLvu41ctAi4kMxXhPA3tpsIcCuSQQOp4uB67p5tc89ofASm27Kj8L21
ALSHofy6x7qD1zsm7rETjh1z12s0Vpp0ErVa3GW1bDNkQzfC9WtRQ2gZY3oivs6dwhPkaD7ZqopL
I7rUWZ90hQtMze8ofJghYubQII7LCvw9aXxSS0xivB+e0LY+k1Zmx5Wq4DMtkUCJM5FuScGe6DXP
wqXf4hpPznSIY09W42zQVAuUje7fk2hSxguhvQjLXe+oxse9qNvnJktLJrPMf5rkGPUoF4a0iP3z
dlGirIhAAqNRyYoesiZD6V8c9kNdluTt7SLt3OSLLvAkfJ2qN1D3qTQfOzK17ZrRruV6sr2wfihy
fNBRm3kmoEpVgV9+TjYdUhziBGOz4Ra9qDdHErHBk/O0aPYKoqXxK0EDYVLkzqI87zuz8E6lU+RQ
xTMrTqatiiawAofRUZoa4E/aLfwQySKCVOgvxwbMQQtTM4DpqidcCdH9QW/nX2uSvbU/IjS9PSXJ
cLIpOZlR03jnKNq7uwNZCPf0YwA++80OMhD4bENWGmEYbuPVPwRgLv7x89HsXYyA1R+bLyr5AsPX
Q9QPFRUon+iypAOXrZOv5pq3c0DZ14M0J19ciMjyjuMla8LRtuak/+qHcT4sUmLxKy8pow7v/k9L
0aDrpHMubFHvZgS8CrDhqnLtmS0p1nxTjqUk1ybr6ecMZA/KdasNeTyYvftR6ku0TR6hMeVM2BnK
4kIP1jR7Eq7bq1cm5pMADVEde7urjvSr3oKU9ZIPogGNIHQNElGvc+SxRa3rEHuK0aONI5j7VZjE
SzGGz54ebkNftLN75e091jzIFB0Wbr8yGfcFm5tya0KtG9ZDUQEMfMyC/FTfX+yQI2Q4lUSjxpYQ
6HFxrkuhT1PHqVf9W18WUg9RyUHpu4t+1Nph20FoldH/mIsgNoAelqYSCHMl/dEssA0yrSX6hHH+
EcailjJ30qQBaGqi0TjR9RJim+/DIsRTjAX88K46wR5pNKiZUKauIAR73jz2ZSBclcFyMRM0VFT4
DG2VJrG9t8/2mMVnfMZbzFznSCWG+fXezgZdbJtBzvC/FTZCKCORW0H5OfzzAXU2D5Y6AX3nrv93
oD/5oVaAQATEzaXEgcwryIoOLSvkr+fdlPdPQ1/VxA2zOJExevtlq1wsO61kXvfW/SHR2atNwY8W
JBpEqV1TD2Yy0L3IjDatq/3L1YUjhoQpkfTwuoGZOL1uNdxyzNGUNVu+LF5+3CGnR8NR27L9h9NS
+EuTl9OVVCn8TMbQbncGuWjBNBOqnPptOkgsQLeFCZhAHc04Iv0Bb5Id/RCGuPpIqyGeFzJf+AbM
HJAfQbeo05ermpEYEJRQNuxaeqgaDNi5UilB8NmehGbnrTAWwoUR9UDBDlktVGngVsHrdNgQI8ZB
fJKOG5zDXvl7pXfEwO1Q71KTy/jLozu2PIwRnDn0NqGicKUgRmH+OIpr65EtXBi5mpKAWve74yfL
p1u/zig+K/vPUPx/1PbomvjqEMPWS9UBaSIyhXs58pLTidXecnB+24uO8YIBaKUKCZ9ufvw1HUXs
IJi4fyc5bNDID6nSSp6XKJ+IhEluVwD9GEZ59k/Ixmp9RXJKVgrZ9FiVZjQ9uuTy9giAupSNfjpr
MjFcKWD+eFI4FWifU1ySy3MyI9GfzJrWWRaNh9Zck/g83uYdGrQs5x+fhj4PUKbXnijDR0OaDat/
wopIqRofjhs/W34VktnilJcGRIQUioY7ZzWtqOpLv7eW+qd9ac0OIihrVGCKjGE9rn+UI1LFiKWM
wrpDSz8I6xQu/PyA6nIJJHBamfitr5LQswZoHQlUnRoE90sp0AZPxOal5WTiO3mIyFdIvKtyqsGd
xirF7OB5851Df/jpqTkfYPInQ7pUcCjwuHpMYy+Am+8ju14xivquEPvpgT4w2vwEQP8m0h3c/GS0
AJx3uCgDDK+sWEKF3Vjd+TmaL4BZqVOmmJeGWE4nv/D0oR/xcqp4ZNHp820UxT34Wgb8Flnu+1WD
2vQV752WoYvatWHBsbEZrFAuUDIni5tyk8tVsUWyhmzXkk7jNEjcXyjOC60ueudsX6r033hfGOk/
X99c7cfDxpz4k2E0knNNK46qVuhtMWYbt3KENRe/2wgWs6RK3yjiDcn5FYArcel4lquM6ocb90/3
ZbyirjJXWXaBXqfwLRh7tsShnk1cuX8fz5zjUufRjOPsu9Cv5ByiEnw0ye5CUrlIIBCK0fpgYhD5
W3DZ1TCt5XjPO2BCBCPVatEbLhaMYUQ8RLCh14ROssaloNCMaaMx9lJZ6f55RZG1u37s/i5JniEp
lInroKp5qxeBO1IMfkTervgubyUu8EEiDx9jqT9pjZoDAZxFMhuHSxFMmbkoVtzt9QfWAw4/Gkea
QfLwRvr+ntTxhcFQ4jJC2h7+8S6sytq95UqwqymxSbJfIP5/6EO5tu7IpyhRUdZ8zdimMMxtiuPf
uHbuqgvBAMyua+yXFAiORPiHvW8etC4FSR1X91IZz+vUbWxuHCJktP+b5GItFu5Vy0gijcPonhnw
Woc85yt8E5c/Nzuoyv5548rgkGsZ7OgPn4RLQCv4RT1ST4JgldXeAwSiWO1zYYer70gOa+lgDqgj
/WCQCffYIJcDt7FqO/df24owG6daftJl3XbYGJM1/bSkg37FDsY02XotiOddpQCQaTNGX6qCXiD0
tqoWL5Zlbyl7pjJ/jsSFuJQIohXcYIvBGeXJeup26Qdr6OM9A0tjpO1j4DIdAPb8ffM2Og2/6y0K
X+RqU4sMbCQfir+16HMhengz1m3okt5XFXFMU7b3lZvHO0H6w/09WbOzaF+5vrXx5F4Ndgn1YKGc
dIP5IlQmQ3+5fW5Z0208qXXV74/IYLChhjLadNxOlAlYK6YGPGsfqm5djip3gp6LCON9oeK/tATy
S96b3Qp8osCGCFp3WMSDA2fEax56ThdeL2ed7oTfVsdKNZcyRGmaHOvjureqAbDVrw10XKXpnKST
c/wsxbI1uCqeSVpGa8byj8u2ktXubJlCQw4rwAWyk9622XQU4mMa5IcpeVJ44mrKizvYmHicEORK
TKPKXMKeKD7QFREiG5O4JEchF2anOSR2MlS4DmERHpS/40Vh7VuGKOGD101x6S3djLK8wJ6esqHt
+WG8T79sRkvLj54/EEc0sUIGqwUFcN60Emt+MO9sHztLp84TJJkfUG7J3U/Qi8ipoNimAMYnM5w2
DDxA0zwwDxuQIXEie3f0lUWH59kIiNQTPMVqDGOnEg0CmjHiNnf9jt1ih8E0ANcodLlJOBr8XuM4
ldRiYt6vbqUy9BdRuP61l9/zqEr8kZyiLoFmbwB4dN0m9oK0qVOn6Si1PqFKdHTml2Zz+VKG/F2w
AtzrrvRoPTyNuMBxUmuMiiMaHMUe6uaO9Us4FGlhoEzmvv7iVt+X0QHaAV9oczlDUC01REZwbCfR
Z/DPaQ8gYEvV+UuEVZTL3GWq2isCYV8PtFjSCjVR0I9AsAOjFPbgbLSskkZEp70L4nKD/Ip5wu3e
VswyjC/rFsKdpCoWE6WjhO+765Sxc9L+peMX4KvGdkwxK1gK4gmuZ03Z0RtAapHL1VvSngESEQKs
2xwjF3XrxjRJgp77jf+o6y1nvu9fcHXvF9d4iKqVSrvudM4UdRjEGank/BcIgqj5quRkSkqByIxh
uv5LMaAZUobs4RjXgqnAI9FSn86nN5/n37b/5HgjElJc8uqKOjpRaXwQM1WtWoqHmSemkk6LYhRe
OtQhMqMu8gmwxOoJ+/A7kbOx2ZJB2HsIo2Yz46oZvpApfxXEhI+eS+9WLk2N+2wcZeNE9mdYi/vn
7des10zYqZPkUYo8MfO9NKuNxdMjaLWY2q2FmyzdBC4xtddqkp8/RpGyeHQedp6r2TqQWTvreWi6
vs+t3hZmWiB58/JJn9s0T2quD1HANrji5aTJ+yqOGBFqZkrrHKYex1MsQRbNSGt6kbFBkG6OBEr6
YcNG5clc9PzirRz4JDrBng+ZXF13/+EzdDziqsZyfXgDhjysDs3GCjG+MzFVtwh8yoKclef3EBT9
phzFF8vP7EPYfGN4nGm3DCrPpicN1T2LXNaM/YILPLTcWidZwdAjr6f33Ipq5rr5rJtmwMljom3g
xjxB9zim+oK3fZnLJs1APZaMVkrnjSAcKH7/h+FoWpO8g+e56zGBWJofrCrOSxElklZ0JnLZkgcw
OrN9fVWVupDdc1H0W5qydNvM4p2uBh1FjicK/IjFEMeip9QGgcY+LW5nYRv4cbOy49XpT++Ftcj5
1g3zZ2OUShgxpb8W+Xm2b12M14dhFnhH+MI5VfUE6wso9RbNLThS2vBbs/sVhmcG4o50TB1Yiv+H
qRV2oclTgwAaNu9hCBLB71HuUuty90dIqpXo+j+mI1gNTGe1K01Gr8lEiiH9fu792h4h++FhWzAf
0KT3gmmOze0pM/fFyFSc6Fj3wiq0aYHxYM6UcJTe0um0Gd/6X7JCbADA8QQg9RJqZey9ZcE1HTmg
0SK+tQUkIFaSGC9dGQPfq4ThN6XktRDKVFvBRC2gpMARI2soVEfqc2dGdiack9Oywi0zlqv2GTuG
MKIIm4Z0RJNbQvbN8b1orjHhYcuOVx55rWXq2apb9YneV60ho9CkhTmelDT7t0lMGhQJiAkHjm0u
/IKTtFqeAr03eFs6G5WdCMPnBavbz7axXvdql3cJrSZRye1qkG6VxeguaJmrrEe3F3FVzatTS3Gh
PMnSsJVuZ+JeDaWWF0AmT0mU9t+Qe1HzDVbyTddtlYZBvL4/vs2Zjo4HYac36XQwwy6Pnx+3dxOq
zh7cX8mmR4xb/WrWMA5rggxSH+gzNxHCHJtZQ1uzW1haHaD+SPZFhKfKe7judtN6wRadADQArvW+
QGKAQZlfAbgpI6YkVyqxxOwt+hw6RS/KgwwvFooarPAYmawulbNqAZLotu6bclSyJE/eRYwQMioi
Btnu8CWf1Lo84ld0YWIhlAqQVDr9qCmnXbeJ9Pv8hNJuoBn97esRrx3rVQyUoFxGsDE/5IGQ4WWL
dp6bnsjCf9PIRstWatYAelDSiskXxk+zqMil+410xkEu4P4oDpi/LDvxHY6xKwsIYpXB1NPBk2UQ
4k6MSc7bk4uhSzIXzucE3TXmcGKVzorfqaGEDKH2h4fTjTehbS3tZsBx6iH97jqibR0e6PvOYIuQ
FJu33aTEifOTDpx89DBfhoQKX3/WRTbPMdNbGSSP7H7wxu+mTMGLpp8BzgfR5dl98aSOmpk6o3Xo
a/9nkdT2h9TJFa/OKAi4fdQ+I91OCln0Q+L5VH3m0xd2C7gI4uQTgmRrcq736bCa+lTQG1UmgAlu
Et4+fxJT6D/QEwD9BSK50v9Ug20Q5KjyN9nbkvJqvkkce6RZlD+LwsmqXxwcBUAtPc59BD90RkGt
9ScTIbtyrFbwnwaFYxAa6sAaNAsb6LWcz/iGNqBg5umVehCOvgbk1vGrkvFXTkAoFoYFoxJvxV3w
U/+VCewFpwLyfCFwCd+eVbklb/++ymbKKJJQTQBXXjTvd9knyHnGzXSpa2tFiPlscNeZO/N/kI7R
JweU6Jvuh2nT3x2jCVPr1v1MlwSNJ4sWUSllza35Qtx2HoxIrYqgbT+1jthAbz0ie0zKgEr7zCxw
waTPQ9Y8znocoKtAij5bepp4VAqQA/zCHzWdY6KqL0cF0J9oaGIKRttKvD0HzUPnd91gwzn8Bv0r
hgEBfmtKXnh2ROK7TPFVcWtPHyJ6TDPdqpCBrgDWZ98KMGUhDqlRQqW+/5hqzPAT1Qqw6ObvVc6/
b9yCRPVfD9oJ5ADEetAwMyZ4uSvvZYEqbI2WDZ4OKAG/nHSN8U80sZJpe3Ae3scTOLfVMX5rfCRt
n1hMBHHgK9QJkIPD96CKoEycgRUw5D3aZgPLhsxdizuTWfs+IqgHGItRsBjXLJrTzZaoh/iMTLWY
XFxHHDhnkPVYLZbDpY9/mWXj2YX0TG10eHc9wcF1b1gee4pX2Jd3C28bZkJQvzK/zSFOmc1m6F7l
djgSr5eBdMl9ZaoFmDtVxDbF3adSDRir1FyMTrPeL13biHp5nDwRosjCeLwhOE164WfY02AGoHTn
f1MqKcFMQwc3n+NpmxbasKhtpCxhWdTc361GOwuxMjS+K/6fDbdlJ6Lcj7E9U+3LDweOn2JJMqc+
S1TCnIl9/nvjMRK1M1H9XtTBzZRfrgJPbKC0OLDnq5L4UawH2hDjGtxC9OEgomQYZ3S8w3YudO2b
+IbXUDxINptIN2j5k4I2Nsschj4HeS/EH39nC5DRtFi+DMDTbXmxDdEtjsGVYRR6ApTEuF3z16t1
Kt+IriP4JSiNX1BQjT2gTqTgY2g6vBlsBbxUitGaZG1ynpshGjleaGEgYLUD2LkHTYCL7VWkvlne
mdALVGWUL4QdNtVHwiUUHeFdSMXv6/5rAhAAU/VP1+geFMpTfSWAkS1Iisk+fNLAprdElN/KQc7L
VVY2sIEZzYOcyqVzddTPHF3yd3n16J5CFam7BoWfEMrISl2TU8qgsCsqPAmG/i1YRmLMFZDHk/hx
Sb2gtlyFeIl9GYfFfCfhuOTaAdorFfnelI0jGo3U+TQ8Ipe9PlAhVpwWiGhJ9igbt1iVUokj4K5C
Y0fV6kY16pyouFGmNOPNgwFQ0Wds3EBPS1j4j7q1ptLsPbtpkr7H0Ungz9XU7zvR0Ey3cPjcby4/
IPDHYz0jOlt67JPfIbBgRLp3Bs94RjY7UKlWiw42Mb/p4NP5nVQY0pHuRa5gapEmW69pbC+IT8eN
GzIJkRmzbI297zh1qeTCPPmXlytFcVEmwWoRUUD9LfsxTI0HwpZuVPXd3Nvgetkr9oaOqX+BsyC0
P0874njp8RRUKgknQKX94X2CVFgaAd4ygNbUH0MRg6w9k1sI+MG2ivbPhSpO6vKdIRfiZH6bYX8S
fcvPjM8dgRfGq+/QIQii+ofsgaIfxIu7u7vfOeVAlK2/HHGMDrUegqPAaqS10iBD8OcMXH/03Dr1
IjqtKglWHdiZO5t0i+aR8KN/vN3ArmfsBDb9LZRp3Vuq/LxPb5M0Xq8xbUr5ynqpkh1tkevaOQz7
50Y9rsUG4r9n8dZ4j99DDz0WmfRh5IJYfaVdSHR3S9fYu9it69fRYiqgql87DeZ28Edkp0owDASe
rl1fnxSWyCMBveLnIStcRC1Js5aTSpCqK9Xn30EIhOsPO3GVlaPzT4Kc1BS+8+ppXBh8Ccb3ASCi
5+JWWtAdFCDsv30UNDmzCWOkWNJstLVbwEZxml2ZQizxqkbl7RtXLsgr+ubSdLd9WZZ9d9w3kdMx
5KhHVcQES5LubCYHjYqHnjUUbyqw2lJ//C+/2QO0NUruAvop6bh5pyogySoD6tmYNuuqJx7x7aNx
GDrF5cK3ZQtDTIqs7NYkMkhPK64S2mjZo5pjGTTD/Ahcle/3rqMenMCkz718bbtZOvI3atFt6g2N
CCPE3esGetuljaWw9Oz0jsDS9WVkmYqUptPiOjlhs3KUaWm1CkQyALmftSKd8eu+0zyvFxMP10bT
y97B/KoKCuUO747UHREp2vT0I9bmg5E7UZocFkv8SW5ICkp1D3gkyquXmxJtAbg1P6m4IRsMmv/a
NpiK3LrXxHOqAO7OJkCIh+H/uRxKbOQLlp5Vzb2xw+QeJ/ouvReUdkA1TcFbUjiZTX/OtLnucCh1
imtkXKT15M5wiAMID5MZFtT9TU8ltGh+GqEPCtWto5gUJ86ALoSJLiBpf0kNvhqmFBG+3/yra8uQ
aVq+UGvD940dx4A2mtxmFtODU67QBISj2dg1FikjJOn45sELxElmqapd6YcHRlbMT55IHjqsPwWW
eZKjdvbNlXOV1rKtaCRXlLjbbj57QIHHYo59ThUraOjheadsrHAyWcI/1dM7AFglMoOobDww/V6t
4SUh5vzboYg3WlxyccUI9h/gTdXTZ6/8Hut5eZQFlENEok7ZRfeDZAGEspvUH+keymBZ8z2PMsJE
yCSw2zKWSdZrQogrzf6pvUcK+wZUEIK2pG9I5Nh8XdYlbGzL/oDTJbbiytGWYFZybJqu391qWi4d
Wm8SJybUTWMyQQAYY5A0JCDLTGwu/O5o1il4CIm6TX/GB7wzWspage18Fjw4AskOlq9D+tC/0Qg5
j+VNCkvsJIGzWr44okWaTdlNpZJwftOxiUjAvKivkW7RE+TV/cojCmxqolgCEZi9ErOWJ6/RRTfV
Y9B7aqyi8HJI0zmmT/SsGOnUM+W2XqHo2t2NDANfVE6QygBkKtEIXBwXpQK5uGLDg+GO8lG7TbOY
khQWWo15ikguEjOt8XEyzuwmlqCJP9EqROJsVvINSpLbA1XqZMu0VpJTssWQlOYc+TrwEgD3Ycxk
qdDD3Uh6/gaMP5eh7LHTV7qmw5LcY9ysT9y5nyKghGF2OjU12Zhfh91gb9K1OWz375do1wEsk9gT
8NTdDuom0hIe1mGUOL6rNWdS1qR8Hz0uezmCxtnayAQoRJHg2J78XbdEmNGBnYZUBhBNn9/fLD3G
ngSd42mIAbujU0tZG7178izbR2k/WaQnMUAUtNtA4Yp7IUdzCeKfsBsDTMp/rphrdhU4rErPNnk5
yjWopezZ0gytLFn98tOVyqUVGscZ4KvToKTu9c3bU5RcDUsr9Ht+EVeA//EIHUkCLr24VtUACvzx
1o5jPOkThQaD10A8xflS9RMO3jUSqDWev/LyH/ujey10+XH9ryuzQNHiByG9VIcomjRcveSfKWEM
YQqW+x9T4mMIdo0MwSrh/0EaQ0FXgA5rTirBfeVOAr1Q/2KFP0jgUq3G/mWNC4ZmkZSRkvH+YPIT
goc5HCeyolzgfO2TKo+TQnfggKoATePo4wjE4Fon0jPoAKi29Bs/BTXnyT5YCAgkrewpUPp2RrI3
2XZ7qAiMnLodUEipm3cpywYPL/lLPJi4xurRY5cyT5jgKica+zYwe/xoOiNEzAPcsHxN1wysjsbk
3LTU0P8IM2igOsVYUpn9WO2DeiPO0DG8xp6JnpI/AAjp5ZhIykCBW2ClsS+w4wz01GReWzlmIoBY
jiVQSnSjHFjhXeiWixNgc2k0/nm/n4eVI0Z1hIiGVgcY9zQk24CTTjWKObJ0yG79CKOavKhGwk6N
D5we+yJ62elgfpCCFwOQ+YSaaqtDHyUBJMEN4IwFAtt2lcHM3IxmP/IpecpwDWdf4VbIMds5/PF5
FSlv17hLY3w09ibPbl+HawQ/X8jnPouQIxAIn3i1DTuXTwIXX10jxrQZekGfs97w6V/kX0CnqvqI
Qm2E3xLMZcPaF4LmmQUaIP6N0qAej1hOA4JySjN88gncrIlMKx5rpyt1Fq+TKDStT77lHsco+EJz
V+kyRTSX+jHhDnWY3mZ5jJk+pgvcujAPpDcptD/urK9FQXKl7tsL7Cv6j4U5HsLPxSbpqTothgpq
SOQ7QUvbWV5InyQpbCkrzpMswGPkuKpL/tRU9ZcRzWzWg41j2oR6e86hH9Rvkv2IqXMMJ8mFcfaK
rThO8Gy41L0lyJJc5Da6FigQyxNU1UXIoQSDrREndnOLZGjz6YfSDaQzKfmI/ReO2+ILULO7PIXA
8mGeD/UMl9qwEt92SjWzdw41QZJoRKTI0KZ+gNwyFJ9HZXwyrV7YOg1jCR7pNrUz0Om6eRGgwtTy
SVaWgjMSEMwN0e6OsXytWPVIubrWthnLBiavr3tFopIXT7DXuCeZ0raxC01dgu3wWJSoJ6aVEjvP
6MXDJaseIzOOvu8Cu0f3m2dbTyNHZ4vZzObgxyg3b+EMqR4ROz8svWN4rhLObOuu4nlndy4bPo8Y
+K+YMBewHUuwoM66nCzYPt7Gc19gJ6CzC5JPELbNRtQxcanKIH8VB9ZC1LRntynYXla8GSejeAQR
kG51duIdAjuSGjj2xOmrdNPAe6nN4K7seTfNHOun/kx04dny1yB1E6ENXqJfe9bUPtnhXY3yeCs+
xp7hx7ZFa8vnoDud+wM0ZKZ4UBdjWRSO1hyMM56iEWlwii07kqmzo1GkJ8PEk/KfVx//UqXxWQCy
hDACHaVAXTNVQoIqzo0OPleiTe5nLEN+ipz2Su3mscwWM5zbDRtH5Fp0ejME2quwvuX629uJkSWX
Ep4hoL1A+mtxCxme7iSKLa4v/9Ypv5TRoKb1Sn7/ZNT6BOmTWf/uQXtO5y7TgCpv4jx71tKWEgnM
jpdzx/1Xdgm5MF4823Q3/czCArZN3A0tsowuI6L41InR+mc+iO0mOpoUpl7Fkbx3UqvTMWM4YlJf
w7Rv0K0eBaonl/00tYn9a3b5t3X174is/kqlkw6YTf49/GD40VFjFbaQstbYLWY5KFD6hol7lPjM
ube4dMLd5J0SH+xe/rYSlLAkSMU21GsNwW95mo1nCS+aYiVIq7M0U7Ojg43EeQpKJD7aNyqhb5Od
DySyOYXUsM/k1j+Gu4GG4Il4JX0wNPiXorL5mRvuB9Kzn6vXkgX/jEbRnDeL9UfIYhf1lG62H2rB
Ldx4pUFu6qFJHAT23h79lmsBzoDsRujTtMu6Z6IQ/NKuWZwO0+lpg2ujg6QZCMQBX9hfdMvZtaiC
zu5nUZ2Zyz254/MCUdwVnPpTvejJWfdIOg8mNdRTNdWoFVcBupnh5/ElBrEIxqDhvaH8JVv4l/Nt
S6nU74AiTHNuJR/7yjYmPnx90YiZPsKOtMr2Al4lq/B3ew7H4WpdZPXXhI63xt7rgMheDYApa+Nx
+F4/F85Dn9PwoUlo6SmeTVlqZn/Zzky/G9Q/RFedzEDz+J3BbaNRGjiOzmqHEvc3vC7kSi+tjCyO
FWi39uvr3h4jTO1NLnoi7XuCd/LYW2lqg9/baPoymL/XEIJOP5ejHN/w5DGgj8o5cXTB9S2ed9sV
VZOd3dxuSzziwO+DlFuygzC+x4ZhsskAoIU03S6HayV52PcaQge7yx12ocP265zZRnM1Dwmgatho
Cpzrisu3dYGURHscNhHaQWF75o65h/KD5ckCbGY8nfI0iTpW4n2//ErZ9bSTsOtn82CICZ5ZwyFg
6gqFCBgMqoQiY10sXwqFbswZtcI5jrP1rHoRrXL6S9dDZzSuye0mvL/FHoUssF71nVt5CHDAOYMx
kp5r7xGIrdyQB2ig6fRxlv3lfpXqcL8zvSPl7FgiiNkRHG9gRQwNpK/kfeDsoCcFLp4oQGab6vDc
H7x1gqT0S1s4x+36kuU9ykc4iCGDPjE5DZvxJ2Qd4ICljlHxH5DMQzjEH2/DdsKMLUrjlcpi5obf
Cpn2jzMrYii0t8GGrgd4hshhsgFDfTaJI3sXudg/VqjS9MbjVJrNFDIKdomnJMdrHWA1fw2Ewz5J
9cdYpzjp363HD7k0O7I48lc2tmRP6GJ2ZaofenGQWEB4Uv+oyZ4QdTso2omhPvVrHvFOFEn+gDhP
tGoPZEgINZVfIEv3SKCSyU1rT7zco0LbxlB7zBUI+3ZF2gUOi2+e2oegGjLKYU4iM7z2t/cdYqG2
4pi0+9pUPJd7lee3vr5a/goPgtKIUWXKEUVNSCkzydLj+SwzQNQ4zlrwfx5f5UYxooeG86fBWgvj
DE4kkR8TKglYXsO3/G3yj/TO4kQqHXRZLDXWKlwI586I1kbPkubzX0KGEONLO6xF2HOD7j32zCEn
q6u/s/CwLHYvfvJ7dXAUbJV1yjaLpKD0n685isL/vAmNhR2Cn3OjtGqFN7jE+eisTch1JB05GtFO
Cc/VWU03VBL5SNywyxuv6BsAvgSJFGRjxPA3DanmohJ2wOPAvX269HiYJzFGEacMcoY8C9G3kYgq
XzKNr5lqzkL2v7qOYpJ/Ctqo7Di5ch/Q8BgLDWEM3Wsa/WTNvwsjxX0j8Mc58mrn2SyNUQyCgeRb
yk1Ty24SKx0Wt00FxRiOMbXi1BzehOLnSFHpTPOgxB2xGXsWMG6Nhk6hbdX9676nb1cChxIhZMH+
RGnQ86tAfsN24/n3SoUhr12Aty6NEKonpEtbyjm8nUzjkDqQA4iAi6GXDlqfBQlEeKFcLZxEJ3b2
NtPwDTRmPcw6legAGAJik8neJjeXsiHWC1chlD/AlK2i9p30jJTgVOqkn4dGUbftL6osrA7ondzx
/dZv5V706TMI41TNnHTOHq3mF6jme/oAM67RYPZjnsZMUieHihjufXhb4Zw3IpPBbEL6aRZ+ipHf
jF6lsDpj60oW5e3MD8AxFW30LMPNcov7dLs7WKBsMdlTl6B/WdTSE6cJn4GoTp9+TLBldtRJ/qM5
dWUkaZvmQlBIm8+en2yRrr1kxgFRPtQjfkQKS4IsnblcYD0Yd+GPZJ8neYsIKH1tRpOUOYy5rklB
aU4j1K8EIQAuoLHtoRhHEntR2kQ8C85KAMPa+KZ27EQ9WZDJ4VRzV0S4dwUNcJihdCKa4aSwFmpr
STBHpyfDgDTDxSejUVw/8+sRbSnN6MpXPdjjFJmybrwgwAq0kavdpr+hHvEEvRytPEsuNQIImiTi
292md/9G5gi+lAQ1dQBg4mWvhKEMXXUoUNhXum7eCDUalfUHxtgVhGIAHHPdrE3MptNmnZO7lKYK
m4YlVfhD6CKT2wrTASzZyV0VyOlc4n7UznfCRmv81sYJefpQ9W7zIplloc9loIUgK5CiSxVtZ6oi
puEyjrVeOEXWkXAlJG/6m8GfBmbeL7lRfqzYIqY/Ko86S+KH+TintF/IqSbBhUuPg/snpBhNLj5i
lbKYQkgihWIm/lDu/mVN11oCFchOZMqjt6F0WCCcR0lXWuWC2S2x23xNsMDe63El2GGSfpwEpbeH
zBwYKy84XlCn+YaDbhCKzea54igCwuqEP0a85E2WC0ya9Riitq+BBgs6JMzJUKbLn5cGnyfAWxsC
XRHLayxUWvsx1umR3sV9yt1Dd44xW88jKICQR9B0OeMrRYy+QPcuyNLBPxK0HwFtRc59OZNHI4QJ
2uZRxOSXitaa+au7G0vGT8Ir6am5T/w500MoOcwGp88+2LiLH0R8b6PohMOQ+jhUTDpDKn9Ligtt
CAfWNRBLughpbg08bQ8ct1t02cXuTM3F9zd/6JLNP0aC/KKTp5Vi9YKgV/F6mqp4mGeUhCgqqw8V
L/UkqK1uGg+tV7z+0L/+J0G3sJqk6xpw0IE/fey1vKkjv4+gINnLXN0tFzY2KOHzIhtXhuZLdj4J
mjct3ixMmaAMoNPLS0SfYNjEq6HSGrVn+l2WHqikF3ZVY2FK2npyU+iqW60yGPlSHgKQOnA0RDyy
MN7C0UPBDZWNgpfcnzmHXiLv4qrWLm0QcCjalKYPhmzIWPHKw3NlZuJPXj2gSSR7HL6jkxE71PbG
yX+LBlcNXk6w75QO0VTlldTbbnTbyEB1L1HFWARn9qpP9xadcJQJL4PyZa/wE9agYqeG9l+bgr9J
7eCxnhgkBNTB4Zb7hU0YmayFm103RYU1cDQMYRASBIAUUDuUWWujj7pnFLH8IRcgDd36cfQY6sF1
hB9T3oNSkNtYjrGGQsmMdJ6qkkBuYfSwYND3wORF7eh9Vgr0TVcHoZgmCKZ+rNzlTZorOOGh6q9D
QUIkawQ+fPqYR+RsOWaJwamHI7LJvkH0ImeTGGd95AlGFrzjXnSA3tzeeIfTUf80lIv3VpQZ6bVD
RdEt7y/udh58fHtQiIaewG/L/N5s7LtdyLIe/tvCLdywsjEoKlBTKZba24VIzSPl7f9HUYf7FHzT
rgJyN0EVD+VFDOVb+5MYu53lVmSAOOHvyOSGNdD7eLLfEn5mfwdID/gaKkOpSIvPlVZ+ksbMZTSr
LHZg8dPTC9zXpqe916ekWQx2+3QG6dFqrly7/gunXkudayoAEQYJOsiSVcbd2h2GRG+s9A+FNHH7
Odq0mXyI7v78PfP2Ho+owMqseQK1Kd4KYWqnzkoQjpflDNEBk5zEAlIQXZyTn7kf6PzcDhOPjCyu
tDh1tEtPGD0YOg9ouijttYMoPXwh6dziJOGaukCKzxirXVuWBxQJvQfApRXUZiZ/4zMVI6APZwng
yX2RsbtYAfOPzZ+hvy7aJ/uI0GozIZ9EPRAJMrl6yBZ3eeMu5NuVYRUAJq2RE6Fl0H2V0L8JJ0SP
okTVdLWNljbpKTY0TeCFYB0Nif3zAAPa3EziB4hwwVQ4LwuqYCA3Jr3aN4YXYV1w6nlH6t+V5dxH
UjykcPyGehsrkVeSk4yxH6mEYSczHlvgfqheFHAyfoboVPRtkvR1FDMM3JuEq1XwvtjJxVWBr1CY
3LAEuLm3RXYAg6ouXY7PggWS0Yjdg4skXf/704pJB7JhnfJPX2YTHS0yolJXvhZG4d8u3XfXyIsv
Uqy4l2BU5GCUqGQNIMKCOxmziaC/VLe6z+b6ae69KVM/g7UQLkzVFIijYU2dCMXBtsDW/CxchVgQ
Nr/iSWYHMkoIJ7QbORLLA5eOdNyZTzExjOrWa79U80rMy8azyB76GBkIuaPdhSLLrrBCP4QaD0C4
486JtrSHG4dZG+ElEWn7Q3VX6POx+MXoSQWv6R1mImr9NE/2YXwIJZI2asS4/UN++FYKPifxzVEY
F7Cip/lUPNqAfTOBOrKGJ4f9yW4NVI7p0okSjc0JSs4wlgk0AHkgKMIUL0vIIniqiDEEuMTRxEEL
ErO6YMjyP9F0nlDJXjjA6dDVYhwvyv/xQgjjY2t0L901m1lL+Xp18vYHWEJzZsUBM7u4ORn9Ja8T
UTq7qyRR8835XvJExoW8N6uESsXqP5MLOhiSSgq/shbxS1y+9QPq06ziH4D5Bwyb3OMCEFTmQyQk
ELS7mRhi0OV309QDsKgSv2ZnAJUGnIWnUaUpLsu5nt2acnY8Uso0wjjITiwfc0nWwqH6qLzZaijw
RiwFNd1NGCXN+TM0XFnDU8bjROWGHfZLoKTuzd9zZj0Uq7rHcw/+1pSzlJK1snCn/edH14mV+dfm
73fcVNKWS9VCQHFt9NMXNOGCUrG+4bbmtAQ54uqdm9bskXYrMjbSth1rAKLER0KTnM0+ojUkPZ5s
NGeggJGYipJ4hOScXiL5PUWbeQiBCPxwcmMnWXgbleOEaiNFqZUaZeVXJmzflDmWcZ/W/NZvJETL
j8CLyMxDD6prVZkXKF/+AnAc1a/XcExcr809mEKS4I8TvOA861YsHgS2AOtmpaZyjlpxtzlbq0aI
CqM0yb2couSOGKUmVpWSz8MuG6dIn4Vf8B8NgIGcFeOS2I19RGBupVutQakBU5Z6ILuvL1NKCRNq
V6/FPuhv6+UAWNbtWRKKXD9dSD5BS+ACODBOBLbpAmdaaVQ5YbZCdRH5dv0191ia0fF+N7FnfaNg
rP7KLqcbSShbUOBjws2+ddBIwaRYa8WSrj0TJVb/8GZSZ+Dum6RQklY7sawQCbU8x4GWEwq2ixtl
diYVD3ZFNU6+ijLeu3wujpVA8GBr1eD9wPMHurIvwH8rgDV9iqyZMhW5HL9udTTv6T4Ysy3ePffv
RVQZRaGTy0645uqH0NJ1hVKg/4CTC8emNHdiPTpAD0YTY0285Oy3b+0h+GaHuenWwH+5EHo5DubY
kYB7LP3RQuDoFQ1bCWeAJ+Z4uFaUqJ/zYn95vtHrgfaEcgSFmdJqFkC/LJo9ehmc+NDwUrZY4EoA
8tO1O2TnDNcbeV40o/mUVvmDPzerbIiy28WOD8yheB1rd6H/c74eWO8Z7PWvBRQy0fNWZ7pZiva+
A0vA0HS0V8RwMR4LEFvHrhApiOSHlmr5DfKYgMZLBvM07BJEKOFdK51BXSucP/VChJrpGNqiZvpl
Gm11fniGR96xJejph+FPlz6gwx5NQZMyN8n7wf6rmjghmbuNYgSerpH7Tpzdozx3q9lb1/HbdocW
pdI3uSZfUv/BzcoorroOU4GXjo0bNzhmgS6XEjAIAwZZRmXtW2iz7UZQ+Afn/jQQsPOcZ534eJUN
LYllxz8uxHoRLT/dAqUKeDc1tvdou72Vs00W6ZFwyWrQfHe0gPBDl9NbHenLkyhKOB3a9hdFqlh3
l1P50NVlu3KvlkZSkeCcWRB/u05rAONpG8ugbrs24vFw0O0aZe4PM4Lun5oHFVpw1X9kN8BRzj6C
ci++2NXU2g/ZSq9TNMlBmEFvdm1Q2o5eINuhBan637P5LxtruzbbtaUL3mHHVMdJqgDy+h8fOaNY
cc1KFVf4tD34dz5GR+vkYGaMpwroZUTSLx5h6CfNGOmKYqTVSnnsCL5t8pz+VHTssu5BZ4Br4PbB
hyl8cnn2Q3g/+R79DloJN3x1l9jVwFZn03ahfxRM3PY9+jc4oeT9wwOPijaT0AfONNoIngzw2EVT
ZNSqK2fYBFzK8fSszxpUfS6zYFY/fVhcoWhFAsnyr/ea84r4NfJ037MrK9UPqRhUryao3t9bGkxI
A5EhVorPn01jI0mAwNsWZ1joINkE4UwXUq/tgY/2ZMvTwEiDffPKCMH4yCyG6+q/U6GKK9cxYTk/
Uj973dp5V0WtvTz7ni0Cpv3UAfyNScu+5T8aNTFhCdd0hUHxMGZWrfDZnDLdEZvFdpFLhsNa7SHy
NlgTl2wP4T9gnRm7TiHnoDhqXzePpSAguDu9LwzQMub9DyfyaoqEt2Oth4qwyQrktr6zX2MCObib
+JXpadXygMo+8iGB2Nwa8orS62TgVjDL8UhQdWc7RJWbSRWL0zR3h7uxRN4k0hCWA3DGQcyfCND6
WUdT3vwDEe7o32d8U8kf2ZcMbe0Q6UmYqrR4qoaDgx+9tbP1jPfUlyb1AW6JUCedDLWHAIzl/XkB
v9ArJzWY5r3MNx5/yEzE/urkm4Iwx9d0q2k1jUpK2RvyroFHWOPooOeSAgC1Fw/8V3UhOMTpPDBJ
kjI+Ero3Ngknv5o/D4MWs61gI/6nDgnX18ddzYQIB9ZMi8kOV6NmmWJgUKNtmeddneUSTLSUvldL
8VmCIrRzaTKCSMzpfuJV9XIQ+0Eo1LcpW3eM8/GfaRsIUKo9skTql4tyHkFYuSk95HtYObXqbqcr
LGNRNgzA0aOzJ1Fq2lEmLkcrpCblL/yEuoc/eVZl628jnBouZ1FQD3vz6ccoJtkmYIsMqXjD9h7B
cd6ElpVL8HFQl7wm67M9qn4cO1JRzCV8Y6WzFiCSDGJ4m/jBBSnl6VYXY6TzilpEo18tOBlUkT7C
CG4+nR68WqBMsr3KQgkbZwJUArG4yMb0AlxOXSc40zYA7onnxIHbI+MItoXHanlwDS8PgOn0MlgF
H2QDw/4bbdVUKvs7OrSwLy7EbpsEdca7fodVDuxDKRhfdcKs+cdtFeZnUCfiSvNvJoK51DTpb9TP
2zuP7fHkNoUaTax9mQ+OXJYF+xc3X70zeXyEbuprgmE7eCx2IWcvVoRm2O4voqlRxFD3pOveY2Cw
k7fhUZ1KPvTKBeC2C7pGIFLU64Ytmk0AKEoylSo0TSz92eHwxd+dfvT4TG6HLGer5JYxmXr9cVrI
Heb0SHzUprIel2psEF1V33kxiJePdg6oSm7drYp8io6dhO304jz0UHVV9th97Xn1RTM1D9ao8nQj
qziJskLPIG20Tn8soa0spOISEP/YYvCQCwLIKq2KRjwUlHDD/AKucHuAmXrsuwMKn3LvYQfFUwtQ
37ek9MgxHG6obWV28X+6JyWpl9g+GwxPuPuconUmK+T5+Xhl+irwWoR+gUOWv7uYAzqci9dtfST7
FRWSmuf/3idnhy7BjBoETaZHbK2MAc9lMcfZ++cq9gxSdgU2TNzBEiMSR9eMc2RvcseSbzo3Esk8
7TPtj8aNruSNdAF9AYtU9wPHdosEBd6oUvgWtqBhfWzhL6Hqq0X8KvqHel8c9gscr5j0fnLIDPjv
NQSsMFT3JBJ5+3eeL4xvhp63RnBJ0A3JOAR2YuJUot2Io/uHR2A3aUwNbT/bFLH7KjtuJNbgrded
EQsWzAP6naZIKLfBJqM5yZlA79MxC53Pr0QMCCeC9PCVJgGBtnLQbFFwz2Hn67k0Par2DkeSUgiQ
2r4oGZaAOuvTTueWdinnUfxY+JLxcNZEVzEKIYtWJIeDKPq9onX5tgQ18RuTMVMRs3TbKvICtYRV
Kxqczi53X7Wa39S55O19MsehSfOCJxaP0i+SSpXFyBZgAJ5JYY877SdGzBOHNFmRvZT6qS9WJTFi
4V68ilVzainbCtdCxTZHJ+4gvdvE/HqD6wkZa34g3QgkQ3lRs6BQEhJ+8YM8rHjlG/jXb86LVqWb
TOXIlEjW7ngaBh9FMfXSM9aLndDitmgm5CdiE+9L6CBlBhI7UjosA9WaMSX7axGYwNtwN7nEwURc
EqYaREU+4m65R3V3g8NtfYz9x6LTyqHFrStEdBGZx7n3zJbkoB47BT85lg+D0NZfpBhRf6I33NuU
rsKwiC9oghwqmsNUtQbG3yhr9QaljhEFSh2Z9u9WE2CcjnmLaafGt/WfhrTnQndC7k5xmNilj5+9
o+ENK+VA7Cu/38KzrVRsdOZxw9zDUFEPSGUZ73kNt9xEkWMhrtue06GCQkriPJDZDlFFh6sMvjS7
8nz91wulJC80iu8Evz8xvNTzBvSsL0qlEpSoMP41QfJXQmWHc1w1xeyqf91zLo1SkG3fT8XLKQZh
dK066QqSQ+iW3uR6vWRNlp1Ygn4a9vtu0Kcnojawkm/x6ATE2srTVBs3XytcfayFOTDvVXr7JrQ1
AqmtiAhvYVHyZq6Dzd+c3Kpssj6qk44zaikznej3gAnGLFY0wupqNpTcStDKB8nYTNgDDRFBpf9U
eYLKPi6880NToAMT9oJCtJklk7VzSBN3bZ73yB/PLzwEVIvHWkCflch5sya/1xAAyQJj1PlYngaf
DM5RoziqG2szGsTraMTLGInEiiHQ+Iho5JZlSEK7Gpuy5XBOAG1wmmKFHJkUBV0ZbILRNVFzL0Jm
WySzTDMp2zdoyZ2y/smJTMdGiydXlSLuziFuTZt9T3uWbHp1mWnn5DaMhXplFEH/FYiy7UfvfHXq
ro71UwwB9CJpSGD/+tapD2peKjnBrqRDjvwrizbismFKz+sBc2xm79vRGy2DeFu/hjjAf3rlgxUq
z+5RdE6O34Zgu+gq9s7SxyZFmdA23jejxS60V22WUek/9oTq3Sysn79pth7496pZlDYAzMbyJeIJ
PZPfz7lmDv0wM8y5j1/sFUwnox9hcEP51X7agvb6pqDGr41SlD+m9DZKyiYxgeR9nQgeboEF250h
hNqnK3+hfwGPY446oM+o+l55llyJh6sI1LOpp7s8zOnsfGCgmgvPdRMcI121JBqlgxSDt8JdTj1v
4qcudwof/0Qub8LZQVQNkHjARqEV0acjJ85SBcm6GRqo+02YhqIZAnOBiXZtT+AjBV6ep8y1xU86
5MkSwchUTCxS1PnK9jz1/4HqJkHQKIximb8jmOpmlZuzg8gTsRxvg2G8on9oG1jGUpdlELWILPaO
xhOJ3/SQ+0iq42bPKb4ZiFjVTB6V3zWlUqIIVaGkeygBIMogByEfYBmV4992ETVprY/wNY1RgxES
A6h35PAh6mfYxhAmKuQQfLBudBBmSEZcYVXG9JjkOgp+kWe7XHIxEVL+jn1z4lqoaonlADVzSDuQ
jXJqLCWAL4ruxaR/1BNNeZW7frRDvNWY5czEIkPrT3s0g6YJHZXSl88qTHncoMSYt/7H5pXKUewk
j/WXL/5qYopmcNs4NDgs9g3M7Ht7ojMC6yLdWdr51rbkdYXBJj/ronCRNkVgUwsLJwf9PaFIzVib
TGJTobLametc6IjSN99n+U31RwqYqpm1TUKsc57ULUv3AYFcnS+BPlj1WlzIIxuCq1he5HKYONbT
JgS91Ikz7sUrZeQJyZojrR8nsBOdLYIjmMKvsCgLNY1CptmAc6XPwwogpxLNPIYyQSOErAVbFT8T
OkQ6nNQWWg+slW8qWxQpyIHzxApnChYKg5NUnXRUCHRpANCnmE02f0gWhX355WcFjqjzOR9sHNUD
yRQOeSlUb/jOYKsNgKV/zkDR2T7D/SJpZy0OQHqxe6GU5qzizcHLThEohABaZylT4L+vh3BrVdTO
QrPjHmy0y7QN+q3y3dKhsyVwXbl17Nbu7Ihmw9YAJRof1zR7yuJezJvH8X9jHEiZzyA+pSC6ULEp
9w0nbawhqIeS7Ssj/L89jIfPaDGqfvKnED0ATVkBGPSqjr63gJmMKApZfI+3LGNQP8FcHvGgwrdK
y/S/kkT+PgB7R8sAedaAGBgC+4eXTYcFvFRJR8QqBcsLodchSD/P8Mz4+nKXjZYkDExEN6ZXvnin
Dzln+d6q7JIM8AmjNYTXpfDyJZtHCASPzi4SHFc37U2WU1OXW5XDpxwhSHSVxzMju2IAcfalBnhR
GY4t3yyljgoBSm821gzl7fRO7nH2IIFAKvrlPeBomOlysUKDsYbQQVfkGJLUvv5lbAA3s65Pcgi3
xAKgxINhnJRJQFaH5hN3NH1IWsUK5JKszR8uhI2v0JEQOkkV6vNo4m0ZEUFUCmv0jUMoWQ7FZmlC
YE0xSzieLyvbUJripdawh7slCxOKPeYeydCA/Y4/9W7L1m59lpgtUDVahAHcok+Uk+IjKs6dh9LY
DQ4ohhNzvymvZ3voTGSm8vDE4RwyOwKlHDG7vToUJ2d3WXFqb16j4TUA8ajJ91G8kS7gBemy4Nfx
Z/Ifh6T6zSXlBzgnD1BjzlqKVsX6fQsy3gm15KPu+qwZQo8HyXON/VOrqFXXBPUsGrgJmbyPLKeL
FvSiBwYCCjrgGVG//StGK18TLjzUPSVyiqnpdIqwaW352QPV2M4/a4NMLTx542gHPzN6WD3kVDHM
GfUDYySF/ZxjXFsOhL6Eie6U2KqEHYt+aBDKDrLzz/e9zE+PfSzOQ2lgd0IJJFn/NyUzevY4MEvR
eV9jksNdoxF4mc4rd4TvLK41c/qzlH8Z0t+kxhudR80bbpfheyjZLIp/x2MdO6HVaYA7YsBV/Usa
q5uNaNrn6VwVXAPWkST6qhV5PsCkrKaiO5gVirxJuF2KaVu8C3ZLWrqPxV9Rcpg1+LAKmjAKrjG1
y6lSRbzRqbU+u2sG+Bw9+tG7Hl2FvytiXZWTEriYVHdwW2/697P0/NFK8GnNxvBzdge84Y1pmwxP
h0Yd5y1X6CYws7iSjPLSsBBci42Q3FXy7lnQ7b9ACUQu+eDZuaSjOHqRW9J67GfIVuCfaC5bXvtw
prlnOE/ZP/IFDRGGC0REmau3vYN52fM3wDEss5iastxvWgESr9Rqks8eZoGlyyCJMD5n25jGhAfK
a7ekLeXCue9RtoPd/PIvufaRJn1qj/ToWbJ0Wc4n/Tff2855X8gR1mmts5rAE5QfAT2V14s32u0X
cUTJkkBavcPRrQ5MqMWCmXbAGeFwfQzXqA5gJEQDaPtq1cKcT2le7cwY8eUk7KFSyMKstQN/UjJq
0hvhroDUWbR6XkkxAzuH/4wmXBpuCVq89UeySBLGLiBtkRWTxNwXJv22F0LT/U8M5FW+/SgQw89j
7lwCmsFErRX4K3pACdnmUwV2vMVuZTMdvRdP1jYD+dTiwqqmCe895YDQVozmebGXrFsNWe0eBjpB
hqwq1sY+c+sITPX2JqCeS069KztwXu1PyCWQZQ5T0uqlDzdUwAcdXhAH65P2+UJoDjwD0iSnsX2Z
9uXUqFnNcjOGYO1iHanrN6zkbjBWCP/CgASz2So0dutqlIcMfcAMBqeYAOkFJfgFVVp7DHMmEVdG
9+1/2Q2iwp5EnSy2KcoZIDnbc0soCWZHyJ4+P/xV9TD5uG0aS6HTStIJPsh/WMyUnL56jNySD/R9
9Sa2o7oAHTF0eQOSPd1qgZlYPsJEfUF/TwG4mZkmeuQzHTAO9EFNcr2FFgJKlXnwVvjtn8X5f++W
haqV9BH/jOZcwTX+JUlvs7wnK9g9YlEU+24nBlpW4GHIg8sj82j07lh/ZkAJUhOq450gTGiuHTvF
mnWJGspM6tig3BxWdBacRWoDZBbOk2KpIn23HJ6LAbuyzvSx4ttMqVO3r+u3RPjgMJawujx/bXFN
iB5B1w5PKV2hc+hhfJCcQIvbc3/91YsCX1Hk+9C3qq65UEqlHtp6CjzqBejvN98ePqdtwuN3SdHc
j5aArHmq5P+3L5BjK1qMvuKqWSVlvXE4dxDwBWmkeP+I4Sgh4BpxlI9tMxK86q2r7UOfERcEigS0
e8TwEMPVmYwjayHl1wCHujYm1/3wr3zePp+JXdfO2kEmJHZw57Xj4ddDoH29DGVyIBnltJnQXr66
TCC2s5Ziflik2E9M1WIKRtSY3ggYq8Gp9qVrmXLomSSaGcVoBofaWpzwMwhivzanbsioGKKCNG86
AQ+nKuBo/cEnkQZGZE4O1eSB3lJGuZGKoUrMfme6dTcayIp7kZwDbFoPBS9/XA8ziNu1LiPEPdl+
DBPXpQa+d3Wy4sWhGCtoWmDX2dUjKDJa2QvtL/TZ6mNej3CrL87wBP+gGXE2vdlDuW14//CnN0sm
gChhvFMBPTp1o6lFyyCzariuIWoEs8uxG5FNZhaBjQcurKXT+ABq6jGHtZwO5zny/7NLdfSutN7q
ErTD8dyfVhA+gFf3m+bv/mQsgYxnvdgb9DyOOizd6cqQ1YValdY1zGdnZ9OzkTnRWv+M03rKhCxL
O0eM9z3QEPiyWAmBklOtGQ1clQ6R4+yeXRz9/pR/+wecgnQt8vHbr6EqQpKYADhfOcJzKnALJSBy
vfd7am+tRxf1K+sUxCoPFq7TfZLQoHVFPK4y5klafHifW3t/tdKPiV6XT1HNSe/szfMxeYQISvEk
Iy1aVJ0enMkwsm5N913OxEljHxCRDZBPdcqvIdLcTFFMygC7ezG5gv2ehGTpW0qbH7KPAO1b/KU6
1/TBzrqqNPiKSuM2akIvzPoEoJEaRrzXBbjNipmU3E4q0D6FiU5iScYCkFIbaZYy2xX4n6bUFR/h
Cvbyec9QHey88BcX6ruNc5+t68qsQPD/JhLmJNLZmEVMcTi22zu1/c2Vlt5I0wE0MMJIS3X0C7Vh
nyqC9jsjyMXMqPVkyElRCIP+PsoUdjn3egkq6S2q5LpsZf2eg7ZGM/Vql0sLHbe1CozbLPluZ8Om
q5Nr21KgZm0OO4gdb6ioLdErBrOYWkvyvsa7hZhuas87c2b+w5RWIGo650Bma/Ab6zGKs4UCdNDf
c6P9MuULzzwa7G1GqfPvw5St8g+RfCpswQDF/txzx3dge40mQPrKvsvM5vpkGSeas2yEMnO2YTFP
8srkBR1qRIxtW3ikSxwCzPwE4jINoz/mF+lug05K5rWxhzakQxgB+rJuZagn/BvQ30ykkSX92DMy
g9x9ifNlUe3nKKvOsgaohrU0yEKKLixBYVSynN84+dwZd8BXyK3Kqll7XC3hdsgq10iONvQhbdQ/
9ZFiCRMUAw40iDtm8ps6eWats1r6BT50VfCMZgTSdoaOnRPOf/STdToc1kOZbUJqeXTQ9xy2S92i
YMQayr5CSAvmvVca7NQmQ/OmHvBHyg3X/ZrlUV0acBOZ5empbAcW41/CF8zBz4X0N4SWohRmdk0M
Q2vzBTY5F7RfFcb5lx1ux9HkohY+V/5pOtNKW/jpbGRiQdmXDls/V6XFkDSW6GGMgD2b7HzYJgM+
TF98eqT+ydKZlJexkOfZ/AnQArs9V1Lvyh9C/qrd/A1tDbiiGmt/q0zZa37K5lYGZoIqvoFjh5t0
VR9Ap7cSPUEdtLL3nKcm+1rdcgdrXYbbIu6haPTQ1tcHQ22JbYp3Pgx4T5X2vFBpecQswYoycxua
kZjnt0WGI+z2jQqfl6yMc9vRoLu4Nf5NlZWoIYeaK3rqB/oMQbGpRVI82iAV1W2ArbRJZmhahd8b
2qa1l+ynsE+9Vbdnl+XX1ljOvj2z2bR3KHkb8CmwDS8kypq3ZNaSHg1/9ZXeLbgt5IF05GUZi+2h
cvmt+rY3fMW+Ly1l1TiIySsfQan45G0HyCFPgeFWa5A+q69Y+N1j/0PYK1VENbX+e9xju8gM1O53
cFVS2a9hHv8saqRHfTYpgpMC5ivZa8gIELRXYhx9PGJre50HuiKA9e13ZBwz26fP8DlOLQcsLlsY
862IkEgMmrdxz3voYZso8fTQUWVOFVtr2c65gxWT9dQWb7zeDbbZpJUT5Pz97RmcWm2vMdx8iiHB
3llMvjP0Ems7mR8CuzzLlnQFHbgoMfYo4knHAHwnkWx6ZgTAIbMMidEA3s4itbWAkOkHSzXEA9ro
uAhV5bDDaLBdFZbbLKKp6S/wPNylzcVEj0jTwPjmaHaX2vpRzwpkPXA5PlxjYCGApYzQ8PxSjoGa
GBkGowGZjoQmK5xplHClAce1N3hH/YKhiXPNl+vg3V7KR9l08Y4D3moz7A5mNBZqkrz4q8lm/3HQ
o8FZGx7zmn5KM1G0+5VnbOgYRVpMgfKiz2N6pOzcMHm3xny153ikFLPT+jrq2rmp2nR3SAYabY4o
0L55txYHPDpKjZ8mif2JjuxKRrvmYHciupf7Wqbmp+WQlZFrSp3HIUh/XaM/oxEu/v95UpWOqrZZ
QhLFJNXsWE0Xcusv7yWUlULYI8K6mSQXt8lfXPglXHEfY1Rl28DugkKzJUswR8CIG7uZQ2cbuSNl
KFvRW2iJ2igu6HmZEbtCxn0Bhrvm2rYxY4N2XaL9hSGXQql8cgZifBxjNHvhE5GWsNhAfhFolU6d
fsBwViGPUO7uXaUkIOG5YZsn9j+P9stW9jP0hI7NQImByE5OWo0AVqKObUtG2xIRViVcS2rfBVAz
79QqrjpR35BDBpmvbnIVIgzUkvUuHOEx+opYAP4Anmao4bG8QRlpHe7Dg2fD4vB7hrT6BBnBSOwA
IeiQag28wh6Nl/0ytBpheklCio76obKaN9WGSUo9nu07Oppi1LMnJMjgLfNeFaIl0hYxmTnSy5Tf
NqL+rAAzbh//LdQdN00Ech3gZUixK/e2z5XPF8aOcPSO5LpDYYxQsSmHwMOZtcZ7ZS1Tl01tvnQ4
bwEovdQjq2+zkytiprF9hcjaBkIPb8k1Qwz8IDL07b15VBGZLdm9ldCoCkmrnu/CsGGE6uyYFk/5
iAtN0jSTH+73MYKbUPQO1j6/pWfdJRxTVK0jrf6L6UWjZJXvxbSi/aW6mlS7mm297e418MLhU1Wv
dXnkqboZIqf+HmAkQeBv36hFNwWQFq3OOQuejhSybIpCzL76+LOYpDBJ7sslBDl+pLPIcSr/51Jl
Qc4ZB+cYJcq62DyJSeGtmNZsPflYm4kh7Kz/YzybdUwdi1UTK7ImvuaQ7l8Pr2PsW06MPJfhvoWS
WG5OxHUFwt9pToUgvm9ncCoOu7KucYONg/19378y2HupEvgobVcnxG2m+vf1d/dbYNHKPxnU2Nz3
PuIcga7G/ptLfdjNGbRnPJN9thjPodYgvlznR+oTgvDjXgjYPuhwVYy3KW8GMcoIgDiHSQcYCP58
hQXriZq6l8oZjfCbx4+4+A2LF19Hz4/rAt16EUpCyt2RwM71YpKff9gWNvYoeMz5zr3hfED/lWDz
t70ikqLcprl3MySu3l9GW2BpD7kqB2rVWtkPTplvsibrPHWP7G0R3YKpXiZQj2va+Cc2o3h1WXY/
s6P8C/7DiY9cjiDBhzOVHJ1DULWlLb0RViaDUX6pyCuVaRwtzp1QbPph5xXj4875xCmlWtDCUyOC
fkxWOqnjKJ28jNKMriGjssV/F2FrgviSl6SF1KlxNz/UKz2Ym9i0UF4umCxyH3E8xeflZYqBzVbo
+YpCJSzb4IePaxTnpEcwDwY8H39IiELaeKJHboinpMyka/+FApZopBXkwlLeQoKFeAEMV5fLlDdC
+ro0oAmMi1Wkx9jkmDWq5tgNhAXGrFrc1Ut5D6OIQZfqAvqAGOATUfYFgbViSY/GfZUYQLM0lvAF
QhdNZVG6sYxNu2LQ38fO890FxM19oMD1OgEQr0kfHr6n/HgZURSju041UH0TIkY5HIEuzs+FIu0I
6eu+Z2iXksZFNsylwPHlbzcvDqIyoc4kgQnoIT2J+TBBEp/MX+3XVTJOL5vnrNEqHzwMG/09DYuZ
ff26ftmBD8+tnYPCLrsjwN345HRzUiAhWD7ZzjokrO7QpfStGT8ooajifTc2eFRBTAamFf6cujol
ySH4jixCELmv+YAG3xaRfWja4fCpMdS7LQOZLvoPYP1A4iFOGJqbQGJsOetyPiM3bqY0a5AW8pAX
55QzjepG03k88R0YXuFDP+pHfbxPKTs23v8epwZOu90bzzCDlKqSxLZbAVS8gsJcw7cAIjpWhr0N
Qt7o30UD39Fho6FGohJoFTGGm6eTl+Pz7XInIl5E6tBE8IFlUw9ODSQJ1sIsD90lI5718kuCS4F9
TlIZKOZmW4dhlFhzKO+jmnlK430SPZCsd4OAHm4bG2fYcO6aqVSYJba5XQUcoRYOuQ7LxXHj0SZS
YdJvMo4OkwHPpsxuXSPYyG0fG5FCVYShSllw+MGBL28yJdS4pMb66dE/dhvdmL7jlTaJKAA3kxRa
HSpCqD3Ag2/l9+EZrj39q9MQHESfG8CpJYJuEGXY+MmByM7WTI30Ng2Ml9mFYZxgU7ePlS30AeVQ
jXhzN0t4VkOuVAl7N+NM2XkFgL90idsWSRpoVOrjAH864s6bgCXP/w8JufFTfHhP2EcF5AhdEoBQ
J/XF25IzsjkI8HARXeKmTapLsSOMpZmlDXLiKXC+TSnAxHcXayyGgLKzdwRUpT6nHdTuqVNn5FA0
NYC388meyA6dv2F6sqbRuTeYcqHcBMZTrgZWBvqXjkD9HmOuNfo6LZfkRZE4zZWwIVj/QQ3Bv9TL
ppvYnhyvwFfJavrTN+/SnpZNiWEpLra+GKG+kZ04iEwUMj7/VCS2RUH9Qb+gnt8bWl9iO+Ft0VWX
Cy6tsiYE0VADErRXAEiUh+tHZxdZLPXGVEVl5fHaQgzVi9+/qnWvhHJDdsCQg29HmKQuBxy4TT59
sI50XJJSsiA8yzMOokiZ6Tex0GiIC9bDIxei2e0IGdis+TS5QzS8o0er46lqNK4dgoQsSCbwqC4f
S2OoQjtcZwi43Rha7+lKSiZQ+vH9GlmsF7fSGggWRJNYnY9azahLGg5df8sioye3tZn/IcrhWGNs
9hxL4y6UOr2E/1+7nljvv0KOTyeh2Io4Qbe2BjEnk313NQDI8EkX3LqDrO55H4+cjPcgC1m2NfxE
3l2Lh3hOLG9ryRfIHtvYs+s5ZaxeZ/pZKDCcPVHXHUmF5W1kY/j2o7A0mqMkjU5/iC5mEiWhYKZM
ccEUSmJXpiBugATABLeduJS/SxrMD7f1T5O0Z8eN0FGk/MlPc3JpnD8s9V9EciAXU8Mzl/1J1xoL
Dkk+rdLeq+q7cVyhYk9MhnKnDfKIY45OTLdmTFIvfODXo63+dDYv4ABfR7a80MXz9WpexpecK8Nz
WtReAymmjTGjlNaswKr33VySSPr+3MdX5GfbimfSF9M7KjCjHfl3oxdJXePeaagEfHRhXfNNklYx
XBed9UrRQFMFCSuDxhoopmdI7esYUmaVhjinQv3cYP3wKq4+KkZ8luQp/XiTWz+vjf8ylQjQlew7
9+z01Qvbe93H47X2JKH7l3111k1FsZVg7ekpoxR2IumkYKG+rYGRu+RMR6yT3oO9GMU+GJjhJd3y
ZzgUJtU6jumUrS0O065WZQkPqNPUWOJj3cigFxgdVITjnIU0R+/LpKAbd0UiBXeSiriK6tWsA+qF
xPkmdEFFZ0vzlIvxBF92pQpvxk1OctVCYtdOh13bWa/C+JszrSEkCMJ44LYXeYZ9URJ0s0BgSu/V
1470WroFzRCFs6Au7inr5mO3wCUCA0Ru7989cF2I576eXHAXnaLcIhQi+ctwRy/ki7/XCVrLRCKF
tLOdEmTkM1S7cDVk6C/41fYSyzGuUCIJVf/Qvll3mcvqksfCvMBYTG900xdEh8X9WQttDU3/CicP
SR5L9niKfsZ25SRe9n/xulsZg7a0asMK1orsdYI4nIQVJsQeW7UrXnUlw/GI6DBd3O9cpptzjQOS
GEHf0EarAojglm/EpdRjMsTxZgn8/TUSUctRqT4yZG6XY9es9hZ7rGsXNpnNhXglA866PnGUeq9F
xJp3Uc3b0FBe2YDvs2R8XXV6OY64W3t/tkoBNKYdxNvMQ6NOHmKArnW4/XIDDtF7P6qFlAhPswMR
SHLUoWiuZpbxoIJozLkaQcniWAbIOSY4OiwGnlk7hFhrAMVxWVaPTlyZ5yvoJRxeWw3VuKCZV93a
T83c+17xQX6bBNOun1TJ6ogkEqBeuAU8yQHD+IiDfTwLYyEh2ES5GMllTsSHFCKrswRlOy/kcl3S
AiEOXjtinuU7FBlFipgxrmE7zMXkNhpLXFqOrB/sc1n3+tO4EFb/NNYNZRM11acxbzQGiloO5Ima
G9o4e1dHL+1yENH8y3hZuDT6HVw5LYqZOWwwhNXJ2iTE5+ybT0GfDXPGSQdMfwVD+DVOdocA1CDt
s1mLCb8Y796OSF+AqCH3a1RbxfMFk6VtPDa/mT17tD3gZ1EYE4aBeTh8r26FZUq2OuoFHxBf2E9m
Vx8vuYvp9xUSjLO1Z4bduDqiKjANaoFomsVavyGQ/Z1Vd2PtOmCZ0hXDj8iUXjyBaGxneVa14G46
V9s3IAMlc5SZRoMgF+uED7yNb9gMTuQuqLa7V4LZehn/GiSYn+AFohIpVq/9SuosWUmxlxayFI9j
eJqQtaDMal+vNou9NEY9poP5tA0C3vzVBbt/lJi4vGA/HYGhsfNTaKR5ud87Mke6LFibTEtdrWzk
8biSsmYybHLhxOK83TxfhyblGKNRpobzSkqJlMtXKYlkWRSUJqoPRzV1XcHNX6fqtv1F76g1XJrq
opuledgYbvqLTe0knE24bDqGvae1HVkMLGFB+hCTAj5reHWg6s7z35VBjRQBvqHQfa6LidHlcHlF
Y5pc3H4e7rNtSGsdgIuR+L8reWFWyJOUKBLFJ3PhIYPPza1cGiP8UwWyhMLgc9Cv1oVF5Kt99Eyg
O72JOfK9qVHK6IZqCogVIY231+zZKHll1sycqceznTAjx3wdSXmQ1E9Ely94aouIzDlYe2mtv0sX
Ed1KbEVJWb9XK6DtaRFdv52X+U5mnI23GsrFydHhf/bLy7kFyotZTn8HnYAG5czGaNGRzQhlyMFn
g4XStzgGsDgMnJK6lWEJwX1v3xkN/+9843zFBSqzZVxKS4EvnGhbj7T+5eNKj/2lKsgC47MO3eJh
mmaX7lYFaTB4/M6V8Fk+5NLB0MUBKWcX1/zdf3jkYWYWxHBi+TPjJ5pdJ4mjRJWLKYC3nKg4wvNG
67aJCxsCM60pKrJvA05v92LE63AIh8czKT8VLYGYcjNkh6tMg/dx5aXyw5078qXEGtse9ztrO/ge
ojQu58WiAc9ZJLSLp3yJESQOSZaH8Lgj00Z2LOLujfq8X69f/50fSclF+mEWbL7h6No2FoNBE8IU
Qx0lBtimljCz6LFXOdFVjRCjCyhwZzBZmA30WKB9Xw0n5zwT4qmRZpOWFOLDmbE4yBJ2ACcu6q9H
b7ujF9UhIiKwMLC5L+tYUoZNz+d6DgwEMGrXwJXEX56ofrXPD4CiI7VW/78IhvntqLYXBTOUpQpb
G8kObSOAPkbFYltPLC1OZLCcG8UNa/DwIa8hf6b6UuU0b+yT4N1M/yL1MfQpl8ZU+jCe/fj5BYDc
sw7SnmB2YhAYXpn/TFEGaiKtbcztPoBYoxpq5nF2xXwZEIYo4jnnj770AM5MVK1El4SiW6nIChDl
NXpptQUoD8xmAOqvwXz6hsk7lTGNUuf/FTWorzHTRY9+Pf7GI7HNxNF+d1W9RWQocEttjUPx41oZ
5Ecb24n38LsJhUeW4GxsgenKOmkRhu9/RYgxZoT+6od/aHrjRvtSZzU2G/HF923JbY3uaxISHrpF
DdysLEcEwtx5D4JzRMk/oLwIemD+Olgh6nhiEg+jENzOXjKLsto8DGY4mC6/hhrhZiI0KMTUjG27
TDjVQttRSW3QNQiLsVML+2ybkJlFodtjnwoBAT9YVab9QqL7JQ8wf2VxAgLrgXBzYYdWqpWVbRMj
K8vEDudyoCNgzUTgCwxoJ9EoYpt5fwoB/LaAOxF1JbBOwc23LbbxlfFox6t+51JsMJ2Kw/eDy39l
/F5D6YtxrcBnAjzs4U+FBNsG+yRSs6U6pgoEZWP4LgsFcMudLalk9sXlFud3pM9gulrA2YbtlY5m
t0eLkZKbnkkguuWAlB2uNckUfrhNkwmRmRG0Q1BONscuzmEsknkIGcxHDYm5CWUJyTIDTxPyr5rg
vhylzV2tbVxSFukjE4UQvi6/75x1OmZbXUjU0gpnF3CaDwrYE/y1LlbsBUVIoiSRKUx+trsezuld
mQDRdIUDj4shoMcS/xx6Mof55OnD/dFgMIod/xoO9ax+DgjmWDFp0mDpA9Mmb7Xi1Bbrnh9e2M/t
2mfHKcAPP3vbrcapI+9qtBhH5LDdW3+vkn+z8iJDKS4p7U6ThVuzwTCyfYhsjdke7K5L0nIRliH4
pjdysIfO2+xaKji49i3gfks+gl1oZ+lRyyrUmmpf+w/RXvFOhmR/WVXO5ZqCqrnuIDrUx1FUA/W1
k0li21QBtYwrz3PuXdpoHPTNYXMQAoTpupdav7Ss5kBBNo1aBad1YaOY5vh2Ty6Kxlc3wgg9AL1u
KsXed5+foJjqZ7R9adOGcFbHBMpKLdnhpA0+jsbZzUFaqbV9qrvMhlLlGwTht5gEkjkmj+MJyiDZ
gBNMXXkmG6aJX/s40lVx2lhEj3VeURmyFWFYMUVP4o8ts9da+tWUj5SxaBhB1htRigQALcuLcEW6
asIUmoWyGqTcBuU11AmeTsCSDAC9GEcZjPY2dV/AhyrEz2C8zEsxUh64toKQPqdQuiX6Ysj+HYiH
FTMsbjCiCDrvaj0V9rDMWdPbFQlWR/+8iB8aXbWpQ8C7CDRiVl1F+NoKzpLiUda/kasqAWfGQb76
x/J8mpDrOFVID1fHreU6aZVYbTkgPk4uCw6CSRq1qKA+qRtRnWWkUQ+IIgwLTsYSUxj97h6cQXYJ
rgp4gP9/DUUYHHkA1xUqTLKWqPIMoivLFkPq0F7aHrRhBGoar3G0x9oEZqXmrKo9ueDfEAYnbKiv
7mDOH8+W/VfT6wcadtRL+ymp5jQwCfnXLjRDD8XhEub4jpTjt3u/weVHFotRbOhsJlU3wpsrJe2F
5FRztaWcDpq3lXHsZfoF90+Rvlj0A1hfifWbEB9Z2Sjvm8n7CKoNWxf5o7RAE07p5kFSsD7DEJ9m
38p5aR33u6v7MM20xauyM7nXcthEaOpx0RfQcLip61gl/Kf4UyJHAb5+kNo77QxdXF2pFXly+/cy
mnA2Gwaa2qRiRJVmD16QwjY+TJ32g+AP93mM+NcMYWMXNLFzO5VziBXGcfH/yvEuSxRWVR0oS4rP
nUuD36cq1hU+nE9Z7wu6btRZJ9Os8cHicvW9L/dZu/G8lpKGYozDP5+fGYO++Gf2mSyvBplg3akV
F7A4kXy8b4iwPuiq9E704IGm9uhZn/soe8HOZjYith2JGjGlus90Th1zpSyuX3ntQxCaaVoMxq57
bWmyakVQxZaHW/mzd08sg3j9yBAsrVEi8fbnYPgvr+2vln7ZRa3o058nha+paT5b4BaJEb4K/095
+07I7rYPnUff+PLw8wjSuW4lHPLyS4EGCObkTjFCa/PGPz+z18alqz219sRg1Vd6n3muG9VYBuKN
+mhepQTL/VQ7bHa7t7c2ryjgGT3tAkBxnEySuHW1Q2rdD9CqkaGdIlCFuCKIQkSQVBlY/H+mYwCa
dyMZONPqLMa5nANOqJrIYaGN2TgW7Oul7dAOo7MMW69Jt0oSr6PiDbxe0lXbScfJGJf/kK5BoNgT
cx5qnuJaE6WOMxB1QnQ/kfXuD5BPDtxJIhnd7zHI3hw6BulOJfkQhWLrG9cZIbdO7ORo7gKxPr8N
5T3KclD+iK05ek5U7MNDFuyN5EY7Grv56xAXLnJjEhp9BwaaitKTe0Jwt4UTPNxKH7x7UkmeBJOK
+tL0iDHucpmp8VLaZcagvqcl4IpojWfRPVziccgd+M58QfQNfg8JAhPlUKXvqlQKTQ2AaZg4CXeX
Oc+Rmh42lyG+kutE3Kla5BIkb3JmYpL6ImIWI3wLBe8+hukwsa/jw4CrRbR8MROpMbIqGmQuc4KS
QU9Pswe4LJ8XRcnMOls0Xfx8w0nLTi0jtvQHJOea0lAJ7l7SV8IvXMjphblLReYDOXEgZ2GOzRfa
bBR76NE6gqTM8eH9OMHb//bSN3fFfCdeI8DmSyo2pifLq58GASweVw2KDEa54dcZmhM8IIXkpCMm
jATLRyRwku1UdHTDGiN5BpukgBgMFv9PgTQWXyi6MmD5mJ0Gw2HL1JRf0nuAbWxhqzfZGlDxRCCV
y7ywgipV2l4+CJqDVW2KrmLPgYSSL9ZG606DAhXGObmEXSUSZBTIheDB0rqLW/GQHKHv3G/06tJB
MB0kG+xCRClOEb5tV6ulYw7SJBQEz+qmavEO4nxJ81IpCpE6Ct2QKXBX0l5B0PJQr1fN2NOseNbK
yuj7G72lZKanMrbqKvNp4pArzJBhdeFAdYcE4FJC/I22Nu65M7iET6jaVjAfpaIPD4OX4koHqKGk
3ilLY7nC55DVYmfO9Bw1fBSVa/cgB7ye00np3O/KeaCuW7trJlysOyyhTDf5AQOoXb0Aci7F4l4I
YPf42uSnLZsQ+TDGZuyaTnC812lgTM2tLvaK/9lDRHsatTXGJ5PNc59HrsiqXUiTV8OJ/Yfe4Eik
TtvDSXyTtSFqKOYD2mTcBadGJIVeV2xwSg68azz5T1HTEkBRgza8lUq4cEh0cjMlozlIpJSPKX0F
VcORjjbiMYQ0o8z8BpruInE2inA3oOBy0LRmiHOblSHwJI3KtXR/DGVksNH/3pgtlPhscFdF3CI9
1JgYz+fjxwHkFjDlyjG4BW5pVz2sCVbUFUuw7O9tlfQPWiF717KJj0qYM+IcIOKRg3kekkIAp+xd
wzl+yYnD7aHO995h1NM8ZEgc9FZJimZEVoYiUO/RRfylnIKg6v6H+EQlxjpTr7ayej9r3HtlCTAN
qUFNSURn0RY3fDrk9X0EnjmvAyLW5fmK/LHOJR7d2t8XCfJLlGWG3LfRW+9Er9SxqTv9cgEq+/lY
vMd0UgjEIUCFzsUccSfPI91lZdfmehxyJsbHNqVm4bKhwwhb04OQw37SeGt0KvOv6x9uVaqoUUr8
wbtSfequZcDdDl9WJefSYXDVSxJTQUz/waLYc5mRtEtPLwE4rsvMjmlPMzy4qTkiZqdrGDz4lGtX
ZxEFIjOTLDlQM1O8KRrDIh+uajPN9Xs8AvVZkmBCO9Nibc+Rf/fni+hcaenvhwR0L/gQp4s+yJj3
/uEwV3TGGZhhuqdXuNiT2shHH2ZqJZUNyyqZcfO6N+JmXt+yxw2dbrT/FbmrCrPVE007OSJzS2UW
dsx8lF3GRYc1pqDH4yHJBdJhvDcQHBnIHKsF5DY3his4JQ3kghXXP3Ieur+ZVV/Y5y5+cYSqMNJA
TWUo3l8x9qiyWCkne3oEcMiY052WiE1iO64iDT/vZShteUageN7qMj4BrARM1vtj0uWd+oc6Vw/l
xAokAPzVouyvuuEsy7UtSnPX9Y7K5kmD0nZ8WHymPZDDCGKRh5fFNZYMd0Z9lc6Na+rXwagJlMAh
BoilkJEtWAqbZG4R5DRwFUAa6koTWgsH3BERIdsiQ8GYLzouwdDGl2Dk+VVr8mSxIPvNmhhfWDUB
nDjbtCP7QzcSxZYcKiBqGZCEF0lMpB6bIAC2qeTH+5txDZWe4TfuJIyggFAp027RZJ2nfUOWwioa
q8SqiJEWQrAzMkEGhMpts74uQW1uaoPyiG7T5Ry6XvETCymDZEA9+EBCIZpwQG1kByrQBihoJRhf
PepcxkP75sx6S3kCJOznq1Y/cV7A9kcCOV/CAIszByYe/56pObX5v8Zulac6ZWS72w0w+SlCilFE
COwrYSdDbHK4mRB6Mv/n9bTSUuQ3lmnGCn1bbk35zasJB8M4/n8f6uOJCA/MNhAKAs/vVzoL2Nxe
FQWdI+zopgZaJNLgLCmMUq1d5IC4ES36ENc5c7gnDNeTFzk2F8Hr+6XznYSvdugAKY8KDV8TIfLC
uuOnMd6ooz9iY5mdpQVnQtGmHJuwqLWw85nuMcZqmVfe7F7k0aAL/Y+OtepcjDJFUa27RXzhlavJ
BKcsI6pJ8pwkGcK/nIrYRHJGoE/Cvg/nC0NzGc+5MmrMAuvUr+nFWYlf0a1k1ActMHz/pxDDDd3I
oI10jQh4jhRGch0mGjOkLbjGVKTw5dNLAgNxIOWKhz1SvjrDzn1adtGDrmwQi+CzeiPFTpx31H3p
ABVyxoeNunIvbExxJZc09nQqhibQUoJm6kUzWMd7YljwboyBixkwhgMmSdjw8+DYs/6DTlVpZ6Y4
K0oBsVQm8wOPj5IvscxzO5I1Kr+ZRS78MV+haVMncyL1jKbCBLCnVI/9wfEsNtrfQbmuzfy5psiO
L51JzVIH0nh5wofOpTh8ixHOz1fz9CJnQnM0HwzL/qS+5edo5CTAwvWNA6BXysGJlFmXXKnkjOq3
hShE1zymKURFXOoU0yPOopzcTGR9SSiqHH9EZToPi0T08GFpYhj/4ZZ3gx7NMP3LkVhl43wzg7fF
fXZ4HLWiMVp3kVAa0tybeieOrU7yWNhkn6mkqrh8WdKnuuIdgr8dG1IJY9eliwVyU8tYzfVFDAji
evJfqF4ShIPl3SqbTQBi4wV/wLvnznxF1kebLkad1w5eFecY0EZFfD+dk1X7qrWdfGNJcRFzibPV
wx65at997HlBEiKSFXthyLL+VkFkioYSVgFtC5ehSfa3NWcODCMgXIYUOH23VD0OZOvg/ZtQ01p7
ycv+DvUlYWWtUnX/lcIXb+2T1SeqlAzByw5LK+ZLZDNs0T91yeIcvUlCZtTGexH4hg35stjgG+ka
ZOQ5IdI1ekbsrzaBzZmY5CivO1sp1d4RVupCQQSYy1Vf3L+JJzgmwaR39Tf8ZE0OnZvgBJp0Yy0A
ATTvuZ5up2WUyzEAI6bZVQB8yv1hPf8wyD034PA+dyqCIWk8xBYHRRWgWJbKADinQbQvDEP8UKDQ
JDaaciz1j0S1QwHVpJtSBVe+61I7AsdSEYiX3MrjxNaCSkYRbiOfJWNq33gzv6HMqUVma9AL7rJ0
aFWN4E9YXNC7J418oGcOOKq+6vTiifeRgyevFhdMP2qudK2qnRVvJuo2I0hwjfRENzkj4M0UkHKK
ei/ksJ94ietmuJvHrwPUf0SbS+J66FHa6uyYbuPDZ5+SjNX7+6Ga+9G/W/etNPKmDiWnq8DGp1kJ
kz36LdB4gn7oIXZG2UEBByArrbgqqgMkq6YKWheAQshw7SLBrBFc1Xx5y/W0TOEt8PFRWeMNS1sq
VZg7pLNNtTjIIw7YFtpatJr5a8Z8qKZT/roIm6H8z9heyxaE7MS2LcSqNK0CAaAXah2K14/s7bpk
k9SLrYUJDlxzK+d/nMrwBH0bOn4yVCIqUCVQSYMvJr91BxYBF91XwGyiJmNl0PGVodp7S03LZlkp
QrkZsR7kuDV/lVK4FW/YQU6Prgbc6V8eJsgnHgKCgXr/ip9G3J4F2PaR39/ZGGOPWQnK5/yGyLx4
qglccgE6zN55/1xNHZ1wKDjtBF9PoHsQC/7j3jl4C7QY94LCQjhn+UgFv3B9iL4TJyUmUU+B5TKb
culSWincL55T6olU65zLZNy9xP/BRlx1C/S7QLs8TBQtbLIGIipaurmqVU+bf5VUwyESCto6W04X
MmoWFx9WzCF9W/YmonQ2RzBzyi7y5cWzKDx9b7UCvqygflopCrRVmDkM/o9KtEc0wgjyY6T+B8W2
GK+XdeTNed0FbTfaQqli9a1YVt2pk5sOqU+mmnUmTfuzLn1ZLHwgMCYwda53nMt6zNtVu1QZTG+u
M/Up5QdKyNJld/KnXfTBZPir3btjkHxA2YSO6bNd2b+pM9VNPcBDrjkDSxU6SWutlUWI/5sNBQta
l488hPLxQWVS0VGha7t6KfoSKIAPWVVJTTLUE5Gs7EsfDWkXtciMFN+UsfaAQJkfVvHbegtmjI0z
ct37AYezk56oZpolmGNRVFpUs8aa/RE2Wibn65M1nM+OS/Ez73JdNl6VrlAVNoGvHcuTxbsXTMa2
2v8gCOxChpjN5UMfSIUPq+d2XLbaPX24B+kft2PbRdAkeKYbFnBlAkAdW6TTZztkwEy0YLvb37Ub
sUQtDxH/QI6Grxm3wMI9en6VPdAg6GgCYqnUeBgNTxh3dEJFjyk/54cL0rvZXcaeTxk0WO3EQ7kQ
0Lm0ILVLWm/dN0sP/FGSJoyGCU4GeWE3AL/eBPnmVh74/PLKhkJDUknqnXIm48Mu9gujV2owlSSl
SyqEPaWHmt8zx772GaYQUK6KsCS3ro9MugnqJ+pf3ybLwvxSsgF0EMjReclzR7W00IYGbhFV051F
qyLBL8FzCJU5l0AM2dNVURJh+5sTZXIR+OzxeLSXKHFc8CbEz5b477ZXi1uSjqTbJc2a/xJE810o
wEP/LC5iGSljP3oNjdV1jwFZVPWXZ/Ob2s0TCM4el3X+WqXR1J5AF7oGAitOswUlDJXMQ+xjljX1
SdJXAX5Pr2lc5ps/zjqfSj4oUJVdJ7lhkPlbj1cw1yZZuvVljOLAe5POZu2b0vy1ZFR5ahDFWODH
NTbiqGJ2sIBwcnn2+6MAGSU4UxscTjrBfwwXO4xTRw63kKORVq9PZUQjMu7TARbsq9fgmcRsMwkL
TH0TNZ+WPBaxGATFrL0iyhPbmW2M/mC+ktiIAzV+9OFC1ZwAq0BRtJm10oGVW0D4Guc3ihfCgdMB
xqGo90JS5Ykt8/4Do+D9Q5KVrZhOs6SJMsoo8RLKBIAo+LimzLx5bU/rS2CYM8dAtwe+Caj3vHI0
n8Egm6cBGYe79tUZ9RoJQTjW92zETrI4aZaITOcG2KOpTVCdp/RuuBz/5l9XvXYRMjOJJ0xB5bc2
nBHbrsOOeg9uB8XBZ8C+Q1RCdfq1NLYyCPRRxWt4j6d9hTamw5j0srugaCtR56V937iH5xGRqK+c
ibihL/nGZyzD0b4unAnY33l57hO3mnM3K90PmYe0j42ghTwljTXXXQL+zeO3v4doXZudkuOTE1Hy
sGETDl01fPvJ+JwIz4XB8ZjyJ3RLqxi++NpMTkx8NT+XhqPXC9HemwEjbaF8ycVO7nc7TesDU4cZ
fT3kS71IjHawDD/hBsDmPS1CaD5+tqMP12F+Ac737FPRVaB3RCBE60L+uSAnZtuwp8H+pRY5Q5NK
nm/MKCmaqgzOzEtBdHc5A72kc3YFaDJnwpM+fNuI3bn/lNTswv1tVAAHbTYGLjdj6BirJoV6RQ2X
BpUTUBu7LtddexCbT28ETEmQFhYpKcF4M9Xs3CDJqaRDX1qXA8AZSj8g1I+vVJE7UT8dscnbuJI+
gl9XfeCSsydSXzAkZQ62qAr2ikueZNoeCDivyAUtAgIK6JFd0Q31h28kyNcBVsWU02oUaiKnqVJN
NowGzt4W4Xks0TAPMwx65/46gmktjMhVP317DD9o2DrN3a+mzEbvJFI09buFbWpPoCGmj+nNBwEg
OHFp+UNC/bHEU5JcBkNY0g0+K/9x5n09orU9J3KPhaL6a2gNYiDsRkh7CpF0FYtTvuEZnF/gUW4U
qgKlOi8rLORhkiYQg50dn4MlHZVmyeZ2ZYdXzMVleMb0hM1B6HLt3rOJ/PtGkjIfFR3Zh11+T8ju
S3vy4cM9cZeKWYirJfi68RhygwgU5A5tdKcNKdEqsi7NBI1JmEjWp4MuoAJPX3mUdviDCZAxe+A2
O5as17pzvxF7i7Qb2YUC+UUThc4gmtmmJV8Omdkwts6GbuIVd2j6/Ic28IOb3vW/WKK3qBvsj1VO
J/mXYllbJ9yX+eqk+/KIScW4WyhVXIRGsbIA1jC8AYPqoqAboDbJqrsiyucvvHub85uXz8TzGMJW
US0DJCJw5RsniBNQSk+4PXAV4VsbU1JNjyVaF0CJ5x4WPdEmI0TKGj7oOZ3saQlNTWoTIzHaXKxQ
QhHNDpw7cL7cclGw1WnnZ9kQ2ByEHriNWFo59xh5LyzLTL6rLBXVoxPBUP82UQqq4E3VbxtStcNn
JJJe79MgJF70RFDUhSX6FdEY5EpwS7vZ67JzKYAT2BBVY0fi8tjV/VkIiRQn7BaZr7zD2ddj6hGt
6EItgHgKsBI+OHFRKbnmENiGMkpi1vngJ3iyXIdQcm8BcAakwgL87j3loYu/pnTB6PpU9gjjmwi1
upzPMc0s0APY4NosvQmBL/my7tkLHlnOdRGo9c0/ifmhQ0VGL7TU5SCo1SSpqnWLH9CoT3gN7ggZ
yNqIs28QNFPnLMKP9BzCNb8ed7nHUc79Fw+fErDK6kzaSPP2C5JHbKL2Y3QqY+s1GUZPpITyc31b
e8wN5RWJuFnS+rm0shyjuu5PrURcBELSgzc0ZGQ93v7zDEftkKiXE7YGcElei9eswC6wbOS6P3jP
H7oPwpIicj9t/LRnm7WzoxMB6YQRoCpaA8ES7m06qusneVo2qBx0BspwOz4/45Uv7IuC2VmNTi5n
GoDO7xZbwkJ3to7L13IoT3Vc1Gb3Y0pGmntHHAWiedzlMYQzLbeejjKEYA5Wx0K2bq3CD1VZeU32
Hss/Sn0KoPka2tafyiN1bscAXWN4lYqiBHMJk2PFs4uBrwoREmee7xEde+LzoIKq3qVbRfH5IKuE
4Io5/iZgilA4/T4TxY/cZUTVDa4H+haVSc/7pmzm0wmEtGfBSOX7AvVbjmmbFEd5+uhxGRZqdKAc
UPfLy2+Al+Jpz1Z3JXlZMie+9TNZi64fCBYIHpGpBLqctplpj4HgsE27t1/dYBYD7LmXs9oEvSiv
8JXbDBWTGgr5f1J4CuDXjqMStgV2dr+suaV7f2acgSWrqBoT7In57b6QE55pGMn0py0VNbQ9IFBy
dlWG1RiigL+BehMsEh3Wgh7UDjGyuyOMnX1wmy7qQf4wrlD7CWAcm3xqYI5UT9qmZJrsAO3XFPEh
AQU6u8MyruEdKbOxjFsv6ASBVDxVPx4lndnOCOfIY1dvjaotrrmDhUAm7NF5P9lLJuKNtKmWL8rb
ATBD3Mzn3NhnHwn0ebTnFR7Fee3EpvmQAi9v81qgn6FRI4bTTweSNgnylKQ5hCNDMFiXELUt115C
FSSI6cfCaCxhBkcqesjol2Ogd8Kth3Kn0YSx1aa7MjpdtdJa5bm/C0a8jRomZXm5Jq+i8y4oUpVX
7rZ/H7oOe3XVuMJaZIK6em93373hD8Em5Mzr6ozvrDJS5tqaQ+vnMaL/G3A/o9TMYJuU3svz8yVl
Hl83z2iHi4yUU74rou+dKZTMgg8oCjVhZXDJ+DKEIFlHAAqmBEwioCPAMF3317+owlw63oH/48Mw
A6y8KMknRd9x4CriftedqQcNkafQmGAc+tC1Sxo7Dfo2EKTWOI7lHV4vhLFogQmZBBmoeTgsUqCN
mjf2tYDXvy7afnHMsVBkeElbTER68VDmdvpvNOGBh9+hx7TWEoJTE5h/JajhU6YO8lPUWW6fJoJJ
iAfkVpW9TpjOLy3/srhzOHzqlGWSME5qsSeGLtbZ7IYLNTTunL1AO0UvD1laMB2VJxA+Pv6olA9p
giuqgSlJcklDZ/uul0gu7KZTVdsqR3ywL8e+j6STMyL1awz12OKp6Ou0Jnlu9uDAQm2ff6ajP0Q3
xD220HRjuRPli9lbf3r7r8A7qxD2ssmDvdPH6vLJWMdGX9pePx2R+IY/zYMT7p2zCkG0lmUrtnhe
QOkIMpHoqyPuDhGoKC65mJPQ5YfHLRIA0spGjRiJVhRgEDIzSbBlvE6ohOz6jtmwG3KvskGH/Bml
1wWKGCLrrOS51IN2tOZOpnoneoih3u/HGooOAjFjZ/M3Ib3oSU6jUXSl82vCm4sNGkwuSVJsQL5M
2oOulRCEei34oeYvOpnQtF6DyBF9pxascu9/8cKHoba6BKYsvdgQij6s7TPhu0P920emhldBIvtl
sJlvPK6qDk9modzbt5XiY4c7pmorolHgFaRJsosZcV1OJjeotURELrpHHgQGm6yMnnvVq80lA8gK
gI6OWWXSDfAYeOmGPJgu6t6ZSDc75v4XlQdkOCiRODCn8IxRWuMuQb/srpSCpRmX0r+wFPAnttTG
OInnys6brmf0GpLopHO1T4s5Skc6SyUjuCXiodP02AoLNVOKZcZR1VOFLotNi4m/NwNoHCuw29JZ
YsehaCuNjXMpPJSyznfwkdmPu9aFTaH6iRhXPyFxr0vXTOV6lQ/TmoU9S/IgIqmch5xlVnixVISM
HykWcT68Bt5iEllCYm139Yso3AjTNn/tdY3U16weu6nKaNlkgmU3ggm+OgpBkEIzLraVdtm6wKyk
+Zangw9ZWOwvLr9FZu528O3j3fMPqJXwzyu/XjwLTc2GUPPkVoQNFsbtXrOUZWsQIvCdqH9CVvGW
kl6frZ+5HUurKr6TSrkgDc8DC6qy0xphinkF9pR4GF4ZpjI4AycaYWaPclNNZttDz/IRjObWyGOS
4F02gwwDlKC3dkOnkB+4KGzdRPHearcQ2tCGUX+RAVq1Y9LBtHVRP7LqiSSaXv8J1at36j15zsue
zBSBkj4Ies5o9sIJMM/AIgG0OEx1aVTZOc1loJ21l9qZkwSL70jCJdThCPeqOLwVuTPSoyM81Kri
x/3Sa2AEQWx36isXdQC+kA48qnF5w4RirzepeWzcCRN0Cm6N7G4VIWZMo4CqE61N5PzfbgZjjCnk
AYEDCIfxp8xl00C8w8X+zUtLCyg3gAL+6hbvqCQIyUscCNNY2SI7i4a6QcZVc9inQ3ejlshDVd4y
uhxDp9HFJ+ekpmxiZ9UQlxw3wEBrojIQ/I34u6F6WMlL9wFgkY0NxRyAI7SSULQxoZnl0qjgx5nz
Rdbz6ApVh7sX45mSPxdmcVhVERDAHLIpYPzuR35w5q5j8lF26sMNUAhJRvO3NP2CaHul+4y1V5ow
Y6H4GzZqRiJJ+aRlR+qOS5ImS6r7u6x/RYZwE2WMYferG8FgXWH0IUUx/Wv5QLHvMsPBjZ63TYMe
w+hZn+6c+gf9TPiVEAh0H0RRaPWeyKNep3hJ/F5PAjKmvZDA7qY23Oyahd34R2eXSawWFB3Wanxu
ide8AbqjlTai3zhIHLm2S33CHiqZvZKwIP9a0UeHH0cGh39Bh8eaazc+LAubIaKMRn8cw1Uh/E2T
+0lCffC9xglJd43Og4iRrr+HkLtrZcUXm99ziKMTkYjQ5FzEKwat7mquCRA5dqTtoXN+ws0Qs2X5
Twjrq6H7HmXzL2ejhYZlpJA/F0CaAZMDgikVm35i4D/iWAtK0cycJaBPE3N9N6mJc7/penCiIk7v
f6FttR2sTBU9QUV6VKzTxTZ/uLvQCMnr44gEvvP9UiupHDbl+qIreEJil8Zo61MVp9JD9wg40Rw/
xuUgIPvY/8VEwphd2WeVGSFkbQGm+bvFxqNEnYu9X3M/5St7dKzUQboGmhbxgfsYrf2Z/6OzC2HG
PDNQoQFIPOfpbh7pb7UBue2Qp3+shhDa9P8YFPiWDBiVMzgDWq8aJAy57Leb+2CnjEsc2ikaxXqY
uDuXtvq02DqMoSq7NcBfYU+IYdKlsu0TTeow37S4Ia+QoXyrVg00uS4LD/utRKj9912yk52YJY2b
7+jLqeI1F67UMCDhC0GM8JSy3RbGbqnz4A2rYtbVqoNmqP7EdJYwcL6c0Cq1MEmah9MxGZxEOcYE
x8Ngacqip5oIZSeWr5o+nqqKejHEYt5jUdOdsSmeKx8eQekUwvaajRjIiMjlD/EU4ZZ4i3FhPLh0
Hl9Q4nHjp3FNwnEJAcUfImffwwRIMQWufjmKiC/q/uaYoT485tlj884sgaST2B/BeY8CU3VZJh2W
/FA7ZbFjkdY9BzLHTFmsTLJSHnxnu0GmV+wbZLM1/xSVKvZcFKpjphSprtf483qV+SzHtQw+AeYr
6DGYZ6RgTmhR7me3qbeARAVVrKF8wnn5Cgb/wbcCDxXEFqjBt1VynCAKoRU9EfJbWjR0kKICOo9z
/fO9h8I4u2SpICEuhugW4ntDsD+ZZuMNV2tgBBTn5DjgtMJMQy7d46I3wV1pMkMVSguPsC7eqNh3
EhdxC3yToNEzss8RLyH4c+yX1DB8KtgMtZrrYgzyBZvEg/0K5ck2C9emg2yCLYFL+Jl/wjlDR6X2
jp2QB2l1xCi7sXoNUDJTFUlSNsSwnFXFNsC2ZRL5sXGL0DskTkb07WgxEsXp0oUbU2r2QZ2rHYWe
3iIi2eRj5pZ7+O1SBb5XErfTuTCGrTbnaO8eUvgpZyAT3bXn6VbbVHDazAzKRaMDtChuNqH60gPq
wwzDu34WsdTfxoLklC06R+7KFgKYeyAA0YGJaEDpZX4QhKZJAgZcWMtBFfOuWE/IelCUDL0MGR1E
Q2rGFO+vbQiJ4sCDfkiwqYjUi/sU+qXZLUKk4gXtgBuDOS7irpqttN4KjzFnfaWvFxsEG9SQNpLE
Wso9qkpiAYSOpg1yZ/jqw2u3mVMtYQJQt5gn0yDv212QQAaxz/wGOec96CJ9hrqvUyoKrMOm5B0L
/RT6c1JgMzlttsVrmEWyd4GwUkiDRJH4pcfc4snrwWhG6LaV6c0qAt8KLb+QaoXjFGVLYPjut0cY
snGxy//v4HDOcyaXJz9faBMbW0SmRr8uHNC+k9mr/NrYMsegPVG83qkHjf4pa+pRcOefIw/Cg028
Nlf9hiHP7poC2KK6E+mYybkYXxBln1qQfM8uCizgQDTZ9lm/7IOslgAbOeO+5g+HBUGIIgW33ToX
wsJyC/bKrAa1g3Na8uQeYVvJHRAi8pfoZWdGcm2ZIWG1fSys5i1usIRepDV92mWD7srAT2iuOlBt
5PXA5OSaBJUvLFvlhygrrfUztZUXlc0Hh3OPNy7GBdRxrYvB0nO2B+QSsfFhQYp1I7isOkkHt3Ld
3SMXjaEXwo0ROVYLS/FQzCD2cBUE6CuxPp2p5vbJuRS6i/b5gtW6YUEK9dJLqXyPjfRIHbwNMHNQ
j3D0aWjeD/VmFDxeYyBo8IkvMVsXRw+lvoW/qF1Xtr1xhHGOzIHgQEICVh4SwARWMlGMrg6wtMT1
feayCam0nLC3KpJTeIOMQWmSCfqSUb5TLUipK0c53tBNYx7ypY3rs32IdkUNxiP8eBz8Or05Mvxc
JxDHFdaFch/9HhAcM7q5hFeqKBuVDn23Vq2/JM8LdmOnJqQfmx0M69d+Mp6uhmGL8KkFtFqXJQ51
z6uTH7jTAq5sz60HL8abcUYDbJVDHjU5+Ba2Z85hMuoYHR150fRq7MYUY4oP/jIs/pT3A89qL2Ds
pjoUiQvo1rYUAJ4f2/jbm5buGtehQUhKdF3n/nKRs/n/vrJrZ9HNbszbh4yFsEPw0yOGu4IN97N4
mtHbormuuHkg3D0dscVYjNXd2yiyd3qjOi3cJ3sfE4Te1//aBxtxu3L72RvjiGAB1qcZvdAo8Fe8
f2rIQHJgB+pOdyb86Fu9chrsZlNERvL2l77PvZbLHg8R763vlIBwxDsOOo/+BaL9/3SybXiA+Jk5
CUVF5tqLLaiTPX88GIGOlH78mJC5hGQhj77I2pzKl5AZhve2dOt0thc1DbTDvPaSNg1PtHzEOqGD
RVCd/f3WG7Lbvkd/6AWDYFRlXOf7ahKOZp8Y4t+HkM/kr6R+/HNquuIyPjhiTsvP+s9+NxzLrgcZ
4tkKXgE2NqwUtSqD3NCtnp4fOM3GlPLUcHNThq2VSjc8Ncrlq2SfNatM8haKDwvRwqyXFu1bfApg
eF3JkyiEFYUQ5HaUyON55kuCSaaIBO+cT9q8PRJUa26Hc6v6jmf0bQXcYqB1q0AKmQqfqeTe3UqW
m+UbofVssKhaAxszHLhslcDzAcx4WbYgYvg7nQpp6HCecQQOnROpLGiAw7uAcMao5/RVVU7ZfNgM
scw9pZxj9LY60PdvndD/N+Bhn67oRIWAyYi1IgxSFP3aR9Z8fYFu87jiSf9/B9CMOZaQyPHy41WO
AwkgIYuRakf8peOh296cJSqiAoLf/nHCK1F9rqRc7I4JYuMcHYKE8/mcZO0hTfLr6RLLVECdSxoK
0v3hNVJzboYce0hv+1+U3hoTzv57/LXDpWgEnf3E9Cob0o75pHnE8nW35qFMfJevk4AWb3v7Ii+l
dxTxxCW1wvTn0+rNsnbshK+VXY/2aDg777QjFFRFeUmgxKOlHNaIwLi8Nz+TQD18ONqKlhUmCZDV
TOdvP5lW3GyFUi1kCNN+HjSIJgAvd2FIRme/W+IYYBMvTOeJFsafxIeZU20ZeA3i6OxkipXDYG5R
hKh2mbB4Cysoyu7eLUaBbRRbC2oGOeqB415yOOLxon15xYGqpQUoOCfZQPEtnjGe+/5sS6VxMtVZ
gzt+xCYbsr8gPqo235vYCW++jgoHWViSXyszoWtNDmMv3MPhOXInHTB5VYh1pnqSQay2mdpquKmR
6g9VzSto42Oqs7yUGd3MWlxisTogwSRfHtI2EjzjiyTOPLWNaLnqSSQBKG8Jf3kXDx+MqEuoiq/J
lQET1jk2NsLpbBdvTIKFtTVsiPlgz4LSXjoU/lLv5gIPtsm8iugvIp0ZAb8TBY6d275cU8/fSzDy
BIrGD0yuiIA+8XEBp2roHCNT3kePWBT74NqzSvp8m0rE2wzEW62CtTesyRpZSJFs1+L2+TUZVm/e
eO2MeJIMU6geNgE+5WEr/01UcXPN+gokZmOaVVH4gWLu1r29B/+aPLYWb9awHhM2S0KOxpxmp1N2
3/JK9qq0Mj0xU1roLwhUwk7Larj9lSd9KCT/p76xJYOcrrsjXf6pMFGTna/swTF+3zOpFxWqwm2u
OI87qLlpt5kKG5j8r5HF9locCbzvjp8aiDeqEEYpAWsPohMEIPpt1tsXLmd4CSYvJGXHnWQmIyEE
WlNDScx5GGUd7WZZ8am0B+UHO+MJVYdRRy6yZxGw9XuktixAydwCMRS2k5+fyi2ua1MWhrDTqMw3
6OFFetFFvZuvYzICK4rCTEBA8ctnHMYe0HMt+tq1rCoODFeHGBHPqY0nlg7USwSBZN2mc4bMjCET
oh2cZC5U6HOF+jyAsmiPIrrrI3HqCxaYtpkHB1A6GOB8tLmBpTiEbO9LXHEzfTWVWpegJ+Oj58CZ
jseMD5VSvPcjHkEAmkntlOrDHSx0VmIMwnm1bO3EIrShsEQDSV925n3jP2fXriL8VwhGfiYm3QX4
odaBArpKnLqvzHbWU9Ggh8jdsZpOX965mfdJBkVmiJNfwETDYV4V1VLz5tcdy6KJABjRjRL5AfRI
Vc7u3r0cdi4iAxU03OnpAZpSnxnrqinRWeYJUJn/BoJNO4t0+Tdw2QAcF+whgnitiR0ZytkBA4Sr
rRN7cQzvp5IC5YKacaA5G3Qnf4PCQpLXCx9ZNkRUyacu5l7XvoidPOwU8EpoYH3qq7IPFgqMQIxe
4O6mBE038FTNkuexokn1vskyuiATUsRksdgDLSVro9Je2o8L0J6UH2D+z7K1O10A++AYHzCmh2UX
1K3kSmon509GUVfBBXIWYP2noi5maeLL4oNZFlFDSicN5Yb5sEuss+0Qdu7A4FI99IRVdeOYzTA7
gF2e4rtEnnMs3NYewKnKkvClcoCCTCW/fglKmBLYAjbzdbo8d/kD3Sw3cSWCPYNnM0PoyOHav4MB
5LIESvYUjbT51db+Qfq28H4+k+bS9BWSMM8hlg+z4QavF658WUNCl7ZaKwC1XOnWwyA1SDK6vRXX
b40YgNAFPVUOMhzDu08+mzYCxlAKcfWYn2BWriNPEwldqk9VE1/XO7FBbeHWlnf8vlZNIBlc6uPh
IpPwUDJqhCEKSGuwQyhzvC0eevnqoTeVvLY/OsoE/ZL/oGPhMS7HmgG/0+QgYha1N8sOoN21lYZP
7156XFV6L3pZpLbRSLXpb2mpe0jhO89h1p/8RSG7tdNDRlrRnV1bf+vRRjS2gbKEaPChFglCJBie
68jZNR2ZB4HKALiR5D89CD+m1Y72IhXjwrmCZoMQ4TTpAvBTKF0JfADGzeKbIsoJoLPPJpbg8VvR
+k8N8QexXs+2PD23hApfgcuYrKR/B69uKwpK+0e3nJwwMUUiEJiqZn6bsvPn5sup1XCuVUK/N/vJ
Xld9ZSnvowsa5ZvnQ1l8Iiqqv/0qoedPvsFbXwvehE+mDBpciJ53ZqXAabiiOgrBWTx0yQG6YDr2
Jwm2ucC9b+zKf7SkjGH4xgDqPDS80l1ngRQR/168jNZ+OTSjHPVGVXpZG9iIPdAGnCDCanRWgWzU
U1RToyVDUZz+XDQQy5eaDn1FTtcsmXDRavdf1CXDXTtqDXYXD+iWgEazpBsR/nG56wzXzh12oGc7
g9wHuC205yRx5SQyICORL8Al0tIqvZtVeXZyXwZlQAWeAGjkR7eD/jeL151XGYTB8AV4QCfDW2lp
NPg8tHRDCZJUb207AKBK8gkPrhC7vOGASVdWQHliLJpB5bHCIjMZgxyUr0cfrYo7Kl4FWaSE4uNO
vqTpTfrRfSPoPIDvNnKBml/9Ss+uyjACk0xdl30NjWdnrFDSdp0QDUZ7cNzX2EArRJr3r2N+2p/u
zRR9t84c3D/NCJUq7RPHZR2BbK8zUGybd6FTN+wjJDl+J7y88NWo/W7prH0tBsXEIm46mh1QrF9b
D5jb5FyNKET8hYU7EPLpV0WrRfja4RBEYC3aIuuUENX5R26S4dOAdjdcOjkeFav8DrXmgTGkzU1R
yLpIReoj73tV9eGD+9TO1yn3mfGMkF0qhZ8XA9nDp+hUrtfT6dwvd5uwT2NZ2PQ7TR5Di+D9MDwf
jNIqzXMzjQ9LU2p0oKuQEKXku2nFO7/l2Plv84wVPxbIQmi6Q8OplQgiA6VzRM+ZZyrgH0Ze6yJ+
cH1PNQZ+0pF5i1DMXKqfKzo/GFWq4bhWXscHlW36wjJu7Gsc5y0u9HVauhQxfuiBD2V8U2bJZgkO
H4zcU3sN+PcjNGq1emk8btB6b0Di6x1/arkEDCXB3X0lHsjTziChsJG1Jyy3jxF/9cN9rjfHmFxF
ZEorv3N/8sdN+B7fyrx6uTR26Gt7aBYgGiocIZrn0Qo0037zvPPHSGCvvijSqwVFcqFqVMsDAF+j
NqlPrGgGmin9eppO7QQWXN1AWal1svDQfCRScYUiEpcsVbxTgb13vmCyOBPoPN6lNDm48lFqtE4i
8TgofZ3CrGGCcBnt9y/PJpBsXrMa4qum54nr/zkp2Lz4yRD8naa+ab6dZFaYebv9pks3KsBiV9j8
Ln6B8NmhhBi82GmR5//Jj2HXnMr+AkijiwNxQo3jEDK8sYG4SF2TOzUJPQ/tGi9HS4vlGtgxUulI
J56aivvNidD/gQ64jg9Wn8VMfYJfVUM3K+U+FBHZCM5o7SBmpyVvf2iZIiCXv8WYaOCRMi9Zz0Y3
pkGIAvYXkbZuqEIhxc8FUZ9zTCm2rocnrjrVRa9IIbj2REZ67mrsLQw+9yaqJxKMbg4VXq+qJtI3
4506PsiYcThZeCgf/Zt2P86KiKROE0aARHSbBXwrtjejrsxYcayd9ObIvSN2CSNDFJdeTigdMZHm
lPrTaezD+ZdtP1D3K8uthwOW0sKg1EKdUle6aGQcHS/znhc4qEOtaFMFE302bZsaPHsq+SHt6LEg
YS7t3TIxmHw8y9vxuHDd0BnRBv82mO2BVgUG3HDk504LjJm5DIYcJ8ytQzCxrDizzeLFroi/0vr8
LXRvCj79a6zzlNaBqe795lGSinAXyqOenliqW2cDcSrf5+a7+QoUcpEics6YW1yq/23nqK2r9c2E
wEhn6ndFxlTVoeUtAMr5sTL96hLLs+40tIHgZgG1rYhSagi6vrPaoxv1TZJ/Yy9fJRti7yRTo2ZI
TngrKgEf8fdxeFZZ68RjvUyfny1Ai4X+Mca/qlngyGVRbUAHPPiqUjInB+IEteK41Vbipimni6L1
zRFh3vTcw+N61TRyhHfjbgNnxSb1PRFKe4Lk/lgnBQqIntLqYLyyx9a578o/IEG9nEfxXnkJdTpP
k1ge3aYiGsMyopjcn4r35DT8fqZQ1Fh1p4PPycoCdsgDcMc6weXlq2J9dsWTow4aj0vXPnvVNT2c
c38iIcMdsd43ELmpWZa7COKrjdTx9zlXBVTTHLNBmlHw+e84Qwjf5mVExDx0dNGxFma1g9bgcvkV
T2fNEOD5l3vWpox8Ytqk+yCfMVbYfZdyCkIuFhpPeZUD3n44hI8GbUp716BMNrEmpsiHiflttE5U
i4ftSe5EnGK6KnGqLrM11SbUoaV+d9ijr1Ad1vRbzOHucLE+MhRAKS6i8wGR6B2L3KQaUZ2+DKdm
Qn3S+E9L5LghLXD0AzhvC5slnjXhTnDxBm6gbd+RrEY99jQy4nI4VNFoV2mLHD5iPn4jGC7C0i4m
1z0e+IrYfKQ9vvcff/LEheAiVKJGxejd5+Vi07woWwZJ7mP6vX711QdcAmSwTF8dOEANyLJmJ5Z6
CQPrZmHs192tSCW+oUmS+ngnDQQ2nYsuG3lxQ+64B9eXceJhSJW5kMeA3wxVkKoys3lixP1U0dgw
gRtX2g/y1YbMhmxokuZS93f4s0biStthk092rwef47mg3M2LCcM3FdhLY4wpPUAgvckM/M/Td7wk
VWf5CtcvMxnhY8xETbqCljUc+i/593T3VgTl57XOykGVuXgFX73KQVQz54UkwHpnAM9Lrt8wSmSK
sAPh107loowQ13+CGUjhtykRUsDPfLurXQcRMjv5v7osZEz74Z8xItnGdW/nHbDAd+ljsRQPXro5
r1GehdnmDc0kAntShUd135fxlyqHg8HasRmALP6nyGo3Zs/mIQfOGL1m1TUG1PBdoBeu/BCtKAL3
u1hQ5CgsS1cFGm8XUB1qjzl8iw+yJFvh7vRNZ9RzM+b73N5HjHxDOh86wrTGhWAV86riue5upWl8
0/742pdYf7xU7cfdGvUrFJD/oKZ38CYbT2tQysXyk8Jd2MmElZqaI/dJ8d7/HK2Lx6JGCZYVnSKY
kgbZl09eUk7ofBTpNWQTK6C+RYQqvZGdKY16sC8wJDjyJmc7ryTtIXkNi7JfF3pWX5VI3MZrqX0a
59aQsysGij7abXaAkbZzHIlCu8ErmEiGLy8+u3j0vFQdSmFhzeVNz78HcZ0EDuKTL9RjlxECZRLy
GOJUU8K67UNI0p1m2ibSU8unEQZD0pVqRfMB/02M2619SHBCgDy2MNE/MnnRGDHOsiwLzrpvikq9
EO28lUZ3PYMAoyoP5jE+wWMiXYOW3qiU203uJkOFDibYHA8CGsf//Yc+WLVZz5CgU6/2B+Y+rHgB
YTbvA2Pl8oElNrT8QLAXrwo1pfQXijvEPwMWISizVX70TxOYsb/R0SnJhHGB3yS/KTQpd2uoBL+F
+UIQQEpRRspGVNrmFuG/O3QZPk6ZDnC02gUzJP8nlzjc0rKvkS+fuba0rNbGJm1BWwcRg/hqOs7M
rjwLt2SIt6wW7OxsW1i3pyg2yDYFIK6KPaAv4Qmi4KjUHc7OVN72wsyOhuGzEpkTuz5s8SsruTpQ
Xpgxpqa8qNkLPwOj/WffGYw25uHHuvfqXjl5VnU8wNKfgvS5UCorWsx1HfAqFB2JnO8LrULvuAEY
cECI+LcQ1ofjZD1A7FUm9BGdKwg+WeeAKU/sUU1dqHhYwY0i6Jfkn/29HwJnuXflIsBN6mbRmSzd
9pYmy1EjyJ3YHu+QoFjhTncG8RYYK7MjJuO1eCKcBDMHuazDgHmvoXTXcFMKb7t2N9TalHEaBNfY
VIezwN11M1zwhtgoyVy6ejab2yZhNHu9FXXD46VbnswD0jLodduIISCKZ9ZRqK0KUHlnH18axCFM
GsK8dVsPd7DQJtnCNPlZjvSeFvY1hmS2iwzcUkpMixmSJMobewbrPO4b0lA4nAKx9mXOrfseoEpq
0aneWRRaI9wMV1uZRD+MywDKUA9UJCbhTKPWMnrqKDIzGixRJnqOmvm/tuWT4RNVSsw35nu8rxLa
DoqDBybcrXL9PKlNdFVBynj0whIiYkkthRyeSZ83ik8qMxu4KwGahpOImWpjbNSAoz2dZUc9smk8
c3w+8Q5Cul/dyhLHAu/vIV8hPqPM2aP+R2dkRtvkCcYYDQE4B7wn0M3l8AOP5scy2afcT8tUqRPO
qNmNEf8hd6ehJtESMIrI4dqAh9wVvM5NOW3ehJrIvwlznEpQvw59tyjg1ozDHD4c5bDcYmBZPpC5
OuQZ3nakDzzHk1R4W6sYNG6Z7P1ONoEX6LxnXO6Q7qxqPmweHg+EPOBnifD2s4haeeqah/kjtJfc
JAYS8SqF7SHaSpkTdTj6Zh39FyMY8zXah3sf5ocNkjdc5YXD+0ts5q6EONg/hydIKobH+5lf7cia
RptnXP2LVRN6WXnqjMM1LQOQBd1HTKvVkyofyCB4YVof5/cRR1alUK1ybIdiazyREUrp2DWsTOei
UfR/Cx/k/R87H7D5djIWaF5zAjdJWAdOOyrlfopFkHyHvywZ5nuO+7emSexf2t0QDA9oy7WIn8sp
N4gL3htIrCg/yD4g2Md1dopWZeUojzLT3WkLPl7ry93FyBMXdYeJw7ywmgSQgKpjZ2PX0dwZNJzw
M8pozOB1KCB+g2xgET8+3H2tzeZme0icSn9o1r/JwkTah/uAP/ItUtfYdjQDF3Ne4y8N8yxc4irI
a/i3uqs8X/W+wKoXn7r1cip/exZthOtRb1/rYnGWjjAElQv//nuEhSze8/l8qWGx4w7c8hjOla/M
/wEPUQFSVN7uynHcre6CsINh+Z/jfC50BwX1hFQ8+QAMcz0UUhB2TKDg37VH2Hrqdzd5Ts7ZIkhh
6+yVemjM0HX3lQm3iwAZuLMk7vNSsYTcQpufmnTPC2PGv6xHremXQo/YFxXrwnyujMDKUiOBjS+k
ztt4wSGc1HB3Afi0HK8TwzXHUMGN/0f42RcZ4uAy7s6091XIgAfGUDiXCevmT0G5V5zzdJOCNbNo
jShEaPljHdl0Q7D94l79fuY8JlDAclXy9o9LtsmB4TqxtcN+CALVs5Hirryd09NQ4luJmCSDcD6N
mq6FOqz20dZROUi3nscX2pL9Fu6gkEz+pq0pLssBfWW83xxRqy+Xd6IOf+Y6szD6Do1wFlvQ0Njx
3u/UHwGpJjA1CAA8SSxVpViOrfHfu1aKg9ILs3nMC7s3p7t1WMMmidsLmmugn5PGySrwWMVvJqKH
IsIPdrhaKUCM+NVbXPc43o3MBx0+QsszUP10westZZQLI5M490h2wyKqCjxpbaMHJLWuP1VDGIPr
HEryo+H6vhTcV31bMn46rHM4oonRTIt539nwyAqzRR56bcAl0BWpZ+QIO1MJQltCpHEUedYGAoyp
8KnWPD+cLsiDOeq2m/xkgJpE27HhzdVKCY2v6nBsUey7PZorP3AfUXBYasZ44GIJCTAo0TckUt3b
52x5xHuMg1iWak9JCh0IX6HfpH9JU/ZXwil+kK1cqeWg+8y7S/svDe1JgQZFy8k4IPIhSzTPESvm
1yUMOswhE38u23FLpKMcI4k3nzAra0juc9bqmxKEAm5tKSkuG0DvPQ2oLp9LMCA3tNuSauaPcRpd
kTVb+Et8tzs6EAY1aWVe5M9L6BTcBdgevmvmP/11VEF307Yz2Sk+7Gewhil8LAJQ/9uj/QPTINDu
+NsqPGtaQ4KuCgdJt8XgwHgbsaS9DKTdHLf+ARP/F+SVyQxhFZO4oZaqzWNqurJGGoPPL2Kxnine
85ydWkvzkqLTwkyTHskvByMiz4rC6w0mjWVMMnwdSPaWILas3GtYCebI1mh0DCKSrnTtClwi9K6B
J8lQxqoeBzyKg5d56fslfYoCB8zjVm3ALXjPTixRQgyDcwH4uha/FMd+p5VcdOFACnGGevKWEUPr
nRYCtaNOo7UQptwaoI1S0k9TJAhfZNt5FW6yndy2CXjWNSM4nf9AO69HS0pVmcT8yxyR1MZIBjRs
X9dIz6fYp5nKLKvTmwh2cQAfkuNTD9jmLED/7DJ1W19i/lH3JWFsQLWy3cqzIy0X39eUYVkN7yUi
vity1Z3b+K88Sj2lMn9Hz1aBI1wC/cRVpMtr+Wr0c0f36xj4cR3chDUxz9AH7CfAy89IuZ5ghLlb
Py2H3c8CcFxfcPlp0FzNfPZbp/0ANfUiTgNz7VvN6+o4nGLz2D7zuq7EoFoYYnUqgCXa5I/hToc4
joVy5qhWNi2uyT8qiQXoHye12HUFr6yK+/M5VbQ17OFzWsdAGmL8B53gEaakjQWsf3j9UHybovoc
0j8a+av9GFjC7mseRBAMsX44zHRwFqpQvQcHv1YC88mZlQSKLpfU4AoOIli4VLxIKLWyg4p7ByhH
PYsvZp1+IpebDH1QKrCZOu7Eu//wbXtjuKtOUA4BxXz9QBqtlNeJ/rMoIQhhWarZdNCCDSO9olQj
MGJuk16x4BmJp7EmRrbdCZXpU0xUppNpxZ4o5/6FEodkmYYcFfpasBfXn5vN0IFx7qJypvSomCjK
IJRcgJDdXf+zMt6tc60wVIEIZTTdENEkXGYb5r9369dyTfXvOFRR9NCZUG3RUYuUNwzlCyhk/Jec
Fp2MnZ/GgZDp5iKOwWl7RvG4Y9pmUTobwBJAmVqmERPlgi68GrJVnXJa0vGsMn3KpVz4KFoeew2N
kmRxi7Cz4FlCRCiil3n2kVUG7KZxBd8KeC8PbOm03Rf0ujg+1FZRMAcnalg2AUr4qc3UOUhFAtSN
rmd1nCZP9jJmMU82yiebimBOLLWJ4VsrXFk7xCeSNxurNEu/gdUgtBhoyIe7GspqsJR/DXpaaYN7
plEIPha36L/OCB2lGpml65hs/XOxs6K3ZWDxAaN21wgamtxjsKY7/D3jz81jj/iozNpCa+HQuxGf
g3OnRFjF34CrS8VgyGbVoSdT1lWWdkOCCcXZWVdyA1v6+E87XHOZgV+7Ti7ZtTb8y1SI+HZs0fX7
bFNJgG5YmDRh+jDQxWGtlS1vMerfFYRHM6Q9JyFob1kvf2tJzW6TMg388w2MISDdYSBRgxoX/CM2
o+V1adZH5F85Feou0dJqVWyrCbnR9IeMuhkmpRM6btGnyumxug48zCgDDoKvqgWtQ1oojNvgVWIi
FOa2nOK7TFNcQcDOw9KlwPxNV+Wzgh0xm/Y+FLYIncx7uRPjcEP+uJFXe8q5foabF2SnY0ObGuLP
0EN/DWMhMNF/ZRdguiNcCkliCFETFyP4kO3vIFOuwIvoX0N+4MUZibT1ns+QZ6Ei36Ny5cqfQoW4
UH1Zey0/2HpCVcBkBm+3QAQleFJtzvLlBrNl8fA8t3HRgmR4rDbJl/KLTFRlZHj83KF0dz/DDkdU
GsJdopqvRNbnQGDmu+rMpNwUEAPO7ekcMUMz+cfsGzie9P/a6V4LQNYveSWEHPM1O1qrUlf2sOQF
pPhAfGF9FKz4OTtglNideukrZvPB5D1cQNSqm3vA9yt/2yuUom96n73Kpzp3XTvPtbbphjQdLG0d
SmfymuHRU8wMBWS+/qXtuPLnqVyKrbxo1ro6pDNKkhJ4Gisc6hO8RxZtNYKXI8cyM6fZ1QoPn9JH
SkfnndMN/Ot30xT2oVXFGhtsCVSjioQsV0Vpt+ltmj5TxYB8Cci113mJG0lCfL8wTJXFdtCSZF4v
UJAjRgow3cgRjK85WA7M0LKMZ1crQeS26Yyg7unB1jeS9h6xjOy/t3x8mrQkVsw4cXbIddFUc80Q
Sc+A+WuKxBoeNP1KJKfnbEERhvdFZt3atbCgy/l/AVny+DLrJ6XBWZGsfReiBEUl7CiH6YwNNL7m
SuRzhEQ6SwGbWpl9WIvfwOAgY7xfLDQsKBsuD7AISGWvWj9cLwNVhq0uWADQVRIS5plN+QRXpr7r
SbwgAaqy2gj2wOpfaVpHAeQwVweJkas01OrOqBMqjJSzvLksX+gQjpLaj/mbnTUzLx+RcdecYELr
bxEHEAFxWUDsO+LwSIL6ttmO6/lVe429/MAopOAENzV1BKUzKKV7ZCrbDC/nGIwBC3OCBvvvIpiH
cEON+/ELlJpcrzYbJ2JYz2c0MxseZnVrZflQZC4Hw3rmC6HH9Od2lNWJUhRBxYXArYljhyinrqpf
JDbnFCk0cki9VJsWVIJmX9XTlGcPmEVE9dAWrwTRSwj/P9JfIr8QZDs3U5lx6FnXUb6+sG4GkoEn
IdwfaSUQNvykxqP4fFQ8peyIrlLlOXiHTKOKS5tR2lQ/CnuLLklScfxIFkbwYPe0RkjnH8phIFE3
ae8ESyKpBG1lTC5VfknyLZQJ6f2lzlW/CCEC+DUMwF0PyidRe6tXIbgSoTwrd/aNt25PFIAeg3tp
o1NFPKnqIETgAPd5eq+iw+YTcgUBr0rwiaNTmMu68mYlcYf+wdSx9vxLzZCx/4CY+qJMeCsx+FX2
CGf9VWJlgrOAKB4SCb0qs453rNsJ3rLw0FF8kbxmBBPqOsn46vIIfMKB+jLGdfKu4+0dOvRSK3yL
791+zb5Sys9uvpsLA+FWq50g9ppeEESngPCVsDc8Oz10S/SYh4vCJaqMVmDP2h1YkrBo4c3uzu2i
/t3r3bfpv6gGccrz0BUNQrDRerSLoiiOU0i+H8njU8rRr+LUIrr5HA6etqv9c7Q8Oh74zFCOII13
OfsVtoaSjgeY2aan9ipS7x+5a7BM4lmT8CyBA5H0iXxgtUy0G6Wnweqm2gWqv6pV7JGaXCH+jMsx
0krGup4XLaKpbgwns3zs5ODOCQq/jKeq1S4NZHfuw6IKunIjfGiNy9+IdnHAx7bWULksFlUTzz57
NiEM8e8IYaGDQG1Q5SamspHsQtHoy5lPdk0Y6h0eReRt4ygFFlXRXleFIo0ms2OAzEp1tU6OTk40
187TLDaP5GeWkZrqOlkZYUkZToznC1A9h3/m1AZrfRFeDaLt1rTiHzo9PvAVjcN7Wze6jCuSHTrF
FzoKzt9C7GVQ2WZErtNCi+fuvV59ShWTmiZKELa5oVI53ivhH722NSYgwskfOCPz/6dyi1yDo0a7
XrhBHD0U2Sq9R6TLt13OVH1ZCk0PuflE4IZn6vGCoJx68hk3NK5oJGA9HGCPmdSWpjO9gDuBLXnv
hGDQm9cZ7fadzs+RM3QvfWZfQBZCMnxS5/uyVd3Bihelv+4QMgqeh6wJaJU000fr1IxaN6TW/+/S
RUwfAlso2tSBf6KwOlOfpeJpncdia0gSh6yhflk3Y7IQ1w1Tf5d68+Qhu9qi7b24ODkxlXgueO5b
WX2xqAPIIDYI718cR0aKRj1oVXsJDHeG20z4pyvgS2+VLKFasncqc1UAcc4Oo42Zg8uWPzm0f685
ahDZ2WtPThD/Ehai8z7IqKl0z1q93EnG5aqyVJgKXlhwwZpalVFdwYUKD+ArLP96Nd/q9MVOCpTo
fX8Yt0X0AktOvVKd7eBC4Woc2dhWh7KxVc9FsF/vDax40NtDMroyZyL+6a/ZVSbPatWULabce92I
krC92pUOGNZYTLpEPA5RXhT61lUJsHE0ZUa00Xp/h33GnF1Xw/LPwLE6Rx+3WrVY49Sd+ooUCeYQ
Vz6HFfLxUe4md/LMpf1tU324k2qj35+7WYa0cVuXFk+f3WCSSazhSwS21ZkdHNxlTUNG2RNBjkgC
4QIGZ0hsO60cvZopp2LPvDL1KaMYFJaK3NQPLqPJp9ghifzTgkPFeZwNwl76ZXpEv7O7wbAg4Ddp
5daOIsHwh/4aQx5ajJgqG95p9bIg1E957pkD93/bSYjBiase3xckeVELL6iu9PUwRXiX7usHUf0/
L0p0TUlJZdYVrMfQkzIb0KOGSGDzhR3UjG8W4PNyb1iGLArfPzxdro2C4MtSgTHxpVROxqVN6YVN
FvkMYJrmm+FYoJ+q2mZvB5qgcvtrUIRRuHm9NVX846x3qcCNJsBgtzm4oqA4+iZXImwFlzsQfxhe
uJDSAGyFcSyY0vRW1olBqhW5hbuTuF9k5OBH5wzwHnm2Hg3HXsyJqmzrS7k9+KJjIE4CdXy6M4rW
AtNHZUsmdbV+CdtgZl9IRd2e0HJITewU30rNzpV+099Nl//hQd58qEsBw26ru40j9rXiBiuUXM9M
LHOBfS9fIBIn0X1SsYfLzWvuvxQ85fupg/ww75lWzFKm2bjsUHQXGo7UjEAytjczuT0J2mVqtUSj
Z6Zutxzlt+ogrXb74jDGdvZ45NnTKOnju6eC4TbZpyhcWgnNW/fYH+hHq9MHLBtG12RV8Zo311Ly
YpoFD1Mtvl8WSjRmXJAh+TgYwzg/LwvBndBp8StdPqidw1as639xvzb6SLpIhpY95irhy/wszNbe
gg758/Xt23NCRr9bdJFtzuh8QXtiqfYL4ZpK6ntmZbxlutdMfaRFseQcUZ2O61Oi8WcfGY8JsMov
SBOox9YddiTFiEJMY1bd+sKxAdl1c77aVX8C4+PKK5Ml2nr0wQSkRysv4BiLx4HTyEogX/ro8sJu
0cjPxirue9RuayLoxpqzbV3t4zbeCvmqh+BN27mZU8e4UeZHF3SAmixXZBXPNXdMjA5+ZZFRFtIF
WB4K8whZw6K/3pEo750UkOKaCJPyPBhLKUZc5kYyCfNXWEc9ESGzRIrfcVIkaLwg/+OBwxKbSh37
VXh9Ge6uESJQIxZH/RZk0cYpS5OyCO7XRgZLBCXrD5LCOTZsKfcQjCkiciai4iQS8/kf+BKrty/k
bB+B4VX498qneyTO2aFEynsW+3ZVfiYg78bQJLkatiCu7vr01pXdluxdljG3drnsaYHw0DQa7iaF
TPEvbab3nbCxiIwvl698tK8ElG6ycQCnurcYgl8J4DJHooU1DhGR2ZmaC3fVW5iR3SF26lr13NqX
UIxC/q08QPTrWQfxkVkRe9XvKJ+Q43p1fpPGASUeijSZJuI8r7Iva/AyPOGsVDYT4D2vAAYwknfv
hmJcJdLM1VccP5AVOhGXKQSmjS9v51Z6rGap1WzpqDkfddIr0cBlm4IkfSagsQyt++7X22f47tQK
hEZqtFNRQiAqlZxhUg9xxfIBDsPjRUwma05TbPQSpdmurIWutUyhYmIL/GXg122ScsynaFJ6SiJ3
+Z3IlEONVNqaHY4c4WmWvzUM90gePiaVkemhUv9VS3f0UGAqTty+4bhK1d4pBUTHHJMbYRBi3Vco
2GozuyeS5qGr53iJ4DKDIzoPs4Bh6F2t1UvyxM4Kj9TPrv0GKgwopzG2VyE+NMbVecoa0fuoNtld
UZC3wb167nimtDAdl0nIAY+V98s4WYDTb4Yn8XmFDJO8vHaioLNZjzkNz72t9YJLz9zax4ljd4SD
7rYnnAUo1MR7tWBKUvFQ9zrbpRn1FZawMvD60U26IgI22qJ9huAq2UGw72uLE2PseM3Q946/9PJa
KWf0/zYV08KFxVqKTisr+N8IvVgW/ut/kTEajAKQmKtiuKvw/dIT1tAGAjsW+jUy/VkgPg4e0AIH
jpKFyXkGzpFzviC8MynF1FIdZpioh6XRbDEJhSymiwzB9sJl3H0M/CK1pJ/eAxB1m/++MV0VjO/3
oSgjygjq7Iharj7p+Cs/aP+oRHxd+/Jszum0aBqKXxCNZJQGS15BrG7Hij6W1cX5Dmd4ELT5oaFt
OR7Y1lcol2EWp+JXplv/3kh4Y/5uN4tIgvrJvJGFMGTku99Uw9JJxUBJOtPQHKhky5k7UDLl5jrD
MmhGKqhkK1IcAQlEpMNMBp3kQi3dW9G8+kr7nyKHhWaCJUIbysBWyAsQurxSuoFkalk79kPn/Z1u
dGL0Y34ZiZeWOlWs9M4PM0dy4IVENIRTo+Zi1ioGEVeGXhYWEx8GeFQ8+evnzh8onYQl7uQBYYa3
u7uXzM09EepSQVVaOFyYhM3vRRndBn6n42PGsugHao6b//5775Cz9u3xOuSSrJJMT0a+ocph2vUQ
/T3asg+jH1lFoCrnR759PGG/M7KbME41faqW3hAPvhgntlnYYy8JGnPF88yxWRF+34/pubTFvBYL
A1XtBBZUIAT8ZY5FymXPBGUrO+QMskgpsX6GuMiYJ6BqPcXfV/CKd2fSxGu93P+UxgZvwj2HnpKt
z78v9PlB7MynKyhcDwwBkRGb18vJQHmC5IumGOsMiDmZIDA/3OuYkiAq8IeS8Id3xnbw78+ycv9m
TDQLX0Ps4AB5HhLI/0g9z1kvYIhqFxPlW4XjWnJJWVaC3pWDH8tTLsgSNvtX6L9osQmTH9TFL6T/
jV7a6P3mMKHhKmUeoGh6ZlOO7aA7E77iFio3rtaPeMenp3A0CyDnqJLdgtYn09tGKV7ZlIddfTcI
hLgwlXAMKMH72bRsHMthvtbxa6oZmTkC4XZKkTnNq01b+3tXzSeoLa3P0z344Iu2dlrnsnvT0WJA
8etu8+MMmNpGlbuehOJKoyi3Yp81tN/nc6KdW0ANgzEl2VyLmU7ONV2f2CqIqAn/Oaa/9RErlcVn
fjxgGrqpkwa4TPH+Z779hXNMWixbK+y1nTV31cfB7ssEJvhibS5WiJBoIQBXLyo+x8Gfx2pVJxzC
1KTSGPpv19G45HwNs9wYSvxRDLu0+G4qUqIMYi00B+l9LQqlBFsI2YG4EgKUzNQ/OMqQ64aFkhXg
byoSBLuLBp3sLbmf31Unf4um1ccjwZkrMw0/V0N3n+LnvO0X7rehE5ez/2CS7KuMmRPWitaJpLyU
lQeBSw1ERZXLXh40dE2nEj/9CeqZGRFMeuLchLWrpq8VN8wxIDZWj6OoXH+mv43piljveGhXIE2i
OL07syRTBSpxyg2agMQetihGnJ/hCNQR3bbIrqz2Exf9cUvrG9PRuVr53TlroRl5Ra5Uo/7+6r5Q
wl+DIuDb7+KJD+cbSntBV9agvHEylHJO3qtsb1EzapOWzI+gA69rF15JB44F8w5MfqJ2nRtfFTkS
aOi4SeHJnWUC5xF0zb/k92QBmCp6g/mAQ6kK0I/cm1jfpLCwuggOHu97Py+gJpM14gG0bLMf6GQ2
5rBJg3J7KCtMVoLpPHZEjSPpccWxPCBX+l9CGuWdNQkADcNK5hAS1r3xJSVC8er2FMaAL6OBTxCD
80xOwSgmzVP7Wa8sBpDLENy0PNrHpg68voWnCf3mJtJgEWs/H4W73bG533H0l3Ty52tCilna5oog
9jksZXZVTnFEX2gKCpplkvAweLg/0JwUlT8nik79L5Vs03LxXXBm0OY7e12sh98brvIvmGL5+D39
YvYp/9fYFczHzpDLuc4sdymVHDH9KIfsATLT04qjjdwoo6ARqG/uP1a07d4aMPmbLz8yfwImQ/AP
cY4hbcYI0SsoRUSXcQEGq9eZmxvIiBE/8j5xHoqKTSxF2sNoJgu/lI4CSuv9UxotQa0bbO0K3V4f
qdtg9nqz1R90XZRgAqZJuawaBcD3EuPkciAzU64BBye89DLFCP3w1KYnyqiw4ZOK1MxKYJiyY3Fo
jaWD5mC/u38uIHCx51PVrHg38GBIX+49iCyoVDeroBIsIz11eXP+pAEOHsGRSH2Q0q38A/LLKtEw
lAR5aaV83zIAbPNMqW7xtztjrN0esUugQDM4HyD9WYTEIyhYVH3rMFN7S8mhMcog6t5Mib+hpaSc
ZxAwN4RfkmrsvSCpCFEs1nZt1Vsp3P/p9fGuS15ThzBSG8mY8aCG7eR3KGeaX177FPMAN3qxU5Ft
mhp3neY1peS8hAm04kRe6RFwCYQNCVl6Z72o4dOhsH+4h4sCQ93oAJFwb58wmZWmPYEoic0I1XmQ
Isu2lO6zbhvFxhjbr0nj4X6lpLhqyCsNGp95+xPtblfGOf/g+W/BTZSjL1pQJMY7CF+Z6onBkaFp
PdmjmerQBcWJ0n9mYVRYsdoVHghDW63KfQGuX5hb41fgak7gZJuYx6wO+znSy6ElukRCbH0iu692
p9P30NPvLJFXEG8T5+ROd886zyIRcXk8CSp1rtInNIGFIZ1qApWi230qiRxpM0WK7Dhxx4P9ZvSs
dy+qbPPLkih+ACAuovpc5jGuIpAWRdlj8g7weIf4ME6L99Cdg++GXEjmbM7T9zgMdrqeUgBud0Kd
r/tEx9zaK/vMVSk2FPLTEg7FFG4sLhowga2z15sSgFFxra2OZOLboBvKc1N14OKKY9LeinRaFZLw
13YA2mjv17gZklvUhpdPc9ElkwlBIqMFwDvZqWOyTyi4syh+Be3FQhP20b15dAgRxsbTJOZhnH5/
gcy614OYB8Ok4rwyqg1HOWpTG+vi948VOV0uUCk79p1JGU3ci9gXYeaY3YsXmgJcwWMwr0mj9pWW
A4OX3dNnOlbyY4MQ+6oc4WYXdoy4DAwlr34dfAXIxgLcVXT3duD3ndrk0O4WDhfXWot+1DmclUaW
B/50WmijxlumqaeFUgQcR5NJqXK1vnuXvmfzlqQXWCEPuQxmf753LwsrOuz1nqAin7p8Pcj6IVw5
WK0rTwdGkCubQMbi06pzZ4di0LQeWozhVVt78+HGQHCH5OqsHZbM78s67LUgWwmc7AH5upqYnT6I
vezxdK4LBZBuGkqa6zsTCSInFtzfiPviHPSmpLqSD1xQZJkoYgZK32xoDllEVyV+EwK4xJTBRMSJ
omGCHKgHCgY/4uvyaK05V0qP7gsuF8/ntMcmuRyGixNidPwQlDrPQ2DA5o03FHHW8CV0LYMlvkh0
YNkNY1e+LsaLwFVB/u1NVXaYoeQNIgSJVyKlhGZUsWfNQ5ish5x/9nUIwpNe8LvdbuCHvr4LEsSO
qZhZ71SnXUYI4hxGHez+lsS1lkaXqyyNvQK1/ZC2/y/2wfjZ5/Sya2bU6se4UU7UjiCUNbxIUV6f
mNBRVXpajwNAjSzuQrwsczPqX0ctXHINKC6ACHUY3HQCM6Q+co4XovQMn0zQUR+9g0TRt1JlpnpV
eX+6j3T94Xi0deprwVFwOZeMfIzHvO0nUsIIMOic4krW0F6KHrzW1oM9GjYnNtTq2ueNF/D5EqVs
TwGHFtcRCvaxJnW37F6B2JCdRb8d7kgZUObJ+nTX2lbTD7PIACNgxIF2KWLYYIBIyQUBfddBqz/P
0fU8Kp3/TLDRfvSxqaemnfKyiep7vjlbX4Jd4M0tBYwqWcXBmIc7OFEBPXSouetRPGdDarAoiujA
znfuZqsL/uagU/kl2Me3QwWlcKV3h3IjsGR7e25a+uhmQqDihj/V/IckrGftdmFqJOYLWJf/9p6s
151zFCWU1Me4Y8RVAeo7HstdkclVdXNBW3Nf1O3XbtPuSJKs79UllegajIJOrDz+Fkl5Z4hhaZIU
Erulbvfqb7OVrtMYNZ1VzpKtPrgeHG+DtRclmIBWaOUy4EO74J2B7+SuA00TXTpeQRqy45Yq7zGz
hB9iLLAqdSqv8kbguz5n+pW5SgzqgHtORfPUepXnvUKuiKaaMVs/YA9R9LTDIQWcZtI30gqvrY9f
M46zh/GIf4fbIq6XjskGp9/sg9QCtYIufxvjC/NhRVf4u5ppAcMBY2+oF7iOKXZglgdqzIgQcF63
OjtdJq34/BgVFnzLPMXY5lqLwUknNjPUgDe1EEi8xAWP+Oh1wB8I7rjPLNFVzgBtfbfoVd+VUPvo
VSgnin3qYgltlWGT5AFNlTHORBplB828EvL7ePCA+f1SeT9YISA8u/vs7VJrYaToFBTBoukQnXKH
OCjwia9YlzzUO5h7Gez44RN/D1Us6G4CxO3yKg6q5LoPAn3dPZHrZyhw2FBtExRgFTtx69rqcTkR
h97HBbgeT4XUIJQmagO1gUB5CgdGg9OZluG7J+4olArLEnU/pJNXaryLxJmexuBaChJ9hGGruib3
KImnEwHijVRqtayO3wZ8uz6RU4GFyq/W9lAQqWKs6kMkJ8n/KzjK6DIb5lV1f2NfchI2aDLu4YaM
kgFRPhurvNpPcBZdyjTaXeYtMZ4GNIdwgu4c4BHgAqLmHBXvWOjKtsZhJPQp5XakgC59QyWim8NC
rP88fBHUX+17R3I+B15dWi+XMBpS39UhHP8jgj5sWedReyza3zGhF/DgCRzHPjxW3R/U3lHK+yPn
2HN6Uqp0mc/fBG0RsEipwgLwSUy13AWUuNI739ysVvQ48Zp9hmTnN9hRGrdGiHKP8QJEOWsoecJM
ebiPmQnmuvhZJRTEus3Fe6YTEopY4ft63NIUDnFT5bkr6MFqXT7oOVPMv7PcVLo9Mzsmjz4Fk8po
rjFcwxop5H5tZPz7acVEI+c7PpTKynxxxY4TVLY20NBz+W134yiIW9WfqKfxEdRksI2lrXs+DYOr
UKGHXMYYSOZF6K248b7m85EHbDHQFB1xzfJsKvq+0pLrUIjBoJ1Xqkpm/zAL7GIyBkCYIIspss/s
p0tZ9cjX2zfr146JCQhwAckZwoQOzKULKfMmwZHnRJJz6eqRUpbnlFbUnkzWyLrpGeWP8BuQUTaJ
7Nc0G96BZyMj2dtRGLm8Fdc84YH5guPq8dxz1e+jsK3/Qno1kMPSokHQYjY1Gj57YjNKQw2nO0Vg
jsvm2+nz5yPtTa5vjH5gNTKo51/hv+AMHEmupNiHX+QjlF0NAK769fRlEiAueotwt+pbW1lhYPtn
Vw9jisFOkrpcwMjCzQp7zfbIutKj0+6bvla36wLYm73uws/rDaohFmbDhWRpVIWl0cMXgT7X8SOl
LdG1HB4Hf1VTcI3VlrLrgnQ5IlgODUdn+il9RJ233C1u8JnOnNW3E8hwNzthrmzGlUtTUX/qC5tU
ZYVk9RjDkAqctsI7h+RwstyLrYt1TVhfm+/+PhbDvGALNr21D15hHhQfAVyvPWteIR2kIxI4d6Yo
zxomdxdEGnMP55XM53hHvMhkxlgDDX/SYt/kmj7/M81pihiprPY7fo4Efu2N+MHxGI0XA1BR9z5l
YTe2mwy2RQAFmqCEin06dlRLk2MsqoytV9SFI+GZZSttX2wrKlZVqEvLSiSCiw2fXCBiOeyRW38r
9k2v3OP1r5CmyayYf5KPcjxrTZpN1LDx0MUDXX4uGRl8C3OaZPZmv/OQZJPh5yw2AmmmrYSeHusT
W2JhhYQ5EC/fWXCS+tzcRBfXRLpRKyaRoBRj9NJ1zeHALJ9kra18/VrszrZGcnS15nnIkJzcacN4
mocvk9aYjMA05MSmTaZhUyUoCv5qLQSRi9Edxyjkt0Rc7AFpgq2IJM7YIe5WT9g6GpzOD0AltBKI
cd+dRHeSqAp2zcb0TUcdR7WgQfQN3xbWagMUbaWDycHA2vFyCHRaW5kZNAPTOHcqADLpFQRVse0C
O5oJE+qWKHAu7Yfc4zIjM/OWyTAAZlThNknIgga+wNRPZVHogSi8t1FtM+f/aaFzx5+0TexaLT/L
6duHjFE9SvZsG6AA0wszTDdmEHeFCOXkN5gcb7RzBC697HPzyGGcCDuduAhi3fvjH+xmjSTeRHFF
l+y+LcM6ScBYykCTodvtp+n3tabcLgdikMNXmf419VWrbW4KFzYgBsRQZgYETcevn8rPn6VEYilT
8KdMQo0vw6+WB7S/j9savzgYZ4xGs+K9dGzuCUbhOPdY1h+OZWFcoJwXMyrx1JyKscw7abAEPDqH
3RZe7ydS1hBfYDtQOSGJfl4p/5Obk/xmaP+MTVbmepqzumzjOAKQjhDR6KUaP2xbSP18vWh5SbVv
0ROycKSaarogT9m+4sSdPCv7SsGUcECs/7CJwHquzYJl6XljcFB7wCr2Vd05i/FlhHQPHRLD4oAB
UyChBQVoP//jilcfwUNuWcu6pXJKmO6b8vVq+D32KIFUV7o8sxxhQXAYZxnCpf8C2R1JIbGN3Bh6
S0iLxIaXCuEYVKx3+OHxzVGJzTA4LuJOtu92wti0OIbP7zxdh/0SSbM3l+DwMZYHde+90u+rzrXd
/Pn12omyKKg84/7RQ+N4XKQ1WgjVl+Vl4HPtEiNWYP7GjOPKU8gphyQyjSWyDLf2Mc8x+RRVO+/C
LyvQRmAmAQVYGjJHCJ94zRnsgrH0PaQ6kFxmXsmcMbDKwXB8UJr3fev7TXx2vFt6HtVw3VN6dyuR
gX/2vdGf73ZQVzy60tCW8MaUae8dylqVnMo1/UUnKEK4p9y30aUZaEe/OAaS4uRePGZ12VuxAQFt
rKMmMKaoCRmiQCdWK6UMhHunWg6o10noqkaPLhseBacrRwl1OAlCOdDbuCvzxiPg54RvQq+ukjLr
k8LphFTfeCEr8haf3CShgGj3Ei8+qwz5xF1eYKBd/SdJWV7/YnI5fHt5hcTUhrXNv8HvmHUkpzWu
oRl68w5YWNjE8JFTMrdqpATRwvdEyDsUOHzsaHKsIWO1dc92uQjPC/1nHPPcq9rwYFCSJMhXS22A
B2X4jV1P6x7cbKuBDRzdU8jvOWEgWofVvX1Cm0Z9KIb3/CBw5W7gNti5khtk7NtX6RdXD/RDjUuQ
LU3dfv8l6fOLu/Ip85SRcvG9xjg+otWEdFxjUds99uRQ9tLc8operLV3yvOG4uw8tbpDj/EeYGMN
QXFF51hXq1kzaWFr/zpI3qMG+gqP+JKVK6lgkezYMh5lEc9PakDO3QKDRlNiSOTg0tRrRB7CjfoJ
c91v0b4QfOWrfY/B/85HdCmpw9JNA0mJXhTrY0xRIDqnF0GP/jrQ9rM10yRS7rStrVB1D9Hs6Qbg
kBOGL+Qbpke57U0Xlna4dhQ9D5SxpX7+EkGLhO5F5m7PfWyUEQlJQeSIerQ1Gq7csm8XfpwxIdaj
rjn8NVHVeXE4NW74p2EUDxYMp6llFI+hiV0iRfoL0CymmX27d19UkDDnnBfnpxe2iSyKbPqtoF55
7y4cK/3MNcfKzt9E9Nug4AVUnsc3U6bRjzwWGN8Z31xhpDMi3VfIvqUlWQEfKJv8D2A5Up7/RPTg
UxfMcfgbaOSy+4lmnceJUhnDpFWO8NLWZF83PbLo0vX/QYV2RdKmKocqWC7JDTHSWMLFJfkt+cL2
TJduoOyViYOuXj4ZfLSfH1jaP704kgV6+y+4Fm31DOpKDbs/7dXRbDZgkwBfD4XvrTcT0/5QlDaI
LMjz9D33t0BXd3uVDojySjvehXVZXuZYG9lP57fiUPt2piG5k/0fNo4osoms/qBSNYhsybc2geuD
uwP9zDRvD4Fg+t4rqJYIrWwmZ2+Qr14VecZIbU4+tH4XfPHKidswJiplvNNIE+XqkL/3+H+rq026
wrPP4hmTE9HD0rjZky2M2tGHL4NuNb/aBW3eRbUOyMZ5M3AYLU1hj6ma3FMVRZOeWrKRmTcenATk
ulEM+Sd+TpvVfE/8Q0q9EY/fl5mLBC797kVhptwp0OmKXzxf4RT2l79uTtfIW72mXGftoqlkiCTQ
B5bRptYpSoJLBoRYI6dpC4SO6hVY4rcmr/DmujGB48qFnXk7/V22k+Z77awQbyMJ1Do1ROaCPveg
1ED25mCGIjoB9kIU/H9wC08hU92P9uQX4fKurde0t8Yf38lRm062VYTc7tze6PJnKwVg2eTX7lPc
ee85g0MQn9Sw61lUMEoTALR6WM7e4CD9myHga5APkqtig7h9MssvPfiV/rKSQpoueT9vgypPM7Yc
MdCcEthMgauY41k78RtxqeUw7N+ntOi5bSzEDEHUbblr1SCF6suHoGBSJ5Xc3/AuURlsbhnvyY5h
KawKWrD2HeDtfc21ZerbFdSYQMRtbeRdXVH4iW9tDVrZW75ExguNBbpu2YgnwczA91qaQYRWnFoj
jhbsj3NWVzHlp9+ZM5FtRVXjxNnR6tv6gStZtH3SHBUGlske1RaI4mljIZHB45FF59q3aSGZAKP/
/O4ZCCxf5WeZm8Ot61TYma+CWZS+y/FW4wKLGmiy+ONu6EQLhZhMRJfvwFy2I4j0EWNotlYqo+Iy
2iK+pqVG3QoSCuWTrgi+sNdYCjTS+Vvl9B8tR/xVySdzxI692v5jO73w8+kPTHKFoqRJLnBOS64G
qXPGsm2hpzS9/Umh7A2x9nRcE+o/YfdCbGwp8nJH4jNKQFt0efkaLjUVwMHiv4DK0oD18OSJiZmU
+fC+c3Pf+F+Fklp+Hk9BsrD5f97MJZAxDQaetOu9sodINOJNGpNbZyJdFhDyt/68RutEvsJPr6t7
8oUBmqYy8OVQ3mbccHl8KpsMDJfhd+V1n24E+fpa7PFN9yDEL5go2XLbX4MolQ04NyyI4Myv9ir8
tBUhRtKildZ+euTxGuybx43BgtDymqZQx1YvvJYuwjvQyr8A/UqUk3RJHSHifemukZHSw65elLto
NqFycA7+9P6s7oZedRnOWYQclLOq+ECHRP7SENyAQiTLjJ+vz7Hco5/UWiT+bmU4a+NVhy8amBMZ
ikYmasovUN3oQUZpB0ML8DgmIhyMl8CpObNpmmGMATVej65tPZ5S2uVe/q6gTQ9HRaheQtjLxXmn
st6ArUkyuFTyl92Y63eiNFEHUlSMoBGj7wWwnYaK1yCdYRuFQLsDVFSvs0guxpM+n5dOTYdm4WTJ
UCvUB8JA9I7Y3z6IlPyCiBaJpvOupETYInrxUzWL4nJi7id9pEHJsh/IoP8BMfGOuy4ULzWOeF+H
AVI8Cnp9MAn23YTA6oh3N9XkE5Noy2rm2pDezhsWmLIIoXm2OJDZ0Hb+Zi0gjPKsS2I0TtDypzhi
vj3pgHOL5/0/dcq7h/Fn5OTr0nq665Ys2T/vImOwR7NHFv4+vCkgpmMJ2+T9clXhapKoU+Zopnir
Gq2STqAHP6QSCV77GIaQxH2zwgG+l2FbviIGyRjaMXyjWwd88pCm5ZubOt4ql234lJIbwya/XGfJ
a/Rd9gYKzatgou7yWs//R4PorKzyIyjoWzxVvy6xz2XAZZO2NQlG8xXndKmUUdGwunhSd2++SX7S
ulNWy7bC8t0f7OX5v/hPZJpkq6VAvxTVoAy8snwdrxD2+5kFo+UgcHHXNrQ1rWRuEiOUejdSE4yU
KIM5UYnhegzh8g2ijj0qG26iZvJT4eursfJf58m56HHAsMPIctxWL/KPWia83jmU1XhhI3NHTVM3
Y5gt8kirYiaoWEl3HinkkRTPbV0+Gf8Owt7q6eNiiLeU8QgXSjh/cAwU5AIw808AMf3ljuo0//tX
HDbyOxvsx6Drji5mmazv+LpVW1dKqlqYMFkIiROEiNLe3TmGn5BcV0+MxnAcu+X+QjoPQIrndEak
1eZxd4QPp09I0v/+MZNPeEnPwv0TxcCIxX7XPTzV7zRSukK20gm6PU8R7dbSN7Inuup7w+KlTFet
WqrQhFsV/xaNE92epbp+Ytygc4466RPPlX9I+FSvOVZfFvj2pWYNPyCLty2kGpZcjeEviMtXsqLl
zSkOtaP9EzvfMcIWd9HreKtVIIx9WTpKsFLYQ5EFjquh5lbMlYiNIarbwLWLfJJL89Ws5xlnRHd3
NONhRc0GffuRYAJKqsgTniyLR1OHObsB1IOCjoRGi0cw41jPfGCr7AfIjmL1bv8yWjquSyKsr0xu
8Y4Zc8XTYlv2elhj2ClUb2vs/YbQBF9svXBgWD/tTXOwkXS8am3r3ZxkRfoKIWuT6cvm/clPz7Gv
MdUZHVMWWIhU+gUZLUk5uoF+Wln3J8DEyD3dH7nDk5gpaH+OItF013WZ2r4351CIpYlS6K4tsmCf
4IRU5yiCIlgd67JVBRr/ExugoSF7xBEOLmuHQSGFCpb1IxWAo8A9x6+1DYC+osO8CSySQm6GeYEw
Bp7xHECeknTjztH5hfNswwbeTTNfIs5JhEX4WjlA33iOBl0IJ3RW8e9iOcSKfX671lU0IohckJEK
52diG8uLfet7cz34vf22Z5efrvoqPCdvpQtOozdJtghxRTdTOvYU9dd4qa2HIUzcEY8WWO2ayH9h
NtIMbYcHgki/eak46QLUP9mRpPi+Ib3QtBgmoKTUGUmWoZ1TrFvrEJ4EP0bnk2cg5/IdjgSVav2K
4LWK+4Tl2H5nYvcIUEOtM/2WrXue16aqI4qaDWxBLGCTLxBdjaO1hePbMJFP4SAfiM0suWzvreb2
5F6hIpnwf8KrS9YQvmYbbfmyM6PEEeLYJg7p2StI04xp1CI2RRMvFcq48mr9i2FQqMk6Tg1M64br
mlt30AW9qCauqOlJ7KqqNDWcqVGsa7MQKCfrmOfVhPiW1z+tknKdlOF30ZMao0N8qykJyDxkghGS
3s0WgV1uZhka9q2GaNruAxbOSW3qdP2BjPxi2OLkD/0uZ4I25L6NfLiTXPLDY77KM7QmsPNl643C
XwrohrawyCHtOnlASCgf3Jiq6lkC5brCEjmHySDgejdVvFzHRbHdfxMZO3Fex1MgYlWPWDdYP4X/
pXvfAjIV/5HyWZIOiQGQ1R2QljvdrfuejSc0+bc9CXN/EY77Fi3nxjFeNkHUznFFgdyIe0kGyK5G
wtyZQct1nywyKesQ71i6iNS2Nq8RK/5hv9tmCCIyjKZWUwnhG77tOpHIasIzwQJkuIKyvxY4JwKn
MCfjurzx1CfJ72953ozVPWzJPuDho6y2oioTHsoW7IoMA/9CHCI4U3+IXUlzXY6Obv7VYqMNsLkn
lh9DP/V7IQnzLHvck40mCAjboL11cyfVS1RviTrrsLpowPbL02RbUQ68C+pn9ov7sEw4Hxv9SBZS
Rf7S1dPgWIMpFSuW9Y1IdyaqqfEJr94Lf/eyppEs616ZdeDlchBMTyR+WOvQ0LEyT5R2EPnhRXbY
9NWC5OR+3MaRhI1tpK8mfvHEfmmkrL6pNcYh3At56S97HsjeP4LLIvWsZNzjkRnTW1k0nvi46iQV
RLFzdqGADuomH5MGIH0qrPv7FBc4Qm2ZDyDLzOGfICZtZXGxo+L+vIvVncrJEl5tAdqv7tHe3tNr
8Hqgg7VAkAL3kRf8dfEyDX82tnCvFfR/5/jBbkPWEQegb3QPBDD5kzUiwke1UM4KcA9E2sJZLJRa
AAJu9t6f57InxexaNnXhLdu/z3zsCMJh9TDfvc6bhoaHjfJ4FH/WsOoli0oMw1+g9lb9rHq563gF
qKmwyYPcpei+KSgrfItDyW1GzqilyW6DiuKeZ5FDXzJqv/r+vw6RUwT2M7Q+TEAixjmebmiR60QK
GhVViweVBFatOJc35bwJoFMELlQKQBHc6pqXefyFk9DfZwuHhw8svWmYXXmnqelnJCcybcDyXC4u
Vmj3m03P4l0FVjbV9abCJrwGwe6zP2MJ4gRZ/3oEH0qNzoQtHJby//LAiR50DZJbxOA8woFIy6m/
GlhBrx9ug/KipwwpR9vsWwEUItNIDUngvh0UNw6dh/tnU9GyC8DLxZeW00+H9nPEZb7+SwoAUhHu
qo1OXD4PG7VzOxUdbmKWcthMBBLk87JCQJpVpvFgAeKf5fZX4RvYfeGC0SqSbLf2wG9+yaMTQXZv
5lXcr/x4zbGRmPS3rB4S2GfvgrL96UcyuTbsYorYi2ck95gKkuEoTQIjG/t778iHhnuNzswS06XP
5cKhKLW8sacTjprS7my+AShnKapYiEDKXWHW+m/0JIrcXEGV1iGmdJ/oqiNOHBwt2NbdSRk0ZV7+
yabtIjBTPNq8YvpbF2NfC/eB+SKiCXsHvUDjLt0tWC/zf0jahrVbu8pKHceUp9k46WsEkIW1AGCm
+69n3Y4hfxxaKKR3R37fEcCm8aKY9K2eSOl28PRA77wIZQtPQAAdKfApy+12O2uFG5ot5K3PrM08
o+qAgKLJLOw5TsgxMQyGLHKRMfJlBY0RB6M1hlCeKQjI2LF677XtNKzMgUBzRhE7+cOiG09WVJm2
3qCLDuhu888JJ4MqxonT+mTUcMGp+INJ5FHV0M02VXYG0JdV08OlQc/172twXiZF5Ionvq8xDqH1
eSDCTjlpf4QMJLEUhxmGJQmvMMSmuXUYFs43i00Kt8uheCUMgzDONEGF+ujpPeB1+VJwCT0id+ya
+AL7uPRO7baQDHG/gXJjWU7n5O0RFHQaUGvPp4QRtQlB97NvbL9jPVrAMpRjGYgaFRhn3P1vEEQZ
lNUUYB8VVPpLuR8CWKpccxfLj5FUiKBSkTIjvp3BkbQacM6iSexNZxUpKBkFjENlMP9oMTOpYlTG
wQSK27FjLw9rO9+rgNQR2bttCyPXKIeAOTvGgzm2n6hcaWvOcbiC+MoaFuwPDwjjsM0oLXAoImxv
ApLZijnYLzg+gcvUfR3gStZC41w+XZUX9BXsSQhOlf+VYBJXnEtMz6bTwmIb1y4fydy7PbG7Jxgy
G52Ta8gg+/UJNN0mzh0IkGtXbWY2HW9WhqZgKZcB+qTYq8Sem2UBs4qulN94vfUy/BSNG3Nr2hxP
CrX0NVuCmkEVMDoq06BBGhHw4xqiszqkGyUN+lbJyJ/bp7DAdfO5xpEeffwQAEVM8jmACoF16vR5
PNONiuDK2sqQDv2lctKCwUpfiuyQfaWaAb7UdUUosFOWOoFNvnpV5HH3ZvPUVrmkEkePSECBBSC5
U/WeoBlTk6EfXMQTnHZuSReprwM5hTypcEyxmhsTgpNsUWyjro9gLDfPj2sHFXv8TAwdAflqLInK
Pav3QpL5LAAEafMQ01t+u5A/HJk/8v46pTElL/0n05iljMqJGppyTLU4UPn5/OO8GK4FL2jL8L1g
xVq8TPePgOFgUIELlKOWTUGeXUs4iueheKMW6BLe1n569zle2uiHv5haKlFyk/FCUL8DDfQapBoa
yLS6fAatJiFKxbs25eQyqgpJJ8e2y7M+/gYZ3OJMSRegBaLfYLmCOUYCkGnShUr0D8XdrcihQOpy
ZyAlo7/4ii8Ug3qw/pNsr4mPBk5Nx/rSQdnrRGS9hAltDNAbwsgLQFpX8Kz4xptynNtGG7en2Uqi
iaFOhiqVLysMWKKYGxEKTTvzUQqvD2TF7ZVwh8c1M9mB7yKKI0HgrXe4K1Fd8OmslLgOxYj4F/j8
vbPGQIgwfn/GJxdRRPNTxFAy6yXsRee5JTdXEVzmrVhNw5rxw+UHzBUFPHtKEdGbxEvCX2B0P1gk
ABZa+lksSRg00CiRB7JLW4xe+vBXXqoQQ8YPcoeCzYZfIb5e00nc2EwcbNilEi3Dzf+eAiedWUd8
0HMBMT6P2NyJ4KQ96K7c6qUcceMTOuuGfzDE2jQNB6DFmiglhXj7TG39CEyI4z+zYpY7pMnmUT5y
/k7uOoDB3EVL/tk8UJasfxBeCz/YTjr5EALSbGex267+ggWetlLTc5Wuiw3Rv2A2LhkrmfIQOyxy
NDe7SvhL/3b4WoZ2rCQ2r8M2IoSoRxhRwL21geWSWdspp35GDtHAA/3MVpLzwB34zu/HQYLTpg+i
XFNEhfALHXB/FRmpS99DKmgWV2F0a6HXG7vOPhodHDEOT4n4p7eTbrBg0tVFC/GKBXXPntwJA8oY
7htS4219sMqN7s1h9rxMKVyxcW08BYAF0HJ8aAFnzMSFlFQ8dHLU+6CcAwilzIXVqAzNryLOtElx
bN1ARN717lxIn46+QDHu+IoHLGf232Oodfi4EUdiPfxhELoj7gY/Ns6mM5arNWmeTNeXIrs8FADR
jQRkBf5vd70mYbwmdaGQvWL40OCLRpZ6IQsS1hkJ3MxCesQnitbBfEQopFIHoaJ7mILwX9VIOKmA
1ngqwkR97jNVlkqO1KH7q7z1/3QcTGsJNOScKy6SGoGAKLwlT9lTFdeuq/DqZgM/sRObngL4XQ2I
PLXaZHr+9ZbtBUdd2j79+m3mGa4o8Z44+fW9tslxr7FL/x8M7I6rSdbvyqLq0FlUWsB5xTBh+xQQ
fH2H2bFKoYJ2CXkKSF8g3/4VAqY46fcM3/kAUMsRT+J5NywfhqWPiOSVCyNz1XllzfiDYXBtTEFh
lR94z+tsVoZxd1HmNcPcXogR7NnrWaeGpepWUkRzDo/Qmx5UG3LXKqBPE28wD3VaWX2wrtntcBbT
L2b/8Yqgc9vKrpS9YeOsdEzJnYJnGDpxY8WdRywclEwxt+LgjVMld5O13bcDn8vK6Ea1p5UcY3Xa
mOjWzc4o4b0uke6bl2QusasCwMOQHq7njCOiIp6YXR1kMc03z8RtcF+IqZ1OWe6KeidRr9DdAoPs
702y87MlNFxwgo6ldCE/lNNfvDueJ+YzRwNHDIlc3AyWGeswQtl9pFmj+aVKM5cM4o6Bc9BZvqHq
qGZTSI7NAsfSYtJtfcRg1JU2C4HQSgdrSIXNAwzK5D4mHQiYK2utYiDahyFWsfgSBPsovEz6OmOY
A3BHZ1gi3vZ3bIZehYTBCx1y4jeOA0yT8yO+k5OfL3wUKRHvvXG1JP993SVd0Z2rh3VCjfcaYyNe
UoxqkrbujaLde4U6mD+DzsJ6QI3oLU7Yuf34W6U8HvX3PNNxycjsOxt9i3eWpJPfnYvykD+F4soZ
jp1GDupbbdbQEYE1qO+sWh12WVstLYfEeTw9l5+8iGJHmKc7H613BqqecO4SISITpNTnDbm8Dtlv
9Lhbbf3xGOZSaxi0+PJXF/cn+sXsxr7nPkcGutu5kpu3vwSEPqWFKcbB6kxszNIrmbWzWhSbxYQU
FRaaYTNkUanJa9/2Mdy+vPUOqr7vykr56U2sS6gZS6x9P+8wiVfwrlXjbuHsH4MPCGwoh+eG7NzD
/Lh56ApGsJIfgGTMDWP6plq0UiRiHVJDf0MGbI4Os+Mm+Bo3g+b2irwWFZT67JKg5xeCoB+UhCRj
hgoou6xZkj2gBnFYmUDHf3yMevk/oXagS2TkNXtnnV+3SqogZU9z8JPNoX8iA5uAIdBSYzpAYrnC
HPQv13y+hQ5mdZzShze4IB2xb3WfR390fGrZPUe+dpwLbgAR2JLAybDOLRYWYbhTS1c1d+zV8kwN
ww2NeRsbh3dLgJJtJyKKEfNWmh5mdE0XFJ6SdEJAft8JSrWWPm4/OdATqWlmssxnf4nIcq26yD8P
l6FmR7YTTeW9TZtNEbAPj1sQwyzu1oTszJZNKsdMbtCSo3OI7jPx321uKL68HlXOXKCY4KZ5bc/x
/chL1/cfp+q6Gw/IIA14MPagIKLBKcgcg1lfXA2d0Aa1TqL910RUvpGtCzayBPHkkicgjqfOY8LA
z1qISwk9E6k4TuXjVQYCZTogysIsot1un5wU/HLrdOJnEJJ1CQ5wy38ZC9tOWVdDt0iH/ZOLcB4Y
4k2nwPVt+EZAln8hvZOnQn9CaDuizuggB0C5Ty51cITfbBSd9hxE+HW9UqViFQB0Ec2QGd1Txb0r
WbT6teP8ysO9X6RGa1chyitLcUsLBLYWkO8xeEABAOxJUUfNTUDUmQnA4Dq241jc0JXYai9yJvsv
pPwhaIHcvTzbm5gI5b06wqcmKl2Tft+Y+6CAxyqOOGOHdik/NNUz6PRg3GCXa/0OsPyl3tY1Ncdv
E8luoiPsfleO1iU/V0hGryRlKlfgeG3quAZKUXxUaicXIPgyEs3hg0uvC7dP0GCHVNJTBZtiepD2
qv8FbV+XOKasLOIG94+0fE7y6f/WY1/vTY8nnJUXE91J08ctjUksyCYmtXjxA2bMC6O6k+P9Xy/I
34JZ99VJOpq5IfDDJ4E8aHlDGNS/5myehvvWwQ5OTo5u8jaltxwS+A0EbvcZRWE7iQ+5S0AHB+tZ
8iqStnnRkDHQNLuPvj2jvLfaCvJUI5KgiocdYTF6vizddZnpCCHtUFiuqHQPZGNvg1X3wBFfrPC3
MWQ+WPEEU7eRnCF1X720PHaMl9DAHxHH4a+4MDTNOECRzLrAtXQDx7hCaNiEfWHuaVTRdJh1DzIb
kv7Kjpp9B9h4jq0bpdzoaKcr+s41ugjD1GGtzfbSVByRdZWgkPt0M8rPJ/pNJ/9G2sBIDr3IgsIn
e8USb825grI/hNEc3adu1OeUc1HCOcttD6IuLMVGqKxMXGUTGFRm/96jcNbd5ENCq82Fh0NDLEnC
IqipkOYfw4EQriY3kV/vUEMnew37R4qpUM4YutVNAiUVYQbP9LI2httpEqle+utILDBottHlsJ6j
q8C9mprE9bHtN/cAigqJQuy/P5NPv2hk6EGjM+VtD/zxrC+3Ujihx4ocxD3xDc/hnLzGTDGUb+2Z
CRFmvxzfORUqG/nJ10E0LyIMlNwlG570fy1qS8RWCAc6O67nKHwjVWWIpbjLDlupeEj1/P5EaOr/
El6foSo4kR/PhEdm39mUjA9EvJj9vThiAwy/asr4t+SX6nCTqmAbUGj6mzDSgbyIMwRtoYQek0r6
HZBxzs5v5lbZWuus3ruAVQizo/LPLGk8Yz5DvGfuI5jBT/lCLzPWE0g6ObXdfMKaMsJ2zzPuTjsg
1gGcOQPDmQlcgegjabUwQnb6G2iMRklzAXtF/DvzPeN3tZacX5BHrrX0HQ9laK6GYQ7TFjquSA6U
i6owc20qPX1PDuLo3fPrEJ8Nw0SJozpWNhv5WJUZMLd5RwRdbH3fekQw2tBh7coYICl0CybHGC63
ydOdqAJoToUenEgwmuQdnUM5bnvvzE5Z03CmIUORhfHGwB+iuHoK3yYIvjjM23kEyLCEC3wR6lLZ
c4qaTS4+rsXieQqzMYe6VzChhdwpYPieKbCo/jhFud/Q2VBDbRr1Mdlfjc3kW0eeAY+sO8VjQT/X
0cQzV/Zh0AUoIdVHDBtdsQUTtBlkY/hdJxosA9XWKEaYk4zZeMalbgHAKuyGZPqQ7XOuwBjyawtK
n6awz/CIxeddnoR0AFi5sq2uXZCMwqWHvrujetAY3I2BaS6Snf5QjQ2je9RlQYdfWX3mETgsPFW0
0AJxTKMAS7GlvC+4M1dJka/UGx9EMJ++Kxloyrm51rFAaQFVjj23Ij+4vwHIsCGcBBUIeOyOdsKe
bZhQwXqCd8SsKyzXgs+yGML4Z0PJGgIJGfXeSY3c9oO1pZa9PryBK88dxfjckMgQgbQwCpY5p8PZ
ehDqmVSCkfNXOR6WDGAZ/7uBkBo3yjGkpfTFLvFlLSInqJ7K9Zgm37gvmqK7hZT/5LvUwz9W1OKs
oEa3b1dOOiDMvT0/IC7jORqLc09pxsD8gs2UcI3HF8HSR/MUV7l2Vsu6UEBzHExqB9+rjG8gOciY
YlHn+oAIIKzOXYrc+rQ7sbNPBUwKHbKQok/UQQKZ5nsRz6s1WJx0pq6Mvd5tQU9nORAHMJ0mGIsP
yPkpsq3zUHaF/jedI9SzhghkzfQM7QBfZJwc/GR0yIiIDs9Jd1xQKq7acXslAyyX7s/4mU/pIygx
SXMzCGSmEU7q2EGZtvvmbAoaAwCsN/qZ5epfyqJ2VmWMWUP3RakRj8DqqM+51JO+aq+wgxFuJmtj
yaaqkzIIH6Vt9q/9yjOm0HuDwZjJO61thAyYp5WtkU8PnJA9dAbIpheWtvsCgolsznIj6WiCdq7R
lTWIX7qImqaa9jxBphd7g/H4HO3OrhCxeF7vaM1MQpLgeDz18bQp5e7SGe9nhkGQwIT7EOabymKq
nx3TfBoItqOkVlrvzl3iHqV9QbE3sybtVsikoMOB/jGcE1TdQqmhGlmFoFYYZWT8hUqxFdsv5nY7
jbW/+1mksLt3Ye5oGW59e1rfzmxtO8ViQegI6AmkURc0mgiyIfat1ii0O5ldgKIJ00cDcZ9EL2mE
O9CyUyqHvaQ3Uz8gv6snTXDZYKTYyyqGlhLN+3BesHq1/gf5C58cnFQxPqaKmqB6EgLVXZLlklHK
YWDFPQ162q3mmY1naNC7+mk+Wak4txxooBZ0el+KuDfRJbAgY72/J9SjXkhFXGnS9KzdxMTL5CCN
XzsZCrQYHNCWeOCBr8/sQNTncjqWZsE8R/VTRaIkm4RKCme9Xk18C7Fyl0MghKgRG3WFAcfy5pun
YbmLFgFmWwtANLV+4+PDKGq2evDmJUa8nHFytCW39xWS21uekImx31vRKP4iejk1pajSmEjJ9O5i
idD5V4Rf6wi9rviadD2M60I8xyKE6uCKcDrtthdeYNKLqIDKhxs0ghHTfMwvhJmitvl1rGmlOGwO
u0BPx2QCZWRfQXBfpCrZv2JSBzwJ692GZQHGO0J43dg0XKWYlqFtHUeTEjvZVSdMXxmobBPwei75
1G4rmqZr0yJH+eWur8erzar/GNMQ63sWvf2qEGui3o06zJykR2gqeaFf8Fd5qd76K0OILIQ7v5rK
Y3KhxFS+nMyF9CGT/hkTDt2J0CGRjUnPjYXVRPOuE1i4GeAeQiou1uFo4GH5YjFyw9wdhP5sRxIF
bDRjBlNEwM65AYei6T0U6mJ4fPkfWqXN/9HWGu6GZr5uByFVglzTeqmiYsYC7PP3sXBxylFi8X9W
iEi3DqH6RiBRir6e7qz5b1JPel7ueBeAs6YaWqRO8iH46D3UknL3Mv8flUgN4CHkf8USiNJkRzx1
LQu5w7tFZ24FtLgnOamfIhjnDxmJD21KpYIP4AwiVWexqDWT1Jrzvd5NFJjAiQBl/pcQQauSH06r
g441XGprF5glp/2iZUrG45DZ+PyUVhzINaQ6+X+q2fvIaiDEm2y+cgRfn79Ujvskud713FumfXn3
ArT9RT7dlW+lsvRj/VRCWcMOGySf6+782JyooUCX2un76nqCAJiHl0ebS4SfhImnqGi0qucgWNll
ViqBnRSw38fz087BukQp9FIp1OCOTiszMF5TWm1Hn0tGST+zGh0v2U8AOB6DWjc+cJD6Fhs3V2Bl
TLfp07Sz5GvsYv5JwLnyLN9IOnk/OSBiLg2l27e4bHbcpiC71CnaOILnCexj8B29Sk7uIc2vrsdT
7gSr9N1xn1azyIxOoqnnkePs/cmgZCjM/BY8ZP8pTXToT0zWug/wMMzpVdMwRhIxm3lE9XzWAV09
wItV9CHnTAkQ3RHjro/js63KDbmoUbebhO3GxPtCYo6EyC1aAQL6NK4Abr95NvHLBk7C9Ckh67qy
6qY7rRIDvinhP23Z3+izmDjWAhst6FJDfe83DRuHa6AoSyxPEqL6EN2tCHX3aqW4x7IbDon1NWuW
f6wHK7DmKKveMOyMohrd9p6ygfSsLg2+oOSpEmA2YQ4194a0Z7NZiAdlnf+dJBCYVsVwbiA+VnGX
waXIivT0m117ynvRW5w+JToTukzFkQHrcUTbeoL3exo269qYDPt5FkDQk4Okc8Jba/TOdI29FGCV
ehInd/YiUYbMFD/qdKNMxUxqo1VxaqigMyuzCfbVMQK2d8iGPuckm92ggJmS+zHDzONyAUIbqEcJ
UVJbfoRiq5B6DKVus6wRPcFHJJ3D+nHEncp8X5Rb/OkVZtA7lgxpXYKelgoKyVJlypG0n64LfWin
12fbzdW4QWkwJf+veqkvZAsODCpOCmJ0qbFzB/5TeYvbb5w86qAvY8zP8rmzddS6P9pm47dOMwQE
YiHYjjGxdOCUUjBcBhbvI5ELk0HU37Onm0zX230lNyp6FGSsopftqDFHN2B+24rsoWjxUnr91n2o
BsjFtCA0y2E8EPKb19qxtCyMYZnk2byWqIk3J7fwSM+KLkBMRymSX9iOCjWJrJ46LnyL4drACBEW
r/7XBVsOVUV26nH9yasjG2ECo5vGZfWjRVffL0p/N8Hn2XRbOIhrm2TbgW7dVsnZRvdMUvugDDOz
AAuDkEJyD+VWAfmrAVVkRg54rF6wd/x3OxLp0B+qNxKkzBaq3aQzETFj7kyEnhlEgskykU0OP9l4
SLGapvkV8gFy4WSitefeuvz8CZe0fqFt9qxz3c85f9HIKKxCFR226r5BFJfm0m8tB3LiYFirGJof
mjNGzlbtcCn7E/8DVfhMav7WewOn/fDyH1FVPUvXFsw1j+B1vl3A8TrhGzZa8Fil4VfA7E8il2tS
MazKhCqEqTnJBLTi7H6EHqF3L13JSW1JAx74kuInUZBZP77n1dhrBXGwHYr3Q/NNByDM/h/Au8ex
++hlJLGm65FSTLdPHe78DQv4KsHT+KCxicaiCZjP855rJrsQ1iMM37bfMDFzZVHRhPNESoD3h1YG
lj/YsAiGVOGrvDxB8kBAZOPEGMBKFJfIuFNirJg+wrHcw9zj7eEokh63VT3jkhSPQ54dNXCpaB/O
h5KcbXTy5lzThz4oBeWxETZ5vMGBq7CwhovF3YM+rHgG0PTCgpQQJYz4tZvdAO1fgUehESMlP1Yj
GQykQSV2WdYeCMKB9otz9OopUt0Df542atQ+TqQ+dGMnnCRezltvQceNFl/Ub/yOtqGG25Zwpn5c
WoMFRlpVwGLOFfs9gC4NElVeKru1DYJEmFBh2r2t/1VFF8ZcXCmtmdXxk2vorxabmwf1Qz4HCRdP
ont4kwk2uemDIGXnZDiUw5rPfg28HGVXYeJj8HvqzMmznnsvCgB1w7GnqoDwnfokTbf0xcOUvHmT
KLFTKOm2s/6DQhIDjDkfyUoGAZeNXdVDg24aiwxsdAKqWJtNvMG5vLdRGGmNmW1pKdGlRSEOCSt1
Qn9eKfxIaAiH7SgiReaCNq3L6Ag6ac9w3xpuBZTaF8a1GS/IqTIvsXoGUygmisYb3PA66tZ4BCGH
202TxImxemLmeuNKLR6a4ULKfPwqq7YdDym4gWkxInzaXBG+hKvDHFSNpKOujcALSNZQiV6yuwPF
paI1Wkcxii1D7L2yZLV6M55+9tS6XLbpwxtsqrA8lKaGtuEESLt930sb0SeIBK+iUD/bG8ERznTv
3ja+DMzZDgWuMVPzG8K8k2tot1npbGy5ps2NJ2e7VbG0+zo2LI2H8k8YQISY+TncEAAPrmrGS1EH
5pGKFw7UX+VmcYY4CwfRlZkw5ATgxCydfxOZKae9sH5vHGw/J03r+Yc8RUgF1CyQjX9j6KRmUDyL
RArF1g3yl5WMV+qOKLonsywfSfLty2aMiV/4uzHOkirf5EL+mRqWbV/Ge68a27fabNe0U4gjvimF
3NQ46WitQ/jOdbSZulDaji6udJCTjXgaLehxh7zzK69kXJxm9o6fYt4ktQka2SP+Ra/ISJ3jkf89
KfNj9Hg3K+shINAOpj4xPhYedlcVqJeebTNUyZDnMwf9/O4E0zQT2XWI/tyNEeBi/gc272bUfJee
ckIU6+TtkIk679cyhnRw6ef4v6AuZ/pB1WadtLgovlDxmLzdwfCladdy7aVTiql9Z8QOb6Yq/UIE
TUYejXe0sGceEgUnnZlig/2PYts+6Y81mh/PpAMUFcFKFj/3SelPbX3UIUXtMjeqzXH/kWbhnd2y
/RGoVrmdl7+digpjhKCVfbJr2Gx4suWUUEnWUpilJTObVCEj3vb7xpQWWjpXOZdbSMjUwXq9lEQX
XjuXWtEJHcFzzsoJqLfIVzoytNDq2JQSXRRExxZR5FFRcRDqSsMAYUlA/ThfdbRNaUOnd1PYBl4W
Mbr5wHW54l1P80vu1DN7qz7KHBS+iWhXwxyw1LODHbGmrWBOVlPdbUQR1o86GP8DhCE1pWX62GNg
eyNVN6fa7liEwrjd+sHZ+q3Cta4Tpz+lkV4UAHgQRTxEWH4dHqtS4L5KHmDn5TGapgHULiioSkak
2SgAGCWjpS6JDlo1ejPtAt3kx+NkDnKbhWhzkcByGDI2mSBsjoSvpNrozUO4haTy6r7TBF+etWYX
9KDkwGTBW/6cfeK3PWfJyThJmp5pCIvxM/lR355Rf1Bfu4WLF2BHtOuZKRP88cBsTbDtPKgdK8pF
KKmg01W8Xelm+YxbLn6yF2GTyK10ehV9m82rRfLp4/+kxkJgKhBtysmBKZgxZYQBNm4GnPDOSDe+
j5a3Nl4njt+sL9jBAza5NCtcrcXIu1OWmpqtWN5UuuhOAIypyCJv/yslbLHjRAvB3kOwaQCB7qYN
OYpj5+u65ZONeNYRE7UzeruVEYWIcyBXxcQJBBxvb1vGoSOBhk+dSZe7K6O9gp7+5i5axHPLe5L1
b8L0ixEgvQdOzwVuVrXuZRoVOmQHYevS30TCniOUrjgChB/eiuEzb54DIlFGufMgM+wfQ9Auler3
Iy14dMMVxA4/K0kzt/srekdbbMJqttTFEVP9Sj7NJuq73e0yDnTbZXCeRoTTjW5eTIuV6YfWnW/y
0mNditUrXP75pln+ldKQO6Du5ET8xi5EdFQf0pl60k0PLQNfFYskiGHhOP/7GWmrlLpUAK+kk/w+
ZcqnkDMTfdsOdMOuWLarUPVNiK2R276Eeqyib8pBfFP6rB+ujiWu2O2mDZ/8Zz+il3B/yYhXFyTB
ZjftyIXVAD4qT7xEvmNmDEXh5h9hOxVy4UbsOfu+xM8+whAVEggt9rKNCQR14aC5iH8kfFybruhp
BWTb2AwK3oDqfmONKZTCbwqXLEoqX27KGaJ61Cy4RL8rHa3yGNoD5XdqE058zHPrCnfLCdb+n3Mp
8YS0j9WrA9pv4ggZaq14Ek8um2A3Fd4r4i1IqoHZWn0LG3mHCpVNp6WRRiCyDtCALgZcearsAdHY
psOAE14Khfu5oOhwx0u7+TK6/hCijYIyGDCitU/w1X+WYL3Oq3R02hcGn4T4m9PgLVE3Sm19eMCi
sfrob8EywqU0XigoNrPIl8t2ygZMz/7sRNsvjfXgCItEkJnxaxX8/JX8THUz76NS1udhWjpe00PM
uW+6NoX42taih0UUmNkZC6EqUzmkBBAwqC1S3EpwU6dRgepg6pZgp4uygQqP4dJRVx/gFCls7tIG
HD9W25OsX2U0mSy3SpXlEpODQNEMACFc/V+7t47D1uP4tyuEGQv3sDynvR2keYUmAVVWtRafhcrp
pMbhqLMiFBDSVAWlmJPybSBwh42VWmHCwTTtmSw/tZywgj1mnrsoppqT7tNiZ0qljuuXlnSQnY16
u6QwRSwY7Aiq0f2Ft9oPEq3pURFc3WX76CIkCv3CsTzzDLDPuYoC9ryX3e+SzMJnSFC+XBXgn5Of
YjGhksvZfy0XnZr7XYLcNkvVjrh1Lm+icRJHln72rFD3gBP/FXq7beuMTL6sANA3fE4RLJ5wm45C
3h68v9ee8zttYKeQS1JY4dV+E9QM400fPcBcMI2xNTXPl8niFeCQtanrueFUFqsm5pyNKgowf0T1
bq1SGxfEjHXLcPF1k9Y6MYz4MV9xIbIKJW5pZEBEFpn7p6vl347EMhzkAdxAfswsmjFxEnR2oAnx
3VEzJuVm89DCX1t0gzHdMubuE2eygzf6+U771aVqibABC6Ye5AQeEoMpqq9deQLK/SYGfwMUAyy1
7Ogl7Ux9DiIiv9WSH3xsZ7hn2/R3tsc/IwAtJqmxOgNv2GMLDAbdrhQc73wMvkn+Z4ZgFxuk3d9v
u0xcxxx45CEAR+x9oNZBdH8KXZsI5amnEtWkAV6FYAEgB10d4kBMbKQM/2eUHwF/VPxC0xGpSbUn
TVU14cbUQ+JFmnpnBDiycdh51fCO9YO+6oFsiQo1azdNjqqg5jqMshbZf9qmlnUZStRwZNLVgA+Q
JxAG1oK8w5j/iLvWRkK32w9x5whTxQGIQQRmXKavI01FtOm1AGZMhALRFxtZTSkqdp8rHTqJDrTl
ovW2GuIuJrwS49MBFdzr3YFf8EAyZQ9GIqe6RH1SNxbsyo3uIZ+xMkHpcFm9NoRwIMIarb3/QQ0s
ZLelV/pav+bCliQ+X3BQhVjETNW119As7ZGp+/GCDxmybrgnYhbXK2FdnVWveLzT56GPml6WrgY4
szHUf3lRs6dNis3k9lDRimOGXKI08SMUwDc5CZQge+XlrHOOc1d/62c0CPg/af7FACR9hVNv8v2w
Yb9oJtoRh3VIXRBie/Fm2SsgSNniJJig/CjFrfQ6EvJYLfQB1m++tWi9d8unMdX08zPwATIJ+aZs
3Y1sM33sJsJTSZv43gR/Xfk2ZoEc/QC2VetOTFqlF/RzRq5YJupqF9x5PG/4RAf0f7tAttHDUOp1
nj6VraqzglmB/zhl6ldeBHmSX+cOvyZXIle132Ee2Qys9TxciurCmsE03rZkGpD6SwtW3Xe1fvyk
D7tWMdLnPieP+jlL4D8m5aiIf1SjmEs+0RU/LT9ezJr+xEr/nZDsApJNHXDewnwy9I6MU92JIKDY
w9SiNGzYk2m5iso3g64jrzDjPA06Q+AhZX2cUpTlvuUNa0HXUtUpn5cu38y0m/1XF1g3kkZzT0RT
y4OnLQz4Lr2LIRMgPPKOOmegIRBvmwBk3t34WV8wO5KuW7TLiP6udq7uVkaA1M40FjvEN5ABMnQG
xmfdRfqa6EzjzmijntZIbgCJ3l7WrLbuMkl4jjQ22ewUtQbhSUR6Tk3UYpDEJyieuCwrsCTF3q0d
dYGA18VhW2kKjhEJUS33yQpoSqv9WnlTwC9j0kqvRXJ4qlJbg/BrRmloWQ4bQX9vC5G4w7+U932T
hToB76hLrR89/3oKciJAh+Ou6VMUaXsRKIIjW+/n67QONiosWUT2fJHeRLmo8Sxx0tE3UFCBu+Vn
r64qcYjzBaTYiiGPa0NV3V/rkq38BgMZHwze7v0gEYSY1RlsDbRP8Yi40fm35CQbGcwX4DLau0Ib
Ox3/gj1pVZa1ockQidrIgV/Qk9+HD3dKk1EfCrNYqw645s652L+4XT1i3eBxzlNgshMa21Y3bZ7J
oIijL2tBY6Y+jbthQzyPfN5l0+mP0F6sicn4NlvoKWec6AxWvm+t2whs2ENhFqDYQWB2qS/j134X
yuNom+mcCSxO/c9NXRJajL/Nl17zBmLGodzo3FqZ9eEvXCSm+X0txlj/tHWEHEEaWPqeAWEHHQ6b
BwAiX9pw6oElXPw91zHPywsk1mtljt+0JUKAHRQrlfEn3xvJZU0bAy7/jSAvFRVT6VTvmVg5y+Mj
K758YYjZZtX4tiVfTJoyGP8AJo7TB1eaLRA796Clw2dsWwc8raji3Bp6cbH32PfpLvVqCqzfTIon
zVooWQN0ST9a79BZLA9rWhGCH3fUYJLC0ewF7epu+mtlAR8IlW5XHTKOy4WNOB7jUaTjv3b6Kdbt
oPot4nQK+NRr+x+QTa0Duvh1/vN3jzzKu5dS6QiWTUkdQi+58IcHHUb8A+0O9YMKm2LXlqV8l0Nd
ruUVpGWbcZFRYEMU++GaniOAA+EQcx51eoMRhtTs072LKPVejaN/wYJjGokQf1YHNg2kXJ53KljF
bKQ8Dcmmy64m1ujipLMMupR3NlEe27WVORkAy8RWvITEDqvQnlKcbRcOYr06MLszOaqtrsHhWJQp
GxhI2GH85aaIx6QPwhVJGY9co7c28GyGwNN6rTWdUppc2URKAeAJPBIXf/zSzxEi7gCtCrdHz/ux
skMnaj7RLWTa9kPNmrUeb9sQkPXwijZk+sW/O71QFzcBlFN6167gLTsTMpcgE29HHTj2MBpnqvG1
KzG2W/e6MPNyf9t4z69Gu9BMEHEuWC3jupWhIPCe0E00zxqLsbVkHMvbL7XHvWBCBTb3XhGYF+SL
c309lKrr9xcArYdX/5NfdttptChFgH0BAJ625Mz/VJeIET69UfItVWzLd5DxSBfT6vIf5owOvmYu
PAZt++O7xV8b6pX6HFAlWBH0oFSpZPiJmLtT9HfzUbDKDxmEOicxsjW7P9eElDTYM2h7/jraDr01
5PTIO9Ugec4Sf+R1IFtFMuh8mzcnl7z8XYPZVNPIDs6oBh/dRI919jd4Qh+zYg+lK4guCrVaBUw5
kDp79UwcQhikipYRGn9LwBM/xXyfTopXXyavsXIlNsBK7ZsoOaWXMQcLFsH+dmam+5Hfv1zSsQ2Y
BxvGdFcGfLcRGEnhXLcZ8yv+qKuiFNANxoBdnjyMfnz2PTNEx4jGBL59w/gRUPokhyC3lF1Ork6+
zhpDVP+fx7JiVJ6ndzddmtExahHyby1gnxzV3CoRnsCbG0aDVw3YQuW1e/C+sprsTflEqG5k7Day
IaD9DGInNtOIBpe7cuVi3jcK4pSv5PdptSPO+1K5n2fWz5+hsn/zwbwf5iOMZCOZT23whX9nw/yh
DiO1skfG3BcAIqoRDx8WPm7Hf7YVRf1P+rkaMJ7tmwfhZRVoWZ519dusX8+UoutVs3YhzJd8cCgw
sib1pkFVClOCHN+gRZB2epTsw+lL5iSzNSVeQ5z8S6KId1Oal/hiZJEDlrAY9Plf4X62w7qbnUaA
rmIEZejGZkpYwmbl5dgjHclEMKaUr7Q5J7WDeZZdGvi7dU2rFeMlgF2zuuLHdWetA75RRSagJAQ3
/KERbn+g6nInT33Wt9Lo9ZI7X1DXZw2xYCBCOSZbQsaxXjD9hWB+Ku4XOWBeFpC5I1V2vu+mcbYS
WXR0k6RnRd07EjtWAJP9b2xniBQPWm6B/nX3Sg50x48B4P5XNyjYcW/hTmd/5eaWcuicEdsbk33b
W0XrZ7S33yOTFDsOafXK8+Iij61QghW70WH/OmJ8Dz3EmT7gwOSe53I4F9kHfhHzHF7yJ915zV1Q
9MMkUD5C/q3SCmRV+0BwHNM5SXjdLT9iik4LJqfH8cGKfmUw0ep7/koqP25FMlwOf36rfd3gw9Hy
T9vzkky9t7tXOwyrtAPKUr/ib1Zbhx95HZIVJgMV88B14ogHNdsUu3Xbo2Coo+yWGbvrbuTsbID5
hCiz7gvNsbK9EFXLiyNpXIkQcgwaG8t0kesa1CaopyxOHRWeAV5Jb1QjrxBsfgr6NX/iYgNyv7p5
J72dXkKjYEkhBLkzqyBaNA123lQydS6zKxly4PyRghFcagykm+d05QjDGYWn54RxgViIbZ9PX5J6
iboGNg6d48Ke7Dhvir1CH1j2sK2i8gOznTwboTz1nXDuPEnkJBVflLiSJEFJhI1qhxbnG52Ym9ey
raZanceKvmaKHYq/teu3PThuvJgV8SWIRS/a1wjXhKAR355fY2swnMO8R5KMXPtKcdRqIrranuD1
eYYmwu+wTZTpbfCWk0HJQYRoip6AKZAw3Dp+pZhhksosEdWPPWeWduIFozX5Sd8oIDmCghkVOxgC
9rWLvyHizzu8QwLQ3u6vZ+lswNP7SVTnzuxpPGaSM7X+YN2ebY685LvJwRItOpuFUaVwiAxpYMoE
iC1xOGNqrGbuyvXd4nxqNhH0FdHpp8/8TTobbndCVgGuzydFduilNa6AWbAKuqwkPmHlDWhV8hJC
iOywi7ku5MhTfVSCtRkYBYQv3XZf32ZNvIrvfR96T0M8RzfkD7IGaHy6TWkcbNeotcANvYPopNG5
KeuZA6mpVBDZTWRccqleq7+ITb/8wR/GyUb9jP+DiNZDTVAbcNl4ov1QWywAcU5bT4oaIV2tQA8R
Hn8XEkiRVEaOLMcGiCJ5w/j7jzGTBoWdlUMbbuvAYu0WjjNqtMmuG2xg7if1y7LA3E32OxDMOu/L
zmVK7AXCE6gKgO/2g0xGFvNZHq4bXka9RVxpuXSF2bP2By2l9iYb9j+o+CgaEpq21O+M/SpHswQW
vHvUxfRN5/bTdJ2JS1cJF3v8LVxPacAnaK6mqegwq+v0x+gpzDzvS+VVJMAdzItoJNPCKXwbl4mc
aGcgVpFBD4IpHzJnVLCkErb9pPJ4UgMwjzsO89sDRqKD74zRn9S/MgrcBV7CIxwjX6zoW6pBWOsV
VVndG5BrZX2DOzqs1vmlpm7AmhtXn6ti3r6tuN2RPM/OXRiXU3tksnx6+0nDT269c1l9xo5rZo4t
inIHTXLEfZSEfA5UyZ0XcFPr1YyhL9PAA+BKU40VZRCIU+4M0TPnr1DAUFFgc0FMW18Bv1ed3wB4
6HI/VFHSRqc4bmsib0Yryw37uSdtigEM+TjUDKq3nj3IMltoOElh13XICyvGvLheGkHgiooI7kY2
N1uUruOwrqaBnw2bBBpxta5158+8olI7itvvT7EoL6LjJG1c1q5byWuc5Keu8lHR2oLaEZxEEnpg
gsLa4Pdgjj4k/IhQyrSxgn5jfZ6TJXJZMXNFzoa7BWNoRk52d6YIDtdSkSpvRJTdN/Lh/xCMLEI1
ZDprwn1TtXz8FwpzhBI+9n46YTPLyzLdfD0qcsYKZF2L9r863joEm9e1BNSpsWOzzXlnlLSXhmys
kLGW7Pqr3z9129/5QWmLQijz+dt3+ghZzq8H5j07vJckK3bVgjmENMWJeNi0h0AhZgSo2d+JXeMC
lkdQkw2+ExmIDAmOsJBp5f+LMxTB3ZWtM6VPAgmdG8bt+nD98FHs30uDuu4YVCU8qglFJ0eD1zOf
GuGZMuVpe8mrciGmtRStnZ+QDqZdmi2RiRmlPuGwRTWGrkKOSlSftvQ+D5zlaqA8aE6YPq67LLKP
RyUFtZcy0DS5d6xC0C8RP6FU83PVvebv+X0HeVq14Losy5ecRfWge5UbygT7Qf1jff4D4HylCru7
Qor41k1MfW57j5wCkYG8Q72TKbrMhmK83favofmVo361Nh9VPstWhatPvkr9DDl0Z/edLjPXIRbA
edKQSMcuEpd8PNuBOTHk74ISSC6bBfqoyuTs0aJmXB3ZT0RFjR00Wy/h83uBmeA6ERxDEaxhRvQJ
NX2dbRFVSCpD+SRQeWzl9qqTvOFFpPaXkVgxcHSkabk+WhC7bikwl+pKge8QsEs4AhELLSklBZa+
+lWMAyw2lOG6k71X5QEC2DLEKQOxwQAwOHy5CMkEf9vczpweF3yPrZrIVdD600+jdI5wIp+pren1
7yDLhF0y1UT5VzOaWcr+dL7Q72G1vNaIMQ4UQTQnQjU/ajjBHTPHUDoNph8CgjoY4X5DLzM5PShK
Mzm598gM5QMwnT+cXwa3aLCevKMAdSU9KpfwsnFFalMsr92QsS/bJdLoJiD34CRUgpbBhU7l43FG
tklvnmBgfFx/ZseOFHU+S/vxUsNcBO2y9mR5unWmCnIwMrrdus9l09AJl/45HjjfBId51SS/WHFU
coOispkenEyj2VEBPD2ywjURKN7AHv4gjkvH5O/3pwRxhYFlPCUihxC/s8DGVTney8Rb+2D33n/l
3v/z3QbQM2Tbtmd4hDi6WGPC4oW1l9LHjijH3KmHF2FRI0rC9fr3wqLE7pbMVKWXiasYQP49QbFo
bYWsd0F+N7PnvzRW9G4G2+cLR/gr5skHum0Y4GBjprkyZ41Th2TT6fwzUfQR/TTKq6D0uNxxQicD
hf1l9+mZRn1Fdzu+faCha7QyZzIA8679E8d6mapYARkQW9iGkrvjeJ0f9po4WKLud1VeaCYVB1MR
v/jvqrWjPEgs4K/czJikrXmLzLZpimphfvd5JQcbpM3iDZZTg8IANc+Isl0EMkqzwJHnH0EK5JjB
DQ6wPzZpzbaXFTdQvv1clSSbJVg3YrW2U3oiv3Uba/bZ+Q7q0cPtScptVMJyv3n4oGqNF6qMHQ/n
i2MczIFYJazKUSEnFBcApHoMl/Mj1wkP3lr6SowQCQPgXXxhdUlTC9uOmeCeDc2WR2u7fNWGojTh
wqLVki5oT+z5YHtZ1Fj3RBmb9EuvLq1x/1e+WmNndPOgENXnvhyLXcJo+nQYuPHxlEkVTO8pOFNA
Hyw0A8N2bD2ETQOPwjaRYwGEOUosgl3TiEqAAMPdanvyCGkDZF7nKEiEJefpjUiH/80xHnt908b3
7AE9kXpfkgXDsfMVYFTJiXo6s3gT0uboGawD7nVihYvwgFRj/LCjBivhGR74kjCOwerOIsnl0CEL
VUfoLP99oiDb5MWuZux7oeaS4sMo1wOn6nmoLPi8BCj1yRkiFhO+5y4J/H1jLhoFD5j3Uu/sEVgO
3K2w4cqeSSZv5Vz9ZepciyMm+O3n9W6pCAtcY1srqhmVXkojY/jrk6MAC6SFMos5E+GBhC0qDhqX
iZojJU4/QGu61edHIG8asqlNjjcvm/Vo+PaRKBptFE15vaiSHiUiTcpvlPL77cCMuFwCs+6nNc/A
OyNSGApOsvjxCbE/BGWBJsgl3vq37lQz0PJNlyL2s/d9iivWhrHJ7mrztDQLJWcVnV+I3DZ4Sdcp
ZQUjl7elPgkUMuq3fRygNNFpnqIEdjRJyXhueBRTUBr7JHz3AOEhZsrNv3mZY0O9WM6DSZuq8CmN
A3Dmxq8R6aHfAYe1epv4spnEB36r3rIuBSPNMhg0z/XikxEolQibg3drNUjsW+lwBiiKv7ynl5XU
9leNemUU9z7kJ2+rw0uVu/aOHEAwX6OEofIB7cQbDA1F2KIycJ2jlTQsvMXZu0Q29JoIh0ZU4ADQ
gBrPcLYTsCbV26D8yz5cKjhbguo03IB5cX6ssroC+Tr0pB2rqY7C5pB57Wi32tnNT0HxE9v4bTd7
RAfT6BbG9V1S0H5OreF1JuEMspLzOavtN8MYlslgn1a63+xyySVLKrc9/nW3pQ+ZTBMw9CapXzD9
t4ZMRSe5uXvoOQfb/zuuq6VSWaQAYAkhOLuf20v6aqO6o5ry2yT52f4vWoMV589rEpsBHu3f/Tdj
BLa9+Q1P9w71UvbvC5c4uFBIPCjgOrjRBRwLBGe4PkXQPZlY4JgVeWe6ejbmQAlp5wY0gPdS7L/i
/v3HllLAKWtmeOVbTF0P090BD46vqL26nIf4DtWOcRgoYIqbc1zgWJn4AobRj56LbgtL1NoQ8fI5
So9uzIIIc46yEZLjGKbZQcCvIZZNj56W6SSgtHEjop9J/zsqFvD3XafQzmq1JB+xNoAk+8KJjsNS
lsQ7/ygRjrmf9DwczF0N4Sy8RA+F/tXU8HkAtdAqT9FzWwMpU8BTj63CIGDwtsSDQPu6vK9K0uC2
HlDA6yBTzMh+ZH7kW7QAgKDE01S9+h2zVK+Z0bIhjpfO8RL3MyAgVxL5g/QYuehYni7BhE63pjnP
/9Rj0aSM3WoSKx6mewdUPrL10JPDAsA77tPO0t1XJ7K0/JdnMz4Kd1bSWITWNDivciFyC5CcBqx8
TJ8jEiQE1HCC8wFjw2uDPBkD4rbZf3X+NB6NgYGJpoRe2jLDDkTvjmqfLe3vhyUfJU0Fr617m7KA
XcW8EFhqA068rTsOkAzV9321Ro+Sw7NjpNbycXjvyuX8fW3Jo7tPcrFdXOsJV6vlBjT90EyOaKLB
bBjb7jR9JstM/rMeWj5Hu03viLM5jZJPSFo9t1zAGtxxvdoVMdKHSUl7HNeybRHOLiCUINDuOlzz
k1dTcAj4HvXMMHpPDOIwqW+WD/1ZGzg8yKjeY4oE3zULIN9KMUn2fvpOfD+aQ57GpQ4f2aluJBp8
axD79PEk2KJfAr/7CRdLrn43Kj6nzBLHiJuOT4t5dWe7s+2N9Ltv10rHfvcV3TngdCZFOjS5Zitz
1AT6nI+N4IjokuwomAPxfhVBtdfRO/0qk9Uf7Q0y4G+FpQyHyZCvDx+jftiAHB280Idb/4pYqoTA
EaiT+rlzhJShxSUlubwRokrWDzDIXaFKnZafuvZV0Hb3T0jEvDd/4jnEhgU38hjs4nHtRmsWfJwR
/j/2LVp3hKdChqgQXqNP78qXCWrXmscGRVNr8ahbTABxrhCtvmkbVQ8dZINQotFgmmnWrqZsoxKL
DEGxlh6v8yfIMIejsQyIQaW0MROOEuKKXSgM6BzK+MpbwvgUJuWdexIluG/ixvg8fQGhNmhbZ8Nf
vUaTo7nWO9Pks0eRltToKZLlMr18+hh9qlCranMLfNsdTbOhtMNrqxjE4NLdQcakxMSyqjsqLoUm
VtTXzwDQUc/b33QdeLnnPB2CoiWSkrektxGI++s8RaC7hBFpRqVxrdzpSJO14PJ/rHM+4z+Hvs87
98lqWlZciNxWDLMeO3NEbYOBu1lvLBMd39qW0EIwF9f0F/YoMa0qixX2nq9FknqPJrUZzEWu/U+S
TllvSOIwA3EXyif7Tovj4ytgcBJt7obtghy9sLesClrmRmmgJ6FebSFenbYYXL2GVhPlCnP+npc6
Eb5tRSaIKK/7uVew6dV2cxnbWHW6oQoaG3GP0MY7hT4U02EKp7MBkTpNA7Pf50ciqm7XZau/TnIx
PdCjIDvXdFizJPfX6ReqorRRxclrWi5EsjloPYTjDG/6Draa21S3iAUYsQASJ7K/fEn10AMk9F/o
W4ezHjoOLocC8IArrIlXLSa/6VdScWDToEisvJ/n5hd6p+0Txo6TDS6KxFqE02/i9JRPmY8SxgM8
4Tdb/Adm4uLTVxJDe2pBQ8/KguBNFL4iST7Jsi0XB6i1H/EDbm6I6Wcv5fOZ5zrEo9B2+rXngFtA
H9sMtU1GkVDsAmnv0fkey1+eeitmep4lKVtAd+L1ypGmctpOzXNq6FJFc9nNJDUffmfRxff+jBBp
061lYjuT0igTdAWXtkF/Q/nnLy7TtH7mOdxXPYEuwwy9/sLUk6P9ZzCYP3L0qqB7xW00UUtuL7zV
eUrZlu6go/Lf/4pJxjBrlyA9WMQ4EBWSXbv+C1it+iHNYcNVmRs3yit+V1t0bz3XU/Uw9Mu1nZ2Q
dyCx2qhjXtsE5MnutYQp/0fWONAwKvL9TBDXKf1Q0f415ogH2GHaExsGoy/GRzUBpXxeQnWOizVZ
T0uom4P5p0DYo7zgDmeUwb/5SMI1tym7lokUakAfhxDRwjjq3CVz2joXBvdbpySHs4rlRaHRxCUX
vXaeoj42xdj41wazhup0eb7U8ow6Ah96JIV9y43BF3/UrvtL7JAZxzbqs4uQ8Ao5HN3ipwNeKAQH
xosVHvook532G2oTOVRo9pu1mb1LjJ+WOWnV8ggy5WiT25mJy2QahN4EnCqAh6GATA7gsOxFd2Z3
OGMlllxszAPjF/4gPqWt9aKocD1mpxNpAM6QTSNsbeEZaKmCfM4AYQC9uGVjOprc8C5/1gRcVycM
ewa+K/dDpHNp1WBvGtj7Zs8SpNLTpFHCkxrKjRA/AKLiGj540AcStzPuS1lOMB4JqMUbtL1r6apr
tDD+dyfwrdrZZRA4Uz2AaU77tEu7D+b9SWEGkOBocvHJXWP/8dnPpeJeEDHzegachgVWFf1BmxKl
3dKKR7jprOXVc0uW1k0aP0/SAFe5pIG73BnTlBpTWaJrX8cx6iO0wj7bbjEakMb5pJhTV50VpEw8
te0NMU44M6RghRJESO1r3BPDaoCexNvUfT+Mh5XUsTiVEf0ZgWxz75yX7aTFD273UlxkP3oQZLA1
YkdusJiG3Oln4A4uvZjqsFB6KNI5dms2//REAVMgV6Pw5ci9ErZmvA55x1Ze02TyrhAw4JJmQx4V
95PhvG8rcWxigXU61TJTPQGP5GfE4usG6RLPXySD/c1O+3a4qKcYRdZlcNrzq4aiH4skKBFtyrmd
H7xk0+ali/FNvFWe99N6Gi1eoT8c45gO92n5en42PWN7JnFu32kJfgq2iygq9hsCPnHFdS/sM4Ss
xLceyiSwSvUKA2S+2JKaU1VvIlwtqClnHmZkh+h6bvGt+BXwlmMx1KHYIu8MnCObUeO5s1eG4jPa
rFIkgCF+buD99oL5lvVMrdO2COdRjJYOfKhOsvPimXfyv1O2N5Oq4ajOXUG1duOobjqq2HDa+7f+
GfZTzPuy2wSckTch3y/Fp0UcTc+rHofElZB7OLsK8uFdmsC3jFLVo0f0tXSp+MPEUeuXBTVCfrXQ
1dGT1sofVhvM0LeP+0+gIewfnZket14SRVdsA9Eh1SGbot2xq/jYy+wILbyEPJKXcJPXXNPBuvk+
NbeS1SCOXaAtOyZZ2pp4sP/tUNX6R+QhlIZsbqKw4M/DCQhkB5i+jyXHw9VMPG3wwfzi7nm7R+UM
i0HlRz0gdHajviK2OxjkVLnbnLJxxHhb5H+NpgceBCH1lcpFPcUMZuUd0tU5ftKBilgSM9JHy/AM
KUsB4UMMNBw1kApSHZ1KrfOR2caZTDjsmeZkdcDtSdYIT41KW7Aa33yoZbg4CbiULEpFtPiP83rp
ETGBz01n0NAuM9GJlLfFgicIZM7cxYjknwCSiFCtjQ4LtPIFJQgXRgE+eWQXqILJIjQ3ZB8+24ly
ZuIenAv2h8sXuJR81SJtaEDHHU5YBeFv2m/OEfxDLQz8US33LdVNegupg8y7a78RmfgJN9EDuWOz
aFK2BdPAo1VOp/9lUp3kDgC/+slMMFTZSRfOH4sSzex4SNlSFQ4fbqDzdxLrSr8xGwnn9VeHZ2EW
fUIZoxeHVo6rqPE0UK2uegDaowExUI9Bg+tuePAhHaIuGwHCDDdlYKTanTvxXX0NBwk8kXVGznLQ
p0yyyyEQ15mqPdND4D44dHJKWsr5/044JOmfqDLWsM99IiyAd0pZbgdQbYLo/Jm/dOSsCZmedH2X
5us7U8JjLMLkPuTWU7dzs0qFdmdmh8G53OsLwYFRmaddXM78jV+jQxb3HvCQqisTmPSj9vhbtiMI
WFs9VK3jRaKoimfz1WY0Ju9Ytqjmer1yx+V7eDsQi8CTOxk3DvH4oinNrDH47jOxMI86wNyzkCBn
mvVs3RydAR0qwwTSQHne2A4klZ7k6MYQA4wsnrfhL30Kptvpd/a5SQva9RU9/DPea+3P0dcsB73j
FOke7j3B25z9FgSUMryMLHyslK/sbSp0f5dcMTM/hyWlGXhoA4K0Tqnb3t8f8vDIEtbTuHZpaA+5
4MDT4EvQ9mhrOHcVbvtoJV591I/WkD45Gh/q8Dw237MSfZuI5DqpNJuERqJ8PkdpMdFcxA/3IsUl
peoc3rrfM/3Co+ZZIcvTdIXU35qc5J3PQoZ0JiZQoqGAUlOSSHzT+PZEIJm9/4oIPuzrOPHU4q2l
yVB42VPSPqazfGuPppkRF4ZDbmQRyVn6eIi1u10dkWYhSwqHG7+/0enHhBLh5ngASkdGlX7YqNbT
UQymDXJT0LAQyRzXA2U6OL65B4yQ1F67ZxrWtCwlSNopr8t7hXF9karj388h40aC313lNRehtpk1
op2unFbOCaRasdPCTIlxCzDha44klJZONDN7ARVtGnI+2X+2PaJCJpwtulvSzyq+RWPzgt8qTE8U
z0A2zt5sVwd1vzrUPzTkWEhIimtw7BwhOCpz1PtWtXQr/0g21rDLww8VCjToHV/5FCWJZSPSG7gf
m99YKPS6ihDgoSfRDimuURM5Di6OVCATWApSNKcgZijyArRR43wBPcMx6dNxl8t3l+Yst6SvG07e
VR6CBLjEaQ3vraUXFFhLsryejQsvjo+M2t7qBpbt/WALoJmRx2Hi0L9nxMfVJm6AW0fk1AzHnyMF
J0uozumrY6ixdl2XWUrrg6OWY9uvLRfqAKo2bKC31urnmDLsHsL+Ojf39oHm7X385bD7ltI9o5yI
xJSzNBxyroKGThv8J6YFgI/dujsLUWy7gXTcr4FCrazktdVM8qMZhdn39Agsc6GAxALzeBtDn7Ju
rNYKCb/I6mAXaIDX7T4+omcf9V5FjfhtW5seoZ8/gZy1Q3oIiSX2WbmZISoUB+wD0pFAYVIbqlko
92MM+Y3kmDmgM6aiQZPSdDTI/jGdhAHGz/TdSpZHtVHN6p9OvXkcbzh03tisMLxDGDfEtZOiPjQO
U5nRynwojOrSoDJnXHkrQGOn49wIxP1vQx6ML7B+Zp9td8aTa/x6jhAuQsS0eM2y9zY8fpeDciUm
6eEmAU5lM62cyav2lgBRnNnv3AQtNttNutokpnmjvfo0cUzsTRc7GokIWQHtSRwB1sqUw+Kgt7ym
Kxf2gJENrR4QF0KS4RSaLGPmCu4wGApHNkRQX1la7cWdcDZ3xlhuNtzwfoN0hGAhuePYh/ywqDRq
ZAFHuhlzbFAFfy3NYG6825SYDu6F1mocOpc77ubd5cgT53BIybV+B9r1uPMen30aD2s7r5Gw8YPZ
BgEwC5SDGR1PlZ/qvuVRae/ddrM/DOFtepPHhIG+XDhN+THv4Bmnf+gxWMQ4JhF6F9Hn6ru+L86c
iqGxJ1fBOPCKisQvZEGw944OKMsBh/obpsxbU/eFfY+/G6ngR4aVEUcLBPxGCkbpnmq7mhmRnM/E
uuD1uTJwkR+FVorvkz/ft/EckDgcUgtw39vh7tJ2YKKKBHKbNefNPg47qhK8vM2swJEsgG54MBDn
ainJeK/n0IzqfDz4Ehv3sKFRbY7icRSPOuEHBdxdm95UicAGnUlXQGibFhO4pZp4ilf9bxGLjfOf
Rs2IsB7alymtzJbnCOb49kLb3VIuyifcRxDprydnj9u5EFFj0PJhZamv5h1cMnz8tllzbSbu85PF
Ir+yNOsnxYOPk1j0rqZJMjGaC50mKXaJYBvETgJqrNEIWWR27QMl6jYaput4747O6h/XLY8ry1eG
UvmaIvFV2a9lzCm4fcbzn+VRQUPHTMhBKEi5HeIiqgHVnd6GwpO8F9zD4mwIeGUFV8Xei6CDHjr/
Zmd1dKr6zm9UHdrg0DwmN/t85k+hH0Fw4tppE2UQNnJgEOpGmLzyIoDcD3oVnJA4kOXGMYuKXqUC
wIxrYU5ELJOPFRAOMgclRz+BU59DxMXVo/l18A6wCdZxfdhDmEfUXqwSwKQrxrWpqws2+3VC2yo6
606n8jao3rdPH/RdgL59ziMo0oTMASdsp2kFHd984L7Cj6VZa/qIaKThFuLquaGVfAvaJ+TQQcwo
IU/6Uu3X8ovZeVx33m+VQrVD+6EsnBup/4FR/txUxH2JUuWphD2hXgcnw5u1KIJL2tMKQcgTHNUH
rhln3bgKBRiZL0/61/Pfu3uxiim+ThKHbP/pqc8xu3rcpnxNvsfLKjtxiYU2CvwBT9z4D88CkeM8
xuQTenMxdL3tmQaBZpjn0ovJsm4qdttEJv6KlBtuLh2spDCmHYKMroGXjqEYk5M7Axrpev7vtZF1
LiAMWzI8NpXJdIeUTIemB13XpJ8yn1TuQ+HBk2/6UrJywdSkavqtpsYCa6olHEpZ8u1PG7MHgrV7
vA4vHGR3jvDISVdRFq5XA9X4Pi6/gm6byLv1dty9li1ytinh8s6SAXaBNEMF/VJUZvRvIemU6ZvI
8SjcuOdZPWBVFIPXKhZI92E0jVGAwR/cimcTNhM8beNbu4kIju6HLZEqH9WbvnIVHqu5/ARHp+4Q
oC2Xk/8ckIa1EkqEOctmf/oyELQPT4Zjf3DpSQoGLGmDDoieRASiW8VhdwJyk5kZZ13UECuu6ne1
swCnxk3nt//8pvcrBZzvIiAH+2Fc56I/MD7yP039mOxSmscv7oWO5SwUB5oZBnA/x3dE3R3cqG3d
TwewweKCRTwTbnQZaLE0vFfNjb0xXryw4tk3yJDluxiHxPpbsLrXI9HV0/XNx7rzKr+BCnEBfHUI
0IOLoAfl7ShICXjWoUvuRZXrclFBVSN7ucCdYtA09Vh3wN64hxjyrbA5+hOYDbgnt4EPNqEAgp6/
OLOj5daJvLxXYDkVWf/5xYzWTW9YbO/s46M+GxjGXa29cRCjE4cIJ/AcqGNGxXrUGdorBZ+NORy6
7sN+2+qGPgUMzHqePqSae1IWc/Xft//+jqWjmpj9Sv42mZixmn4LvtdCqW6NzX3MmxKw0WV1Me/O
nlmPi8mh5XahVNp0VN+xJw3Vbyg1fANRZHpJhe2ngWwzsnpWFJ9TLuLR9F+4lhh/DjYlcJa/dyui
ue5nFFfZZU8mLoXICd0L4hjOvhSvXuumdoe8BgwYTtMLSxnIIsoMELN7Qf693CUhxCUTCvoLctzy
ILdgCqxQBP9IE9OTi+PoE6wqXauGllmdKoMC++CadVKHUCTMa0du7r7yshwGWdPUYq+/nUUDXwQC
dsrOqtY/Ap0Do2vEk3lUPvlimQTPVjonISYNpJwL4z8PkfAJpucUj8Tvlxzue/bnC3oRWDmlykj9
pq1YL5duOAojXg6TLMR1pocF9SjYCH9uGaYpv7wncm0bQqWWxeyTUiuXxuQ1ITDMUkjF/43uptla
HnyyO/gbTtDl7UMWisQ0jWlHi0JT/At+D3g4HGGq/Fpsf8INfAM5J2ms+nUXIf24UypYON/Q4FIg
0cRYpY/3WvoD2tUYllW+0tAamgzdurukGr2QOPKRIvo0EufHkYmjx5BhSUsnsSpAqJEIfB0UP9kx
1sm+himSNrydCpmMhGzEL7urTu9DDp/kpnG9Cyj6ZVHvOVfHwM5FhGD+ba1CVX411je6Nf4vQRRr
MyA6E0pSp9VhNR3kA3RWE6aUxIfUe1hLvDHvgE19uBPfrMI9TERvwvpRdGmMMd6cnQ+frwCzS2T2
5T8gla8/g8IpRYAO/zjrYTXEhIw+O7PRhcIO5RbcQjOXbeMlB2OXPcT5X0l8AvLTcGnsBiStNmo5
O/nQaOJzjl3d9pfmnD+kiIGQmHFEZmJ/8rnFQpLpmZBAKFPeatKCMpelmWg40BEdYY1JVWjumVsW
5Y2Rf5Us9bE4kUSN4LrBN6g4pfvKlGtzQpvptmaFbvVKj0arxsKXVX3C4dEwRSA+QW5/V7/pUpcH
0BTBgMFNiL+R8l+i559Rr0higJc8GqWJ0fCfG5zbqsKjhEXROzk+qrMZiMTlf2WWbUdjDLkjK8OL
cNOU/Z5/L2l/B62XiOEEHc/sCIGVzHg81NB30opAMkKZazNP5yNrFUvvbpcwvIAh2GzhbcQwpzlN
rGDyKAks8Xc7aBWZLerDJCASQfoq84yANWEoFdG6NgZBqojyMnIKi7eNJD/EbabHzUOPMjTAAwuw
LqeT16N0iGc/CYJnHLJHWiiz6yVXLFfXmSIQcWNpwiJQ9L0sT5TuJSWDXLpZFeJyORpeHMglSmwU
xgtFBb0ZLJdOlWGgNX9YJtKRnk8DGv0EJnotiMprN91MKHoMUj/0GkvrBhClxyRghzIj1ngxlmVD
klfJ/1ZM+uLKyxvX3EYD4sRs3CwriV0Vb0XH/r4lShzcXqChg/NcEUxFnGudKyxNK+lFyMl8Jcuw
iOdv/TE0I9JWw/pxTQIiTBFFIj+tM0OBLa3gOKlddfyvEcgUH3XAWg6o/qmn6Dek0LYcKeQpwOlg
V5QPSi6b5vv6SAyKlrz96eMwgim1ZQ2UdIfIc4BQn0YqmoIFQIN36kRqhaRYpXnbiW1l60rpR8Tb
tu4RlticIbKWWd9nlruJaqWPb5JU3ZeJ/dmwHS8ZMnWUSH1YfjB5cTrocLc7MRSu11ySWAer7puj
DA1LD+ZsV8zhzMB/euZD43HSuqUdsb9b1OtmRJDOsj4yvcnTSJtt/JePHq4qEAlNpTdl6nZLCcZS
HDsV0pfS/JUWuJywLO9J5a0y4GNIuSVGQqyc319IfbFO80NH0qI+RYQTt8KaOW/X4FvGf7Xoiptw
SegMIyZDBKFtPBiKdXh+Hec51iLVO5fsUrjs0lI7uaqIDc5G/0/hJrSmLCeqQSISVG5SuOBPA4SY
S+d73QkCJmI+nxbnOP9iTgSNiJU9QX4O+XsDfbUQI3eUv8pTH0TW7xxx2zu5IweX+pLq50AXgx96
jobp/hIA9F4m/FxKMQRAGKVZCxsuPSh18pNZWqtbm9IRVn6Pqo+/oTnCYbjh3xXkc2XYFIez0xIH
x3sxlNO2RV6XbWLJ1eREw4BpVNteh2E8f3XRr2kW/M6mh5zGEQLfkSBt5906LeoAE/CAMkh8NxES
JASA2N3GFga1zsLxkUeFQ9+28s5OHtfh98llIlGUNkOt6HaaAHM1OZiJYIAZa0Xyukeb1Cctjs2R
jwpXO10K0StbipRCX5Bh+FS2fEB7y9o60fGMEqee1GT0KMxxrqWe+j1kxiv5S+uVfEOXbY1xIGpI
wIrpBWVqOtALO8+4UzoASlpo+b+LEHorko3LtDxkbZZo13RVSIXWzq34a4GSBNRLhnvzyaDrubdk
P3u+wGrcngPHNZkxA62Snw4KD3uQZgPE9JLAgykFXeme80iP/K72eAhD+68w0f686wPuH8hbExqw
4DDsiCs53iwobPTKI6Otx8WXWG/V/qHRJr06Q7hfrL7hYBnuM2YDZ1cNYGG/V0I1tlScpOf312EJ
AiC5wlej2Xe/HWmCoXDIVFf2r0JgpDRv4qRQZUwdT9W4tY/JLcOGVLIAi82wfV70Ph3Rca1uDRXB
XDRedsXiD5T1NLnNqeNvK/Pr+kSZn0OXZYGVtE7X2y/KgCAeet6iD9sIFlGX47Z1vFysW2qbg6+J
kNypMKnDijBq0QNxCV8xKogak01Ab/K8DQp53iDkakouai3PS7OscBGazRcqZ3iQE2ZlewuAnxAW
hg1G8uOeevxzNvZBsDkVZOkRWryFTASnq/dkTizd6Mc78MxJHICwFysCToLC/G7gNQ4kJ0Tl5gGG
3wnXnEeD//kmnxkuyrNL72L6FtNocew74DrSxZm2vCvBTBAGCzA2HeHK7MMVPBM4UI8Z+0kwkGLq
buAd1OmTZ5+8A7BsgjiXiMgqoPJu2MfCLslLgsxqIA8wY5y1434OmMnFYuO7vn7Hc5ghWcMzPjEg
jLHEgtDiaDoRp0jPDE0bGDrMYpZySj1Y3TQVeNL4t3pitWdR0QKnyU9t9krrwoTudbAQfxh+Rp9h
T4gSAEXCV1eUbS557ALMsrfyT4UZVCApcFvVvw+VC06G535luQ0ERON9z0P4jHGWC7dODiEpX3cC
Z6+am0HCqCqniGwwa8EvapQwsX8xFgr+FWDHesaESw+2L4bxUuv98yAAdclQHLG6fwtytDGoRx1u
xr7KYIjnpf3Te8FLFDANcQjKFQvnu5MEvIkGouYaSLeIL/wJTnU98Nh2JTDKfLMXbXvEw47MyX9P
dWAZinY0vQ5K5GkCbXcDqmAB/7mh56UKckPDkx0uD1BqUfTu7O24GWwYWXAmhyTqWSA6Emrkedfw
zJ9cDJVGetf1d0xCpmT1Bim9L0Ph2eUGsFoySQxPSq8eTcRKgsZEjttOvs0GaPuCOUuWE5YJkWL8
ZNHtHPTYQJiS/7gsK0VzryQ8ppksu2IUXvLqsIj9jXmT4jsC0RAomV3B235YsZ5fKgEbZSUs2ul+
6j51HgqewWh472/RniUQTNAYZwgsVU99PjE0St/r8ZMZwnlHVyJ3Nlqw3HAEPvT5cpDmO9NQadeD
q/rUFzwf7rs9j/Ajr6ZJ+KyaBc/e88419RsF+g9OGES0LaATMOiAWtoMirrtSrER2cRcTGQ6aQ+k
RCHipkVJfpjnggidmRbRvjJ8qvzNmSBI9HNLeimnLvGXD6majVRP2gw1pLJlgHJDNch2z//aOzDo
VGKAHrTIul0FqRS5rq/0HO5TWsA0aDRVVXqorTXe1nuAErBe2kGSDlINSn4D917ZS7i2INyrzjzv
g8cnLvPVIQ0IwrYiT1pGN261zOGt5OevXpMW/EkrF1Yb3ZFG7kAkFvVgkl7xou2gcmC37q+qLVwe
DvsMegFsVVS8+59Gy2if6PQ9AHcyQuGuFH4yvERxjPHCHvZYDcRyEsP10VMWf9dIwijOtj4TwtMa
ZgwLXQ9Jvk19j2Mh+pww8jHXz7tbb4cZFeLGRzmgCfZOj4XQQ5brAqQDGe/W3pPb9XHfCJUvQrnt
mQjFS1+8EJKqnX0rrgwA5V+2DbIVWxn/Gvkpfe7XR6D+9oHFWfAQYKuKuPs96aHeO/w542+6NiU6
GJtDxQ2GXAv6p8jmpzyOCGpTwjFBB7cpaxhE078kBJd5Ph1mHn7eRPWCyXDmxsnOggYdTu0MYJ6s
587hnU36vzN2NTZX+vnXBamFKWfgKBzRfXctHUu0DaJJX/yULfGXfCPqnzEeJrs+cVFQAPJ/SzvO
razR4oMFQoOpjMO7gtzfB8loOBLFIk9frAuCjcZqnCWDIkk2kee72NO/o8mHI4Lw9pFMnsmYyhxy
Y4JLEUj6y/wI7lfTiPAlR49NM8i34CPrAl38kXKHgTQxFOqRjyfvtEsw6TYRGwCMXGYFfmRNnVKM
Go6FC4iv1sWFknso8mYcUbqMpAkaRCXCR0WM/5P/y044QwKvluAKjXgbDdWTLHr2AwEo5a7/dfMw
meYAkn+4KYGW12LtAJv+Xb5/8vugMKsyIxovSQ/SL+hqQx/kSPkd8IQ6GwQ7IqM+E9CcICMwEYgY
6gfIqVNYJ/k3okfkz9G14Vhn8VvA4CEqoXysz1df+vYVbZSDhuwQ6C0IfZVdi54GLyIR7BBAiq8U
5f7hFXOi4/UMCqHTM9C1vHZqVVCNbTs328eQLKyenUWOWKghCr6B/OF046FTJ8xpxZC5kNPkVoYd
KlbKB8aBxI5NYp2vyr63jEw3IKbpvPfYfb1eL3aLzk8IRPiOSQwh1IavitlbTI5AML3p39YOwEHg
AWyXzthJB394ClczXcgQtA1L/V0ujaR6Tzrf3g512rThe6seR+VbLXql1s49FY4Mc/C9lg4WfQ2T
RWKjMDaL4KLjqUNM9dvd5alIir+b/YS70YspGl3f2FO0TWWXrB6F6PNcYrnOreze7yikqPBjRLDy
UfiVnKRcRs2czGmEzEcdV/c5UW9i6tNo3DVLgrGY0U00toQdp/ykDmSTspNBMYM0XpysAj25PPeS
oz7ax8mj+78HBj5T7s9nPD/kUUlOc8n6NFgcQaSiUknDL3EU/t2750sttK+/JwMgL5uds+YrEl59
/BbHfh9r8MN4Q3KvLVjlfXadHX8W9mAq2uQD4b0d41R6+Vs+qfTRnbGAS0ZkvH+cuyxkjZSJUChz
39fO1597elCJNF9bnTz7rae/fZGqKQlJ9lYfBJbOs/4NL8gIp+HcKFsbRkBBgBFlkmOecUx9ewGM
DGKEBPpQrxt3ear1GrAhkgj6AU040MTtDOLbZw0O5NJOOfNC8kcLrsfn2GC8d4pOxlru1Au32gqZ
z94MM+OWNG44EwQJ81Z/DTw9BK4iju5ieO0nnnkRipKqKXm1MWsjoYooz6JWwR/ex7Hfgu6WFwvl
FLIXIjnqmTLr4FX+7jhfCiZEpIVWtxRpObYZV6BUpT23S3cEYMIZEIPYyTW+y2zd7Wuwj6n6U8AI
Se3xGZfNVviVGkmHOZJCB1Of9cLc3LAXuo1bdjDjVE9DBuknRuEvjDpurllqVdPPaCDVfdr8/hU0
H/58lxy1CkUcp1cl7lP/Nx1soPctgiDlQS9+D4lI4Cz0TuyBs502Y8414o6Jo0MUBc0yuRGGJss7
EgcWuaZG0NIVonWP7mKh4vbUm0qVAhPINQJLed7v/Zh19c31mGorqOPgJ+2dZwcLd401vZpkb/XM
jdfWDJrlZDcgp7ZBiMFnDj3Iz3bgpChywD0ocuus7AHmd6vJvwc1GqLcQUcaGvncmbm9s3HC0OgR
3fB/JoiZEgiKsgDZj+epoDzYoX1gw06YjrmGfZSr+eOUdeUFGdnG4Nx4yo+lvIpoaMMnrqyK1pmP
dBG+jqF/ZdqmM4OzjK9C3aPpXkSJ09yrFMgtsQXO9AvXuX2qkBgeFf5DIIAn3DbrvsuIFNjflDbW
SXyZ4ciKjPoSIaKSzKXv4T/RMdn5e160DRd/CUF6AaGzT/4uiajLfBpDg+PL6aXOe6FgdZgdmPZP
wHIVGk9ktrQNP31d4vUlvPkLc1jxJTjgicVVq1u/pE9dvFJGpPOIQdsnzIV8TJphCaGobxlHsYf1
MskR9xPwpVylY9Mb8/VZjd5Z9Ubh4MhcYehN5UzprU8/OcslEmjN5d3u6+8duz65SIGGpGyvqLBT
iOVqmSvjWSs7qY6NaVU3AdRFwKl6vF+Ax9pY9SFdEnUYj2EUY3VV5Z6ytpRClZZxcqSZtcJSFEJU
DXrxOXddL2wADVhHST8GHXxf4BhBwlL/EksbqzviCuoAhfFFl9ZLyCLipv3UeVYLz/3rgXxYFCX+
PoCIEiE5WPNC3lEDFyIyAwsOQEOYpJ8BwcmGXBwDcSymZvHmtnp5s4dex4o7wcHMq2bjeahU1UDe
kXXVESPWqJt/GUMWyOdQ84E1Hf+2wtNNcGauvFA15SezyhY0IozqGkm94LKtFw+IzI1p4J0Svw8r
ljjfYsxnQWpnkcG6EJ9ERH/bAqG71n3oMHFgcFpnGpg7BEbIbyzUuvsoA8x9lI1TKiXKiVxExROa
SuKoIs13uVkRAEt7qq7kJWacJhULilyBmQn+NJQRwMHVTMSp7fSIn+sEYGTuwoFIyOJjrMRWVtTA
F3bYbH7FV0qUwkMhpyUCXJ1EP0glo+dlXpwtLvFId0dLd1RvZgDiyr/P82ashQKo/USetrNe3shn
9U0FqAI2A4YLcLaQ/+uXPhByzXlbcU3w2RBcOFkNMHYvDCAI/lqU+fmXlE0g/gp9aZuaGQRUiPTZ
LIC/pCsN2L+WHEhwFmQR+O+LSmQJDxSZmENa/YjepkCSOR46BUm1G4OY2KrRPv7o3+qSwwowZPUr
I9ApnuY/AFKCHbp014X7XQxwP82ea3mieLReSgXlokrZn/sbgmkBMDRv92VBI39vUBx9oBij5dWq
8vAoGptWYueuS/KhJ6ypEXzv7V4YNIbk+8ZOx1Fw41j1V3gSIG6zACEpmvt0llF8u4SThJT4h559
abwWHPlvTriU28J51P+lvFp2s3O1fuoHBG/87mmxK+ivT4UTPrwGuutrTrLpPNxXenlJ6tSVV9ao
mNpZyqUny2bWG2DyWeYMET06XTqZ86da84zWPjrxolMPdVG6ZbUgQ1+wy0zCBCn3AGZRmINKJ5iM
V+5DExvgqTvGPB3gTX06fbmdEP1bwCHARdlVWzKzEjNV35lCr6MLnF4QSqh4BmD8fur28ygxRnDB
Rd6DSRtbqe9KApPUDD/qND2ih13AWFYOS07KbJx3t2zfZVn73A1UwgSS6nZoaH14Hql26V++2zO4
jdOhWv1i8Q71J3l5HPROZP3w8A0cuhZ3vHQ78Xv1nnYTllg/CgoUqzzXtfD4m2+oh/VtHU1lNe8l
1Cc+tdvd4y4e06EIqeKM/xrZb3hddE7nsIAy53wWEygX6oiomL8+CNlm6vPUZBzf+m8hAYaLjwfP
VwFVfr6nXFubO3tDbAva3MZHgSWx9BaIYKZJJM4JJlXGd8BYJRJNzcNleC6qzDYLr+dnJGMsz8+P
571MRjoEHtFCquooGhjS0iI96SuIPdZNOoDV60oSrdgbd9xmcHKkaH7Jmaw1g+F47HEauQ2xLq0l
dUbnMpUFnoCy9W9yrF/+uhLG93t5qvlx2gh0Hr+ZSrgE+eNulvjPiMgTSHKMilUp6osYyPySepKx
86HNfCsMhzAvVLTnTV2W3pnaEgqpSsGjoWbyx6F0nR4tmiAEW79yJK2+z/btButKyvGfJS49+pnk
1h5aLLCcemJFbWCR7hS4mqAjPtewDVu+s2NFqd8mnTMi8FZsq3c/QlaQCg3LkK24N8XUanpInhBp
n7PiLDh8UoV0KaYPSof5yR3mjJyiSKRK9gFXg61zsPnx5Gq9FVHD4t4zJFBBXMH9rHVsuv6y1tKB
V3woboEb/Palw21eymwEpWqdyHqTbHCPCXq+o2npxX0IDvKHhO5YVtTdii86kFtZzTymwx0CgwXj
9ECq54pIaGzySFgOKz5r9EYLETNLlhBwNhaKKiAzCOkNACXSGi5OHNPRPQ3JZ94C43PuJ8ktFxsX
vo7xvKb9cr9f/V46Amq+rBPJjMhRpDeg01rG2euaUrtGPjEvFW9DtlzmeD65mBA8ih+MdnLQJ+Ds
7IXaN9NkXHXznP/xrP+hJJoFSV0DugbudbbpAh9ygklFIzibuqKloEm0vj7fI0uMswyKECckaUky
Wjut/6i2VUAGv2Hsz9bz/CZX4TUpxQ3hiBR0Zr9CGcqXsoJ9uhZq3VpHFEBZnT2FHlJL+ClpkEu6
AVT0LIJ9rv1CxYRYBLHHL47UE8x3raBYn7oifkj7JpERHFKLKJZzJr6Vqc3PjAIlEaIiNpmLuLC5
ePRmOEa0Svfns256mHZbl94/aPgYBn4H4YcnZprRKyum05qoTCVjF9rFXBFq8X2exV3msfCgTPAd
LSFA48zLDV57VcdNBkxDy9M/66ixpKNi5m5e6qqV3vfdtAkkqf7h6dqIx6sNWCxXdyIQ6xVdo3u5
9s3XhZge/hgd1tQjbFzw2ofdFGuMFSrEcViTYIJW66rMwR01o+E8/8H2vsXyOdRauRU7K5bThYnB
gVgnSAdi4q12QOX3AIghF5WLgXsKK/DfmC3+HXXtAi+RojX2ANBiHDugKrFACAVDqNRuGXHSJfuq
L+Q3f4gfDXNsdHIkz0q3MNltSPBbB23gTq4eEiHhktPpc3gonapIAzNJE4EtxLrXQa6EtXvKToJU
0zky8upccZaikoJTGojpWfwizc4/riaPaanybMUIqY5s9BCfhLFNXNaNbPYv34CP2BXqvI7nJZLs
mx4d1rtWFRTbt5UR9j5bZd9IXVb5w8ciDV/yMnnD3va1vXJ75fdUEGgczv8nw3d/XT+n6VfoERde
df6Oy2EpxJiWEhXw068EOk6SrVXcTXQg1NUAoZTyNFD4Jk74+8DLzMFnphGrAhz9anZzaluQ8w/g
jfYezhcu191g9HvyqLZkfKRRmPHHnNaCsSoCCAkKd2hTUhDGhZrzmN8MtsmP+caSNn94HODf7fZd
ikGrHwIaHf8YcMSwbJqNaKRCbmpBaNi9DfK9DlSbmkEOqmUokfTrqsxiM7/m/MP+zXM7ma6BfPBa
Si9uhO5Cx3m2wJ9KdRI5kzUlA0++nrf7TGc0bRSdrR3M0vhuf22yHBazmYS7bORNAgnkLTmeMYBG
Flt9XvjxbtHN+XqyYcmSdqEAZKcezc3xSCM/GuNCPAZJ3kN+HVf8uZVEc2xDGPQSL/K9Q3padqLm
gwnRsiMqAxOssr4RWF5zg8C0rp8GmvL/FQcZzWwv0gWHnLC9l2bFvDVvNx5bKPY6logr17wtyeen
2WUnT0wGG3KErMFXfB1ylHF0SJFCDBIRKR1dFGMV55ecuLmD9kWK3E4U6OgVIYD+rcWpOCOc1X4X
/L3DO6z5ogytLdlgwT3IaO7Mvtnpzir2dIGTaTHD6ETS1ATcxcLEB0YU6mG1eJJFFTbNAPN8nZSs
x5fqXjSBGyL3bqPz3C4ZA+8iqC/BEe0ABx/cHZKADdt9r0ImYAbjBhdT/J3WyBYsd0yEKqCO1iMy
zUN14JnGMr3TVvOWn03iWbIyHLfj6w+hWVCLSHusEnwguBFuwdWeyXgBVz8SvUJIUvrGtRa7uGUy
vJeDQk58Crz9LP6zHcZgoCi+ru1SDnBRBhbU4riP4DsUIqFiXPNq1TCaOUYtc1WVBd8Q89/zvyr/
ILrN2aFiLTmokFsnSjF4CncxjMITZXR8bRM2ibj65IQvga0my8KeR8qXj+xnum8MS2qQ66/wZhd2
vJ/1FLAsgJjUiC0RIynE9JKIGLPHAaTjzx1WzcKPr6G8VBrN/iGNHioog8orYVxmg9MDrWb8A5cu
6vf17akv4MI1H7zADlz+H72ruYDIqdWtLSqQo5FshjCAGdEYw5jTJoG0+wqXJVAdRMdEzZZOob6U
ovJOYVkYxFZqoAMAvDVcTHHlyJLi31C+NSXmFsyPRcf7xHVo8E1g9KXsuOC92RrdUlKuOCpI9ovu
D1rUlkALyJFbMZPxk71zik/1FKx8Ve1KyuG9ZB6y/dXfrfvGy5Y1U09bVCwBGIFpMe4nl/jHhK6o
pWkKDjEFmZx+Tcp17QtEnJePvQYuWwdgNcqCLkWmzpYZrsX4pANm95E7+76Q/e4Z4fmxX0v0K82Z
MOHjjGt0MN5m56xnLxCa+oq0O9lFyajEADBk67FPeN+2J3TuTh6N5tK26nVu5Hjwyzi5YzoCaowr
GrXBpehmeOt6f+yqaZ54FeQITSUC/Ux1tJtWvaUprz/1it56nWABUj/MjXy46CS7hPtoCgzxRwFy
fpgLk0ScSO+xkS/xpuIp7nm94ACbsOLWnZHuKTMXy3GC0af5HvTme/D9X+rpA+G5V1vVK5Me5r9L
vGBUAq7AgGQAVUHTfyQlcPkTPPLys4UgREeafbMMgkl7TqNFTdIs2odz+k4im4qsRJf85D3MUL3+
oxWK3Q2UngMC/Kxi3XvMT6wQfmLmrTvC14n4u71ta8iWPeR76NJKC6yySwrY2KMJ2ywa4AHOhRY2
z/b10IeJnXfGlYpT/NmmAPNhGL/Q45jjUKKXEsaO12twkp4FgiAxITDYiu0ZJmTYY+POpcU7molE
kA+6TMOOT7pPGHe6B+BqszZE033sBz4yCMziV3bASC+iBIh4GCelBsnQnj8cWYytkNuZI0QrkQld
BrpQGg/pKIRt3xMpXaf6KzLKUlnxS5Rod4+lGftDKMThUGu9LEgFXnfIdGtWWtySmmdouED22+nH
UaESg/2mBP+IhEEwnYW8zJc7d3bssNQzT/gLyU71x4y4TAjc2eM+HXOQorKg8lTAV+hFcZGKvvyM
1rVa5qP6mnUm8GL0bBpdG2N0HRrPd8i1nZsJSZBZUDyFgpGEM+p9rj2GJ8JWxq8G2A7Guhprw5sL
H25vSLNNsmoNOg+jRMqG+1tPIumdpUCFz+9D2DGK3mmmj0bguyuhlJpdm8vR2zWsnYmshEgYKHbX
+BZGnrNAgL/K5sZooBHy6Fz6bY9A5psnTpJqlLuUkhes9s6uVJSdIYbn9inRn8kNKRhcYHad26Ld
Eigna5hGMIwkbVSfhM3SCaS6Qu4beOIWz+i2jnJV1p52Sq8YY6nSdVCekUceGWITB40RTo1DpOJu
471fxgYqAEPCBUsdHvsJU/JV1czzLEYXrlqcWiJHNW+Ao2T49hgmJ03mfVIB1OudOqZnyy1RPpgp
BPZtT7/TuSJGw7HDAtuWdoJG6AIcapltz6jL6u0QkVxVJh8O7/dXo2vaMGoPzDIOEtvcrJG5Wbj6
SCc8AloHlEC+gf1kIoU8Lb2XN1W+I/sxf/U2TyFKSZRwhbXX02nVFt4Dd5bkP+lqrUz0ri5PPAG9
6QOuzZ+C8qwB3Q7e0ViBwYmyKHwttcb3cZ+cga5mSs4qy+IO2u+YYVTw/OP7ZwB8sqg8BS5HvyV6
yQHMAXEvCeKdevOUO8c4EoeDulJAeghgE7voaWmInl1F6CirfGqVdlJ8zfQtkFehfb88Kkhj95Fu
omVzeFpYjEGQyxqYSAIirW11y5O6zCvzFX5gXnAOygMhynRVYx1EZpCKwJqr9N7aZAWCJ+mVMJCJ
26pJzOUt4j5JQE+STnpl90I2qKt4f9ZoHgI6P0gmFFRVOi1KyNTysTbVnNkNwmKNiiLo6PG/z6sH
actFPLieT0U1ajdzTXlEUOI6eINh2YJdzcfYSkIW8Lm8DUZUcY1tjtNr1QHTGoIst3rZ/2qaK5pk
o1BHsC3D+YdumJj1xubJV16wyebYMz/gOHvyOb6SWw6cP10qMzGj+mjNEWazfsQdGlzGGQ72vlAz
P5EMVcnLHl64FAFVK6OBxhs0awDEoSrUAt15V1rev1aLMYIaUYnb2dsbBTv6gzmMuPd12MRUA6Se
AvQtRx/Cgi1eil/oY1uxnvSatOEdI07+3lgAqQ7dVmgHIgIij+/BwjIQCnTDqTKo6tg+E0mEL0mQ
nj82k4qyp4d8c2Og0rwes7tlQjQ35IuSg9UU7KDSsAx6cjY2tDyIT+ghvIKh+7X85AMsylOh+Vmd
gQDpwyWeCnQPukq9tUcUVcpqAJ/JvxB9xW8+PBYmUEM8NLlAL+BIHbRrUhWD1oQTP8qKDDunM7aC
QaWPKpZlMdq2EW/fn/TIUHTxQkGeXcBMORTg17TQ9IjkmkY488IwYePfSZeQ/XunwLa0yB1t4YYH
Flgz2tk6qfaQE/rEPEIrVNTqavZc5ay6zDXSDCycYh8PDolGMBuHQHKvL4tg+5AcsIJYMmOIcRnE
qyd3m5ovU7kAhLoL/iNmjQhUeQ0EXCm8ccaM3Bh6S0C3KLUr1KLJUgTuTrBBIjgYaA85QpKR/UZ3
4eaw97kROhvpek++CTlRnmv0E/XpebBpz3lY0yapQCW5OsiVlyt/gttpBMe27dt8kHv8P1eJQ0pn
0HrcavEbsordray6NyPyZpkof7ZxkgzPHkwKAvu/lXJpZWAYU/snBJYXYWrsD360U1uWciYE+Hys
HibHvI61LyksqDvQ8tty0YjxMJsUrOR5/Efzgs/1aQzaJYUM01LY0PzPj+LzVvPRfNgXAJFXiLd/
cOQLHId40l1U8o3za/fsiS9fBvQIBBYQsRtE7HepcdgQljoA4dpbQgq2GwCHQSszrHT+kXTn8AYa
3S3ZTZK4dKC3R1SVawnx8eR++rw20C8Ygk1LPVAgfldqg/HNl1C86F4XzGoFTbsBL7C/EelnSkl9
+yl0iwVDVNr+meBIER7CFYiybqQILVi5qpeIknvsOS3yC3/kGDK3LgU1kXFA0VQh2hg3KfQjLiEv
H5CkWn+CMmoYu7M0Wnq4cYizxDltC90PNS6Lq9cEDQZMlm/Mhf/hTe4oh8EsSUP0d5TCQOS10k9T
JK/WZX6BY0OjTKMs4ELGB58+lpKT8GbKXlL6olMf4SUvY8H9QlYzm+heTjGrJLTI2Wo2kMrHJdmW
7ktcIKYTZZLXXG3mPll6PyKG5/d+bXa9Ya+ChiX7X+LIxYUgr9+qL+1+OAhaBFb6BUg9TWyLayZK
QxvWF7QOnqkAA3ZrwHxj4x3Un9p2N2A3gMeEXCvG/mtWe1fx1QdomrF5rgv2BRpjK0oCitoK+05E
7Xu05Oeidpf9DsKd0+VTW9MlAaREsJJWFMDBMSKNNRJfphgrSVGrFnuYL3MndJR0cCWVsSwniDui
lt8BxyL8YoPbZz1899JNYZ5SKKxX2tUFmZbGOKmSFalDR09/EPRmjNEgukFDl1aMF613RLLIKq17
HBwHbor3oMlqzYZDTTW4a9Qs7LdDrkOUPyIs/YLEZ7Y/ozVZzLOY6xxTyDDdab9hgTH/4AnYrfAW
guxC4fSByFu2THCLU7FgEghK5alyV5x3EHb2Mg+c3gyO7MT0b3mlf69B4LIw0Yifh60Ywqjkj4dO
JDBtqerY54TVEAUSp47ZG3SJUNKpBgwNbcYFEDu/5MEH8fyve8lvLWBILpLEFXIbsRnpc0vzSFPC
reYa1NmGJnoVlmiIYj1B+w0Nz/xkoB+tXGQhLH/b4RaMPl32vBiRSy9iZ7ma6av/AZkEAFtwKuHI
eQehPqyRseaQ+Je1MQAOxA+mWKyPhgKroJIO67uqqZ00iWBFDbMnTqaawr7dHtO12m/QHXaK14/p
T0XWQtwfSdcS5TA+Lwn7li8rRukXEovrKMwl25wC7plA5jf30vFykyqDq7nnQHZGITEv02JOZHzo
vC+ElKuTsGHKuIXlCZPB2C+aZADIJG8NmaKr29/HQnSHRIkqh6/2nGKSNsEGBtOLzsTgUVwjCFEe
sDT1R9CcH9Qul/Ot/tsfiSkOeAHOyO+yHzcxZVjqsXmOsFyQrvXxcIGKPykCkXmCr5wjUzIT0LTu
JsdrQj1OKYS4pEkLDeSfmbA/2jS8m5jtS1VK3y4i5GFb4ANOf5dFIgL5RRMhUFV4FzdLhy+OZurB
2M1QFdyaC7u5s4dMxZvu4pNYDknlTwQPBvtWublfgwCIP4DEXpIZKRUNqStr8DPSAoSzGZhBlO37
lqu2Z3INiKzoBnUjZCmagkpQgIbgKruV1i0iNSH6TXzHWmC3agNxStxNAhFa2dT2TaG3ollTqgj3
bKJNy1VoRQI6z5279aeMnBRff+xdNwCGYf8KA9gUH2Sg1EgHbqyP0FoUAMkhtuCBqJMHXIkh4gwM
nsYol3m7VFF/ubBmw2HAjk7hb8LlpbYjld/e/XCcAeoVxxSsZL8dovlnSIBIsfwAE5ErN4pTEuBR
LE2cT0VCtjyGy40G/GiIAJ1Y1WWTrsEfJ5JykfCsw0p8RgIZKO0Nnmp71U3eIvjkaH0Nk2ryoi0+
weGHEsa3Ovj6ebd+h1BuW9DjxSZmkmEYiazhQZyYIn9488WG05lnFnaGQi27El5YCn5IxOnEAIIp
tF2gGR2MyqkFq5veoRmvQzkXC7v2aZkshD3AD22h/yd4O7bl90aBQT8qdtZEnn6hGHemYG3/hL+G
scLfgXCqWrnrCH78AUugbS0ero1a1+Kgs8TCzPUZKI4x2xPh3c39+BN8rPhq1qJw4HR4No9AchhC
c4Ei2T5wvYsgBNzgajiV99lAoESaYznbKeIxfGjEfXIngXI7ICGKHdy5iRdWfTJGQ3DjlQxO1GX4
4cNNfA1xAnzR6ZE92mPDjCSQWO2ROz+NsNr0JjFRISrT4TyfZuBgGCVpmL4tc7OoSTdGzUmM5Fns
GOmocfnpeC1+9HehLzHiqu2otXWqKpREykdmjjHbKq4AIkWN+XuwK2GSg3uv4DKEfYqjT3KNmGpY
kNVrjrgGXKFaLNuowUX8D4/7+n1/a9y1I2jyPWJSwJ/aYMSI6EPYc5fINTOzT6b7t6eKEU8zC0lr
PnTFGvYf1YBtCP7m7sH6g73IYoLa6doi0Ns0j9PO9sFw6cNcT/mvH7j3yifwv4I2xW2ODMUhZbZx
Y6Lm3Xwn0QWXYF8xQdMVHJ6Iay7ZLDap4paXEeuw6A6/fqVt3rlQAoMD9t6vCi3xZy/OBZuCPLfE
dkguZziPTtZXfo+npmEBSfn7sLtw8woitrCq6DVpvNltOTGUN/lV9e/GuF8jxW2YgnJSk4BUNdnC
ccEUugmd/YUgve1qV9RZimPqQ297Gm495OQ91+JHk4Gr0T1PuYr+mb9BOCTRAF43XjKQMlmqkNS0
0uKSNe83ymCQy2/DCkQWych6mowvXDWFdap91QlVOh+maQfMMYrhbVulazFZdUw324IMtgeaRFel
3mbXH11KugwpnDpiqer7YFc1iuwNay5jO/30udhZksQOke2C6OTqJubAW7YDAWAwcbPiOorjhKet
SJY9+AL+rrWEwMFCZONs+M0/C798AqYbtNiQ0BzdIDOg8Cz1wfvY6o7I1Br4ALYW3YQHuZVdThJ4
FC581pHmRJTEmgS1fjx0D+gesfoA/xzX3Glk8ZfKooDecJn2n+gdI4Y5OzyJRU7/Y1b+rFWLFV9K
gT6SHM1hRF1FBoA8NcnimIbuST7WfB1Ju5unQ/6fsUycktPSsC+KcjEvTvmBLWfYB0o+4xKC4b5u
TyPk0T5Zb9DLKsaliwtQ/cW6x4HcK7okkwWo+QqpGLxJDdOnf+5sNTDa41xQ+w+aohnd84w0oank
LNGzEUW0eKZZSc7xyGlMmP5lcxA/KDWoou8/ycTp3FTCpFLmasaacvotL5NwH9AZgS1W+bH9fuQk
HBDAvBOb8KX7tXtfIMm9FQ3MsDF2mjcB5l6PwChZBqKrJvcq0Xl8VsE6hSUpMen1XQ3LQ4wKqEtB
U3bOTzS3U7hjdZ48JVah5JvvEmXhb27fJskNdm2JUgr5pzTPOuRpCcIA3fcOBQvn+p32VVHLoITX
fDsfDRB7MylofwlKcnryEEBocOmMtTWmS5Bd/2lCUG0cLCrS6KiTopjEUlXi31aMu3OJI5fcbOlr
kPDBryUAUjofxGfMmY/y1uISG0MKDpvARsTxtgI+Rwdsgmywva97PoWkrs1KYtDnNnDGwZGm0peg
/nz+BV/FkuOoUVm7dA8b2RKX9UfouEdLHkFpoysQwhFUTRRfu+kaP6DT9nY/po00hG5qeaGtFgNn
tzCxg620mv64D2QnJkaoIFyY1WvON2AsOodhTI1puMeWxO11xy1mhfcL7iBX9tERd1A0Km/z2LrG
dE0+XVIKM39mAlpH3xT0wczte8RxCWxVBhgIm7LlUUdnDaILEcZ07rfHbhz8Jv1TaNQrDnuVOEF+
yi6nVTNZEHCROctFS+LlT0Kq0oLqX/1jgtPXfspYr+bjLd3x5tuRkJOHCHBumk/TN7FqT78jVIHG
aigNwyrhkaTDQZb+ZNJs68cCBW0DSFk7Kwv4ar0EjcVL8PqG3FudE2g0TAUo2MEd2ZLH1eKVorT/
nP6M7zSxRvMPlowE4ON/9vG7awMrwVe+mqp6dOJ7m/rROMCQNVpD+CcUsSKCyGKQVEvbjJJ+zPyY
AJz1ZaBxWMsdnjknR9zQiE2RectnqnypOTV7/Rr0m+ICJPReGQT3kxATLKB10y4dDWJYHrlE36FS
b8hJ8WaPiZem1Rc6neLATYkYnSENSszJHSCva7DO6GkudHXOdr5xzwBIt2vnsfLGYUQBqOIws0Ks
hAPzcGVPrCEc+Rzs+vnERw4b26asXqgNMA4KnxUwIQ7pLGgnOEC6abQzCIjZruqjkWUj3Xfp3Kai
uy/b8Uwrw6zA3FjYky6G/Pr++ChR69129YgbV3ULiXuZcBm/Sjh3Wyq/6uGnuRqLlwmIdMdSuncm
PIT3ALloQkeyaCs8rMqO2SedOt8h4Hem7GW1YdyFx/MCAB9qpKaDyykRbalfW9lQcKYAINTo/vFL
Nuw3sXT2E4v97Ir53DIQ8NH5ctymgATeIaV7eInOyZR8FLPWLltQ1UrwGxo526RfM+RfOWElDlNG
hx+EdRDzfYeNGPKhuf5NAyzaVVf9HHYWJpNw5PrYvqZ384W7T5zHN1FrjLId8YgQNJfU1EZTxN9a
n2qWRrakdMnHGViWEzAXQt3Ge3CBPhKBRD2rCaIZmL3hy/hmGdyw00bvmtRCyNjGjAowAQdmcJvp
5UXu2jalBiXy62Jc7SFiuM7I1mVgNC83brPLZeelyUKlnxB9lFQ9TBBRs6FYxsoyLqzTQ5vTfhL2
HjmsLq1ii+WCMkBsjlgodJUd0Q7HU02dD6UIneyX3NYqfGeUGMWm2PFle2HK1UEGc88Z8XCQ2IXu
2G566TCHWc+WFvCSosmgSFEUw+3MPLiBKx7HodZdKKXRVoL4GwBywW17o3hO6UkBZlZu4eZQBLko
vIDPCiABXg8qabVTotL4r4eIILwRUzdHgJ6FBPBBjiGsZyAskC2QgrEu0sKxExRJOuHvEUMtXelx
KaGmt4NnGyIqOq4nGO0QuDSv8U+MwGFGK8bUTK0jL72VbdMUSUy1i2nRTTiKAY7Ux5O4Pu+WkQYE
GD5BDGPMIKhx/+Z39TPDtyPc6P4+ugFV2Zf0ZBK/ACl+wyO3t4yIGPxZHQQXNPQwZfRHxUvC3C+o
MFp1lyVerFYxdFSj0ZZo48DPfvKrnIJgV0W+7KImdnOughXvsXweknFyF8o8CDvjqnr3EsPdWnL6
asPSHtXUsxcKdKnTDQ9KytvaJIo+7JlZqGG6JZBfs3NnoXn1FDHOcgiqNdgSR5K5yfxMIL7wtAFd
d+LR/A5ec96YpJ1zzG5d+0Vf0f+1E/CSYmvJuDxwo7T0sgx2xxvz9v5+zr4la0CzetJVImblnRRq
vTzWu0XouyxG4FM9O3EKHDt3qr3fcrLp6b7apzAt5sFtHzpcU2u/5Rw0BPQQdZeoT+tjmI+HBU4K
IPrE4rqPZigZ9qBGh2b6CDWqo1DGE7QzMgA0CsVEoUQ6VkFauNypRZF/Ti71j60rbHWY8lJE+XCe
9MoRpvt6BuVVksR1kywA1Drm/52sstRRt+IKMs3Uu3bPIjmhReDvTwrjXYdL1lZ0hvTbyTYCKry3
vfGmVy2sY/jSSYdxXYF9S3yIz49apyRlgU2l8somdPV0Xgp0XPwysFxZ3vJ0QoiDYzN912qQyra3
TYNjKZ52Ve9az3LatF9ZCKNa57kJWF6N3wxQeAl1PJ8bquH62QAwv36tD0FyUyw491LpbhJBjcWA
YssCo6ay82o707bqdRBnBqEEiQ7219HxqUIhtBc8WSy3xO6DJ02U1uWHS6Dta+q6AoPzJOvPSST8
cXd8CJj4nbiwSncCMdi4TXgrrde3jsr60PGEDdF0Y+pHswiVF0YIFtqGwvnjbMusEJqjPZPuVJB7
ewARvok4yM8GWPQ+3RawyBLEpkmuGBFaBCgz8kT1vJRw+SRSKqEY//Z47FeVUMZma1kCwUVJhW9a
AI+bZq0Mn5ubh4mmCUjPN1w97A2KqkYcCz7zSYKKnwO3tTJICVuD/olL0b3O7DepeyYNiw6vLk1S
vFxjBaZMDqR2iHCUj5uKFklJawM6dsMwQLvUQQddJ00rfpEJKbzseqbCnijm2IpfBZ0SqOtL7Nls
l4ZSOimM+JjnDWFQ8A/V+9PvkWenF7kOV+H5qy5LGrhOTOUaE3A/XY1AN/Pht1rzCr5R/BQmuDiC
2Rw6E4kQYMU/N9R0pYVr8wxF8v0PucU/r6pssa9lCPdLxLZfregPvUW3hTxsjJU1y8I2ui4kYhU2
U6pAWtDYmI/fTEmyMWLn6/YWlSp/3jdQrcla8tZiMTHzhd1QWTOJdUbDcpeboWUhuP/4kjR7fFKZ
cTHrTSaft2AnZtjfm3fh4aQvB80MQr7g9ut/UDecszlPL06kg0rLpdGNzZbKnd0zIFZ4l561Qlza
IhKVWCYXz7bnEw4sQ+QqqDmuWCwL6fR0TCP/ak/Ik1WjSpsA4bcNCBpegqUg4L13HYeQ1HI8EU9O
hllRjjWv8AJhS2WUwIEYT3bAyePoAxUEXfZmxw+Gntg7AKBvoEi5LLur5SbkNthSdg+VFUF+rceZ
RW2E+Z5FUcJo+bzyI0DAi9o+nI9ykdBtJQ6Lz7jvyBYFCDC9T4tpFTOsTXGDPAuHF3kxlA0+N6aq
PQKnRAlvyvhosnASBbAYuDEj5ss/0qvzjqtaPamPGqog9rE819IuddtpVIoz0jFI+tnNz7w7ggN6
MLmCJtqaUpti4npOcPz6ZKTmYzbXBEVjl57hA9FWCKtUFmZ5CHRZiQ1FUx28RcPbP3AzslK3nk/c
+/H381yI3Ok9t6de/2dlcEst0sYuCCg9dszlQCKZxKztChG/rH8Z2HlZP5z7eK40Igl1OGNhMfDC
0vuKjumD+1yujHJ5oCeX1J4WzqyFcK5B4ng+uebnXuP0L+4TkcLm80/6E9IroidJisFGBjZV/Gxk
7FuD5Omr8PWhp6v/vPmUZM/TPQF0FhlLUQgXZ2vZPcQ3D+4feTIsW+VX1tpgoDXyL8KMUKjyRXRb
t29tNIpwwy6XKVi1umiNmdJQDR2kL1lxj4skuvH8mQ5m2kYB88fBwHEeIr+CHz7/MQXCdffzf3rl
NUU9h/B4oj60x+r0LHhFRjIJFgy6F0sh77QSEt9cXQYR7AbukNuziucGXccu9a17gQYtUryxQya+
BGBcamx3QDLRMGgvBbQmrb7CbeTLwea7jixoxIQZLUmntxI8rjyggYsi1Olskz1D3ucYT+IwYNDt
fBQ5OWYe1wjnN0Y1WYrGDhDiWJycH6c49iUZ7lSVApSpW0kn6upM2YbdTMBStRcknoOnpEet05Jv
jKQ0iJlMrCfO7uGz0Uoxatsnnf1//93HdFLGRgSjzK6weMAbgx2GXJQa5MUFl5u1+dA5loQxT3Dg
dNKl+ocgPbNR4to3lwIyYQi3WSg1yZ6L+82l4Et3fiWI23ucXaIsZuw9GmxabNzcVqVF4XqyFFO1
zNf8u3e/5uKZ/KV4HoxY+jh2rMbeiVRgFOG2MSWE/fIH6t3UUnpocuBZ3W99f3yrknxXm7CrLK4x
D19JuXsHNmMWQRm7IpnPPSRyChD4yp2+i2m9RqqGLIVnJPrCS4AXZOTIzYA5W8ihQbI32A54cUl5
6cABowXeJRGr5hV3+xMWdmcoNHFb6MKkwacGU8TzBx97cU3/P8iyITyllm0omgUDBhXdTWZkTv3E
FzWBPMO8BpRL7DbPXpHpyvnjUjrnWMKVYmYKNsUskQr4i2CkR+V/chBqwdRZ32oxDgqL62E9Fvu6
GgEYp5wVYerv/bZNe1VRjAoJ4vniwOtenbAft5YvNfsGrxcPjLQoOdOXvJsym3PWT0WtamdpIBkY
fz9xlP3S7uH5X4RDEiT6fLVw5fU+EEf4LnE+ni1h/SHP2XxFmcA6bSti+06hqRfNTjc7uiL0Ws2Z
moSVOvUxmHz738d6iomLwFb4MHT6n0V1+eeGi9wxEZas59eHIsswDom/V21QAs1Y4DUjqeifhz5j
ipcJ3/pHS6JjoAZu15s8k7LeVdJNbTxUqmh2fB1GcX0gG7zI3fGZlnXMH6r2djWGI29hLVXYAK2h
F2DjUHaJTMgl01qaabe5XSO28eX1NQeaSVpyitLgBHvDofxlRLLaGU7/rmskGMcGq53TJ4pGp6VD
a1EdF0i9jsydy3oO1KqITP18fsWfL6Nhl8ypwmuPwZuhPHad00nLFxNyamu7KCFAL4c7ePVr+PRY
QLjB02HXVFQpuGG/gHWidxwUJSfGPPtPdX7msoIRSc9dZJoKOSRdsPqUwoZtRQL9dAw374AkJwOP
7o12arQdzJvMSMRXVwS/jx25/aMZ9+/O0WV77spY2+MhcUhUsN/vokcpQ2Ld48XZ1y7WbJZZqHZ/
Ew0dTeZVHYKa6EGX5uGNMm+TeaGguNmsw8ryjphtBWOv4tu+sj08/GabLXouF1UbUhQcMAILEmVe
RjgFT46liKMZP72dG0NdxXdMivBZQ/bi7kQiiaMj5kVJHtFmSW87ElKCGDx06MI61YvDHD0wCtx9
PTtStmChnbHvHvvz/GTH4FVfEfCkbjvpi/zcj2nC4BQrNA0juMItL61i8k8u5b5YhI3Fw8QINSuR
oRcxRsQZ4tM4Mc6aTisJyEsfq66Fsg3IoaPe8m1T7YWB9EVvkWRuGnlJeruse5K436Wm3VuP8PsY
aE/ftPbj2ssOfw9Fbg38KlGhqwG3qhHo4dfCHzi9i+bRxPaJRJcAUAkTMhMSmEVkf7XBh+HY29jt
IoG/RuYW9v+ax4tyGyQCIh8sdjPx3TGTbHgdLAdf6rw8+xJqwVEUkB3mlEE2QgOM1ncgICmsoQ2t
NZ8srJ20U72X+Eoeo7OyT5ODXnTzWZMP2yhuB0Yb1ljt+QPDJeJ2G1D7zNoYOowQNlnrOvEq5oCg
Eu80p1G5hb+PD0MhzJtFRcFt0Ca/UAyeXDotcNBwuFGmduAunh4cT8u2lDB+E6DAt7ECoLyEgv6V
woAjYVTGF7kbb7nWu3li50VlUmNmYVxLJGo84BtY7yvn5rUjiCCYj7bWivMZetrBOr4N37bAExgI
5rpWnZGzvGjLzYglcppe/PKuV2VKvXOtvnfMx3OmL0GEErA6OEaF8nKsVlkZ8AS2Elh/nuGaDMsq
+S8UaPH/LKkSe4jW75+ZDhnxmr+K4a3NFMM5oKt8AC8VzZB96VmZsLwn8Li0x3rkQfzB2PSA0rGq
/5MPChfK1vyFRZbmfs0vjHW8Iu2bo27l0igaU6UGEMioGPBm5sfWuYovvUbs3Gb8qpmplbAOmjzy
jfaMXQZ1/ZfRZWOLv6sv3aCGwEtKInkMMBePfbz8aji7rR6FjKUwjmNEpijd4o+eQqDyl+vQvIzn
FugLoUhdpqPj/zWhuqWv/KAWVEWv1gK2qxNzCxnM08C2rq8GbLAI2DDJ8ghDTd/Yo5cLjzCTHgTL
f2FyGGIHwEmcMV8GczMeTeA12rtxThKvm3BT68H2zTJYa7gRNNwsiPS9bCfLp/SYHZ9s8mBhLPOj
RqJ30bZ/nXMT6xn3i6T6lVVDPb/bqsbtRSmhnyZECeX9QkdhVR32WvxFX6OQfHaUd00nv7L5JpmD
VuYwBaWpp6fZ7nXlKxozbVtmQSqiEMX1jLObCMgeEGYEluGlb4ZtLGaPD/tYBU0XTc5N8iaGSYWx
z0/MfJ+suvTgxcWPyillgMbzCSEfFs16b+Y2z6tpupiEp1Op0u1YiqxCPP1MavZ3LgDa4w7TxTS+
e5CcdalGoz50CheKOf4CI/SJDkDDPEqJi1/2ul4j7m5wVvTx6t8RYtuEuODLY6dI5MBCemBM54KQ
8dk9Z1lQwVuN4qkoQobVIDlndpYRITfk4DJpEjxBYfnQc+MkJ0o3Htci5rPvlM0JIslVWukMCOVD
u9PvGIPUurHU0f9L/V7TBpdNGEZOxTyx0XfsTwUoOHQY4sjrbI0xZlb7zhOe3rojR7qnFMQIloPL
ZrS8jJubwoCDJVhhAoxW4mx/AsSjd+Ejg9qL/HxVjml30RkHi31VY9A0GYD1fMU5YAPvVvxHpqY2
Gr6//CbMiJ00qp0gKxQL5sbR3SDE8ap/cmtifwBBsDE+0k3WzpfW/NSiepkPweG+XlfIzlG41zcq
5UEmpIKo3m1QwfBs+Re+Ve7G0qMdisPwwSBINTdYvzs64jiwjQ4oyM/u/hOeFZ0u1H6KepBI5W41
B/rCbsswLahuZqELwj35EkdTDVINAdso8r0aqXgmdhMR2s6Ab9o92tDCZry/58MP6wbyMLLOJn9s
f+u9cvTISNLKzI3mBQl0dbuOm0v2yHj/QOeblQ6bf3AA8Gpnj0FNJup2lKW3RLVSADQqGpdSvyMp
uqRr/YAILkP040qYXSWCysmk/qMuSOCbLrpliKRLCgTQr6Hb6We+nHV8pL2aWm8FScp6zJjIp7uQ
1X5/s4CuBP699ontkaLWFvfTvxkky/dLZT6cJZZPbRuQYEdZFBV/Z/UABdl5zQPDS5Kozy+Jl3il
Xflt+8FhOinGlyNqJ4pmkGTmItf238AMw0R5EvMbG7d016E5mBuDX2crWy8rvLX0NdDC/a+rHVyL
WtNZKMwD2ZOyk2HyIC0UL6MpAolQj3NryWsKYcsUQIDEgk5KAiSYIDxWiiTwCqngUCUpfu8PmdKY
HV6yWjm97+uRkM71gE3yqG2KfMxfZlLd3qVVfu8fwSyJ5J9fsP2xdyaysuUfCz0rwGDn9mOvP/4D
n9OkyNACF+KgF8AmKopZQJb0MX9IgJcxU1aqsms8VSmi7w3OlE+ktk6YfsVX7Z/MwMSxOKYLt5So
8neMu2i7XBgbXZ82v3dtTDR19yDkFmq1f8Fs72K3g+JhXDx2My1iCH9UEil83GYVfOW8lNizkP24
2580WeW08R+6VS1RW1aajPn76nWee4afYTda4rTGHfd2h1xUXr5PxgD6SbMmN8OkaxpnVPEpNR9x
Yf6NW/q3zc7HyHn5Aex+e/Q9TZqaFcF4PFWQXVhqFLkW6LOxcWys3cx1WuPByyl9zMVpofFZ1eII
YYHNI4zP/Tv5o7SYaORefJzPafpuxcXOo2j3R2f1Hi+2CL6xfiMPCu4FtKR4msf5m6KnJNNF3R4A
dsOixDTVuY3xugr4JspT6PxP4y/GsEKdaxSE8GTg7aEo7R5Exe+0KR9aOYrN9q7qb8uoj3K+7S0h
tkB3j4cgEqi9lwtIj65G9zlPMgNe8zzBq0/yxxXPGXOCEpD1FZS647jBGASyuc9bhJUtt82Mh/4b
4AXeJuQtp4CqwgSQJ2Gp8CE3OYq0VGJ8XkpeboabyyjsX7f3XKTRdeR8kLa+O6lbqa5gvEDg6UGU
1jAmAWZRg8d63/ak0gnIYTtkHb28Fb2IfHpaOx3aT2wNZNMb4ItrJJwlCTz7NqYTI/7HRA3n+m/P
aWfRi7XreU6IRWibTSfITfDob21ePIi0mkzowsiU39gW9WeAP0cKNQiHk8l9clMDRndKMU8oYHK2
1cv5zwD2FSl1Hufeg9lIAr/ucgoVRd4ly0xvS4GwGhN0AU/sT4DmLc+gG9RmuepL269iC7wGOphe
sMgm2nJXRrIBkGUSbZHtbLnQ1LSQkGjKIylCl7W7dULo7EXHJmTNLIrE2SEsqqCMkhmZIygZt80C
e/QJnJGEo+yaBbm/rUt0Zg5nYwsgDXORQgPk/J1vf77aiG/oXpWU38xdRbreCMA/7cfWvB1W9kaw
t7pQmwqvP1OU+tUPUboUl8S2Vv7xHTw9/4zBkB6AZB9zrvLC5v76vQHEdnOJnh8IKWIKrtd2T/fT
259jrhwJsDKb3qOVjT3SwHmUC7051SG3gykqYOLfEE+OdiESibgTl+zqEpNhjISTAbLvwDqG6bKN
Y+ierBh8Jy7zzbCsHGHId4c8UR0/H9LsxwDvuPYStl9VqepBUl1QSqXUuHYCL9kRjAFiUg3cAr4U
eSo+hXexA2hwZdLRHaltjNtok4PoRnY3NXety/He887O08jpdXPu8c4ZdoPxi8qtCkdnzSC/r6XQ
8Yt6OmkM+xDdhOC/GVWOkdEw//WOfapar9dGJUzlftjGueDgvo5CnH9jfhMbaFcygya0ygtNSG7A
UR+Ul1zPUSwpYzXS/DbDg2rbJO1XjLyvKApHWvxc0aRlh5MLtyjTzLsxIvOplQD3cLyZm962Trfj
Z5amOQAXQpM5obl6WwoPwoya4af3DLqRrVXQjxglXQ3iCuq8f/Xav6GvvpcQvSBeHEjGl2fSUyZG
ydFCCtBl1yDkIC/kv3xplJXAzHef3kn8C1wL+SdFSIFVQKONt81EJWxDEV0r05aDWIZ9g5M4bfRf
Nlitwt+Q05I51RBurBBsFjqxgtzvJF/wrwsqrLYkgg79u7ihmLZuKtF8YKwCtbH44sX1aPRx7M2W
9fFKekJwbVoGtnvMPOWe1ftba/5LX5VdmInT3zJYxopaF+i4fr52EEOn+0LzNKELyGdI5o475kWI
54Ag5bmRMhA1AAzhY5ARZOmqtMGokDWaYx/HE7l5qbTTRXuNa2NCS/o4Um6tcnLNDpHPYmXE/FeK
rm5tFLz+lX3TcAKeFoeCLL6Zqz+1o3TWvCfTAADqiBRzix3yFHQTc3kG7bUk+q7+z2KFopgdX/dh
eqv+wIOIxaIwudRle8FaDoCi4rjk0VL6uSXengKqAQxYXlITFfkpxm+sdOlJ65kAtTyS7YtDvnr+
U3HHmzXPSwRUKQqjTZ0SK/EO24JcZvDK+JjG5VSOig/WCBT89fmClZyF2ncjJ1a4vKLxQaMUUSVi
wuTip917ECvFQOMtAn6gC0cHH2mduqtqXSBg9KejyC8G+63XdaSiCmXwfwVxmB3W2gmKieQKhbTv
glnrFoV0fBPMZvJ0+TQpCrVtYfE3/L92etJ2WzsjZSEoh6QO/qH0ao7XAbK83UJOSlepqdzBe4xv
V1BBE6zOv/eIHewiN5+oelH5GKQyt7DQId1uaQRw42FcNCOcrkr4v+dY3eb1JACIWF2PxmEEAALa
o5v03Ow9uaY9GPSKC+MRiQ3987JrbQ7FrF3fkKPWSOm/v3WRX2ISyf1T8YH4GsSQJ2sxgFQ8e25e
mRoAzkWGPT9SBcVax2yFk+UkVcOGVdMH/SJfRYvZPMjee7Fx7D5yTEgsi6say0RJEABWqwOFf8BM
vTU8jwCU5IugnhrTVluAk9F1wQuZjYv+gb5tQlqbcSsyKhyPw/dDmEPL229O9j0uhXSH0mDf3ZMI
GXqzfMtoF/xgA0KVYknD4ve2sMuJckV4Ci8zqec+CRlbxpCl1qLYP46XkWW7+G8IH33yZy+/pOBB
+v6Obf+ND2q+NFltoh6lQYjOK6rNOzdw6aQ61jis16U08nC29MpgXdxQrsnYMvuM73yKWCHfXTcV
c2rplpOzvTZTpx5fgt65J3urDUhhAuWfGAu2RskT2yTYEHdYa8QRhlju/cOY7K19uOjEZGTwyAwo
tBE2XODg41nfk/o5NzLBX8MDEIyFmqwF10Fb3zavTyaTYZ3y5ZbDULvia+JsrPdVMPcnTf4p85tQ
YHl+zY9IL/Eux8tTmKkw/5FgiJ2Dlrdtk4n/TnpswhZFtFE86kShVVfxUM1jXGu9w7zAbDSeXx03
oBwCZj3owupH1RPxM/vyZUI35cR1RgJ/rRk+DBfxgrLoWgFyhn+hqAY/ticWx+byT88VRflDSomI
sMR+4C0AvoIZ5Uhs1IJhNlsE/kXSI9poyPCMByTIyshzmCIfkO+1cTX0AsjQr3n/P12qoTCYEAqi
dfn838Ub1iCPhoWzotP2T0f2tyHaILvnkrW+t8vk6DcNLYbD+fE1RBuPiuotkFfORacvFwIjGOTK
CRXnI4JkP+cFT5/SbWQWBTf+FIhRsQJiAGS49dFleBFskeywbl2Mq6tAPeHXkjTYbgwaAtRDVtyl
fbB2iOmeP9pb26iVfaCSmsBlfBFF5u8EAe8eitstv2kgLmzyRYPeCOzMhSybHPeMhNdcDR7L0DN+
8QG9xDaFskAWJvk98Sf9y6KvSOhuVOTKeUSJXPvXR5bcnHU25vPnPBv7c+k5fVbpe7dd4VXrHhtp
NW6M7VzNgGItwtcgoZDSpxps+oZy5ZmZLUzoGTIGuqeTwiXo/7iOopYEXBfMtDR38/CRT69t+3JI
qgdnWTwNBo+rlHGF4Aa5iksDqt5ZcuzB3qh9oHC+tC2Dje61q6NwG2AQwJtaLUrqkNZfqKKpu6ug
5POl0ZrmF56LrsUETQK/t4dEi7sx1LuYzvbiHqNQ9r5BJjtSUXzZ+BNwxQI7GLWyyQNOkHToQ5oz
l9VbnZnom5C9uCxtaTTe2lKbqrarggzRUSkjVLxQt916ooYCF8XKrQV4/TgG5mMQiPOkPtE8y+u/
ihV9oTosAWh3inIhxSVypONMMVjeQaefde9KABkeAnEQ/moTvx2s8mXzQ33YMw2Q1SBzvAIWr33K
Miw0qDztIEhjUKGUyEvSGiGJXvb+ndASUNyyS5IkR8t05aj8OHf1R68L8OYyQv7ZSCEcABRdEWRr
gWvh21/S3kPFZ2CMRiue4fHptnZxZeRRkCUbL/5fXuknDyyq6FLSUWCuS1QVOr80Zrp+L632N7jM
aSse7RaG1SQh8iI3wOm+mgCpsTbtNx01eyECc6krMsUZTBv6KlVn1Vz959rUrBtDrV8r4c8JYCUJ
KrvzP+2s78CmBV0cuDSrAOVDcoWbCnVOwG7rvL91nmSRtI1wyxjKcYU3UHveaO+Dq2W+7m5ggcom
VG5S5E2sDWaDO30vk5/w9gAV/s3WvOAxFpUVZO6qsu2CTOt2a6wr33Rjh/Uhm7V0wRZJ6hMknmC4
w1WTIQPyhI123Ick0JbwbcR+AVvivfDpwLIR4npW91JJUQzNsCalAFffIetRQ1rLuvT3wT10SOFY
XZ4xuyVV45KtBLrhWTtbxdYkl742oFKlOShFLekzELVUqaJtQ+uXDnj3/xnslDNsaemUPJsJxPSE
O5Df11dVIHJnQ6tSehDjt3o65yhdZorWhOJAgWRAxeSIpU51B9sXDqt6fa+zsyDrh0QQftOnbGYx
i/T434WkMZFmOknJO1vWEJ+LrXGUz2q/XX2dOlbiQG4r8B+To04Ko2tMI1E+6lTiMT90gRb9aRBv
cMrOiKL7rGdnF6AIPdMR6mfNuGE90hS/OMBpddozGN8VxWUXonNwLtPiRyz4r7LIVu7hVbQh6hbC
n9Hib6ff959X6/eS+aXTvu5NZTroQIuAn2w7SWCSsrbrW2ZoOqkJUthvUuwpMGGdsTML4Rz5//T+
qFsIfXDWd3nKqAinaVwYOnGQsfSgwz8tRvJDIfIrfDQelkMBgxTVbir78NugSAY3pG3tags3lAhF
4OzTdJ0Ooiplgv+DkrAdCWlLdfFkhTwTeKU72OgKGlWXYsRn+kGiznuZnOMK0XIEso3bjVk9iFfy
bivWYQ3KTeqFTEf4MFoqQ4S3bkYiPOHFmWwTBg7THgY6RY+N4WtX8kjeShf62aPn5uNoBBQ8HOBy
Fz1AwR1/z0JG0uggiMwaZ0WxyuYAFt7O3MnIkICa19dqGmqaQFS+nvH56hofsuFjPgihGNHfQtCI
U7kwvHH79rM+ztjS6Da8+qfmJr8h/9SaPPkqITv9hu/OM+UNh2PXNdONuvWTFUJEAxp8FdqCOsZH
ft/aO2ojEdGgb8bvrb/M8rN6lQahwcnP2Ik9i+ybOZwl8PoVH1mBD/rNWDVaEbL8Av/6BY3RgXgs
2xRTlJ12dhhdTL82Q4rv4nguYgQ7QqNAKFp2HFwkd+IySD6SASivdphTysP/577hmw1yuUIWRGsZ
G/PDXNZK1i21ydwz2D6E+aJajMpsRkbA2Z5raQWqDidyoZbyCilLARnNITWh9sFtulAEznQpaSsk
KyxXBZ2wW3FwyPSPgQFk0gFcteCym9pTyHNxAstPwPbTz1ZIRS4KR0x5puDqR2NnQZ/sf6xAh+5K
6+JLYxnrbBjJXwXHYDbwdhS7toDquc3N58fnPgik0lcV6vgtaYLw8/DfslPgrcZoQS6nuAISnVrU
j1ZTh4hB/nfy0vsD9TjSQHKvlX5b4ENSYdiaOJpXLLHePYokgfWXNNG6YeWFAkH5E3mAT2nTZeCU
HqUIq24L1TmgM/FPK1Svy28QK93RcpYwkeD7R4nEyaEwRlJPjJGhXnRWPGxfKQRPyIrkF83Lmi3d
K/2JklPVyL86nihZV6nB/J14x28LYe8nPkpas7e459HIOsLWXhbuBvKAogCku7V/54A3mwEd7Ny7
6h8YrdbBxLtYwXImv0Hydia+ocdEtPw0BS97rg9nQ0ii9dCM0yCw/8LAZeJa6r553+C4XUevJGUI
wKukdkCn/HXfXVzZQvIaNKYlx5LW0DOE/U2Abt/Yhr0N9aoZ0TZ96IOPV6+bMArB9BB0nsYv6Qne
ewm1qfbo2tWqH5gGsDaHBOyhnGsI7Es+1e725DyddUy3PVe1RhE8pHSFIvij+/2Rj5wDt0odnbk1
kIROhAvK/XcMBL/0zMxbW/3Y4nl/LZznz81LwATx6zhihSSzPDzkaRdRILyR/RutUA8vqsnArYmd
Q4nfk343fEg7nqE6pYMNNw+6bPU1cjw/It0YdfMBLY8nRUJ2RdYJ8j7HoUxWwJmcys6J9ylDdUVG
wQ4LFpI90VAGeljusqw4N/rPC3l5DnwtOj63g2V76Bz738dKjH28I7GuL1fDjW1tRFf9dKkHZB7c
SrEnyqYCr1LXBixfQkIx1FCUejtT6PQg3G2D5vEucm9NTyLg8Oy1w0ASwcHiqGi/rW/9UC5qRSNp
AAL2xLnbEKAy2dyrtwIlwRq6s6DCm86w9wh4D0EaEae46jMQwBzztu2ILPfZj4da4FwkhqyFZ4aZ
Q/BwITjO1LBhsxmge0CWde8rfFcNd/vrd3marzulc0+Iixzcl/SXOas5pDlEDGz0327pyIDacdnb
7oKw/f/ZmCXLhjekyvRXLg883daX3xOearjCM4s80KcEs6j47Mm2UPiNXxvpUgSoJj3xPu+CW7tz
Yp0oyhT9gLAAQjlgLIBUQxheVHVEBfvSNH8St5DDU3dntqvvPOemXK//5nrZDstmgZqCX3Q/jxpq
wePzpaLahXfBlQJKP1U4jYCrCsjzJBP2IibqW3yEKTECpF6H1haRCSAwyGm6pDTDFTs5DJZloSI4
DEZrUw0R/Drj7tVAqZk86t2ENKIYdQqq+okIlyBr28HIdCPF90fosGLnFSClW6nj+8vtaKih5vo1
QkX1u0g0B+Uxfs1WyT99TKogbqDongIGbDw9HPL63K2eV+d5HRR4o8esf5wHU7fMPcSXU4pY6A3Z
DGoGcMopu3dCTQE9KKxSUNFxmWOeC4knAcL8efafMLJCwshxUHjPvQF5WTxpIRfIKxWV8LzEl/MZ
gMmZNFMem3Un/Sv0DUOHv9utxNPxZQXN0WKTH37Y8JXTxIYtSw6keS7dUl6mmVWU4LkHZLWca9Py
BIj4td2FIWL7e7WqpvIbuhQGyfatJWAMQdUvmQmCiM46oQxqa3R2oIV12s3tcYtjo2Frppj7Tbtm
JZAxGr9UjQG9BAdxJLG6bZoSRMg8gXYqw6UYhek75U1Y2C6JnwH0+5p9sqiYtvOBE4hOCtATc0lI
T3I0+qqss7yEpcrojbu+Z9v5klhnkPH+cUW2u5wbGpVj+sZZ77ReKtTLz6Sycg3H/mWtipJBpfME
Hj9cEpviA4wGDh+ryEHK5hfxLSu+TJg7yXZJeHupvM5Tnl+wLPxTG1kvX1YcJvfvvtJsDiWKkEhx
vLY19mFj3TL/oVg7oUfdsI4ygzgpQlMEAOMq2HDG2g/Sdgja8guaB7j8r57R7yPg/zT48fdpUGyI
i6IYcdFliVSqojwi9sbHzVW23S+z1JOzyNyCtezU24b/q6FHzsgcGeGAtlSgIEXhnfRCRNj7kaHZ
G9c0r87glayCqUkB8VbZPvcY7Jg9z9dcCvFWeHM3J6PSv2YH+coeboJWle2z7QGYcTmdK+FDtOC2
vAM2L2jOWR7Bteq0I/WLGTq8pIYkXNX0Aqjg2Vd6OCc4DuXtUZwqdMUY9A2NjTSYd9WQhhY8EHvk
1TUWiLXX+uxg/kv3yoo4uQLe6cA9f3PTH5AUzUTOhvTywC9N7C64zgbnha0klRSgEm4kHW89KJzF
H69wGfXSyP3WYysdeucCG68DalU+YW2fSgEmiMZe4h78FG/sLTzoDCpw09sOKzNyHpgVdFDrTjCK
na93HoEksBfDvSRP4MrSN+vQsTwtZTNI/gTSP2t9axgKeEu9XK8mkiuVCqNdCdXfOuAipLwq79UE
pfE4UCFjbGhQK1D6AT2U/QFaLfAQFUa0cYBnRYirqrLYNS8LB3aa4hbYy/LNFMCoYvl/UdkXNmlR
K0zrQrFIcKRgjdbZly8XfxxQ5OpRxijPElKRknmW0xa9BKuyB3t6vzK1Tt9Cya7qUC1czq5O27tJ
sMLl/c6BNg7xdzF2daTCu0QDju7/oRYFphQxdL8Pd/HT4HwPs4tCHfTHAkGzebSFrPVjxVY62oMn
qRhmWo62bKAqi6vlM4HpHqHTDAFlxmFU6ygM7nH4d1EWXsmSbJBEO4R0J1JcYXYwL+/ZMUXVnHbI
IhDTQx+I85LqG8k0Nb1t39X96QDYfciWZ6bAYJuRpYo56nhY91C5ZP0BF9dig1A1fLNhQB7J6G/G
7CNdoZ5xr9WXafKXWACIzWxcERZm74ICglKCAZa3CgtJXvyJgu+QKk1G3L8Il38pKyH8yQnDDUkq
kF8hs/voEvPgpmQuejV29FQVvPQI44wO4+lBbT+wTmi58U6PXf1uX7LN5pPU81cJhmBNoR82AByy
z/fF2vFSUKKf5GiQrJfbF/g6zfo5HI03YxMpHSEyv9tkI3srMCmP3CNul2NykqCZYngwnRtff/Ss
UFh1GjO2AEHBXPFqW1bxZ6VirzA9qJXNiD73VV/6c4vO6/K+L1ltMyjX7hpPhe/8JIvgj7lSq6X3
0iT+ERjItZCHPYXkVu3ajhIdET/W1Vbvzy/Y1W3yllsNU77dqPsEHqGY74DVOs7kqtpkEkJkeweU
z9z68S6U97T2isWVNXI98FwwZobyME7yfTjDV+CcaoUOzzPx2nshrlA1twpK1hEG7WvT66/Eazmt
akY7BkoMKLCgMX0RwOOWClV8eDtQYg8koo4YEECGAKJqsKznwOHlQGeULmkwyPPy2mEDvotKxef9
D8wKY5CvFXtxpjO45kCS+OJX4vw62G5fzFnlvDO5fb5Qh924m9PJM6Rr5gNpdxFzHnuiPdGqOK0Q
NvTzsn/WvI/qHf61+rkvnXVuGQEn8t7AszOS2cln/bav3eHJKqmptb1FNGWbM63XJ+I+6x8dO55h
JITVvIBvFzGWOpmluGDOEwFbuXvS8KzASM8vjF31JX/fxE5b1ryV1oUfsgtNn6uHey0VqVXU4B3T
knAS/Pbi0ereOASWG+ASg2IiK8yP0VHCEGk2iiSsRRAF0yZnmaPNlgRKIoSjIa+yoWRdpqY5Tj8W
b/o66FaXTvSBm96hfOVzk5rtIqbhgMxtJkQSem3IE1qjI8+N0OjgVHvPoIQbs4xkG8/KnSvDmSdC
Q3P1xS295lUctM8ggb+FtfDOonYvbKC0JbihayHE+81G621H3QcfHi90axyEYYMgcSpYzqpmFSxw
8JAHhAlZVaypYEOLYUubju6k3sGQAAVPLgK//Lg8u96KqY9EFZnQj3BLdtGapqguMTvWbf3/gfIQ
UoGOv6pVfxvMnPR7EDWtIzpYdAXJArCgjR6qkMyE31DYY3ZwsaiKorLHVH+OrnQDOySFmH3fzlrv
4iERPN+5XOOxy3kIgV5OMZkA4sADGbenDStfxpey/Gb7TKvzKyO8lLoY2QZ+8M7aA9Ywhuukaw1o
jaDEp43NSwqo37N38zliEjD+yzApMMJbpt2tZ2+6fbVD/25DLJmJqu1JvypMN/EdKR1wzaefC2tY
2Jn2AKtnruCnpjcKqILCixxx4EV572l9YX6/xq6p7KsdIlpQRxqrVV8C9rNSbWr4pSNPL6PyhY/I
PkTOEJ+F7wXM3i1NRwmeRv/AiaFgRaZCgIg3MB4x6E6OaQjckkgtemuiGzs+jadHZETdUoaAkVBg
RylXpj9M3Vi0pEKiSJ4XXpo4nL8JZbS6nB7yTGOOTKBVowT56tjsOqKNPvUY5vlQRtrvXLuihhfK
wuaKe/nWfUUHdqXl8UY02WL7rDpJTsh25yl7gm0rDrdpShsjfHgjozlaiLg+gsNjUVJ7J6iyAUa6
m6OpC1LNImdMwCKRkak6KuC+MncEbm1DjhvX7z7+GAZ6XyCUuqLLGE3ddUJr4mjyFkI0Hn0i+pVs
fNcPmWpqrypLvuN7IyHXSHjm2/o8DPZbG5fXm61Lxp7wXnIKXIk8s5xrJyAJcKbgPDQ9FZ8Xsaw+
IDMcI7BMumCvIzGQZF/Z7RhDgofe/yNkE6kVnNAct4dfDgnJ3I3nBie1SIagwV7H6nVSj/yN1Vg1
P3K8J6eq5VCfXonyXIOqVyUAufCddh8Xn+iFw6/hu/IyOP1KxN6xjfBR0JqsVnRaTPC9zn8UKaz0
xb++ENNjN0Cev+UR7Ui8KfFyIkj8w/Z9KW7QsCkGXOrUCJQ5dloUg5LCGGfTRtg65FfjcJK/jHVJ
46/cBibeRAUyN/Jww9qMyhSCoh7UgII0nqVdBC2VkD6OCZnrg41JJ3VDa3CTRCZEMNffgMzncwxj
O8MgSybYhpLWD48h5otoU/TmRQCkDybqSvIlVpvsJSvm78ilzB3dvVL/KAhA9asd9db52hbMEGNk
sDDsd6vLSZKqNUkrc3GuuakfhhCkbI0V+hnl8vXKZwTV8B8tDV5+cg23KK3LZm3RhO1mGNEuUtZV
969P5gTZBUO8Q6oprDph0zEnH1blLAHwKKALUf2uEaVjSZMEP+kON7Gh6REBH4y7R68xEQ5e7UUK
QVu0VWrJsT1odrqGiAxbiedrASNKwcSl0oMLYgh5OJ968fBHfIs8vnpdIm5W8JV8nm4IFoCtabRu
v78qh7+4a+0qQ8wexroGgzKqSJgSKSWIoroziPXvVXP90fmNWKqdAqOeFLcHByFnxh51+EgoFLPk
95FS5/MkrGTnu6G5lppRGBlImeR0XSukdLYFG/hlClBA4Zdi139kdSvdqC6vCY/0Ql/24tr88Qry
RE7P27xngH/Z2cNr6DVKpehgWHXPn9kGX85F3W7jrj7e0AaH6V8qP/9psVqfXOHiq9n7aTLRYzRB
4Bfwm3D/WJZfTmYFkRYwLWyT3/iVGc/zeivp3W2KEnDoDRN/hKO9FrtNkMd0ICBkqiAQloXKMQtv
cGQ3jy692mbOe6MpYb3ZgQ4CR1tk0U3avLdw/aNie1fCLE/Alu/Bamc+QTwfSymaDV6m67Xns0J6
zeZAUmY4+ksLiwEdR+HcKdK0lNkjZARLfafwraKlhsgxTSHbuODqBTdcYeRQLbG3qC6pFh1qwn4V
88wgIPVdjIzvMpjeX8q83a7yJFrn8yNd59QgPWBf4HFIsPGQ3p5OsnsGEYZoK5SBA/4LrEGdkSh7
32a7XhN1oz/pMiBza07HmwcGYmchKe3bieyH2Z2hgJ7S5sRRGxTH8EP3ckRSKOWBCg+7tDEaEJYH
JLfwPyPq3JLzN7xvQhNQyUKExbXdXzIFOyS2xgdcG1TxCLbg0YvQEbmk7wu3Pm8syTxM7dyD0/YA
wYKpSyfMAiltiqh6tVUiC0gNuDtUsIIdeCBKDD41j39iLv+wLy8kKOKJPG9U4amqU3Pw+zGptKCc
NR5Zs7lNLoyAU/asJRpbdLAR5Elqxps8MTFdX4VZqPJDyY2Lg741cajQ1yhDihy1QT/c1wbfSz9o
t8KjAVkPaDb63tMlpzzcgxUZOpWk+v1vG8vtMWV5joMawaVaUZENqb51oesbU00n6wSPUQ7FHLtZ
ZCxcUvoItbp1BqDkWsAScZKnCsJjkdFMMre93tp8wuhdTbfwLu1nYofQIpdHstlXnQNURel2U7zv
pfiAHsVWyqRRbY7kSH+uc7QVBPT6nNBWO45vDhEcrU7yumADYtJpoVC+UtVr5dgkhwUkzE3OPXQC
H0PDEHVbDAQQZyr6lB1IVvPtv4kgINnFrRrSwvOHl70iqJHsBDRoyrEgq+6UyAymr6x8UnceNIRH
0SQZHLYy53KXf79V6mthW1x4/15LhGmmixmdOXkeIfUdWYpT6JzChFADd2LUR7IgGvS2qH+AncxW
0FWCjesDla1Pk0zyRSOcM34e2i0iWHanoOJpm3uHEnoNvy+aIOec+PPShBLYzMnvYAd+GipqBQjC
1hIsiIZh8t4ptLOkdAT9kmFQa0U1Xmg57yIaFWc756cJpjF15QawtEpzvTTzBsU23BWTiJKgQ9Fl
bHjncAkBtujbiT4WwMirPcA4Qh8XlMqOcZxYoSb88Xu04IzGLtUpIOC0XYgfay3kBoQhkx6RE+6Z
LJWDc53tm6j131aZkvEZdLkAArFuh/qAilYtf7yEooCFPagGA+S8JQdzA/ll+Slgvc2zv5J+PNm/
6bCo7SPeBfFNakQPNK+OuAqL+nl7T6I9HAr5bam4O3jFbEqMepPiOPrUbjD0YVGRyAhNVm3hzKbv
LlEdqAKlDv0h3nNoV2ycQtEgDRb5GPtG84AtdldQOYImNp50Qibw+pjyU7BQTttX8HJZcwJNInKu
uYS3lC25E7YxKC339WW8TqfabVjlC3jRVmhWeyk0MxZYVPVfg4bY8ibHJdIiRzn5LN5WfbPizIs6
bQPioPgnPjrLkFg0A2nsEm8eIR4q2GDN4W2Nhzpm8LFdg8n8yvep25Rv8CjYmoCrms4rHmAMLhTa
CGVa6o/aBKc0UO1wEqi0LbjTmxaoO6gVjynMPtnDWQn09pz9uRW8bKT6n39xu7rTDzwWWtvMCbfl
bgURL1++N/4rTIZ86HsxNMBgLpzrj9LCSZQ7U2jvLWljNPl1B9APn3kUdb9iDhBJNRmHdzQxdS8J
ZpEH+yd/vokLGybCqzrGNIZLLCcgYj1Bdf2IaXCkR4bqhbhIdnGsjvjpxEj5fpyQ1TxJhP3Vp4Pd
LxXATM+QxwpgbXEpk+S1xVZ2sde8PgD2FEuElV6/oPezKhD+XOE8IRm9dfs+X6c1qJ3qXIPixmlS
yhn5PnKC/kH/jSpRisynUtDaIdxBTg+QRPmmGdja0HSG9Xbd5PGhTP5rRew5DLpv3bonRmzyqIMN
HlmNqawgA7aoxXD2kDGxoTGuyT3rqlT3kK50uF7KsO51VWHpa0KES/8UrOVehmLbw8ARqcHwQhUv
d0ZEE8CNlNvXsRP2bGFUtutLnWDQ/gEyGj5/b6zyU0JuWANF9f5XUGdVNrjlHGjmY2isUK9ymlZS
3UuByTS3f7ZqbigngajWqC0ehjSM/L1sS1NXSQVMFE9NGqgy+atOUTgKZXozhnbdvCbN2EBLxyUu
/YmI2vebqsAqwipwMf+JsPCS54yuVFcrAp4Nqsf17FTnTcJSRCQnxBu0TPI2Tx3qlLCHwvYpB3Jj
DwTimKwx/xNKlkCzsSH+dyvbWxmC+QIsvQrJCbYUsUZQ4/XUhBMAGJSEj83A+MQYvlb+JD8mt1gs
vqWos6tpt9SORNU9VrKQ/uB7iKiyZlEGb7b0NC6R5ODR0DS0yPmgbSBXLCFAhUbP3tL2vRUBzn3A
HFAxpuv2mLOYiwh3UL08E5b9D+DcTmrJkqsHHA1oSHfHSO4PTWUuRZDm+i9dsXEsVqJ/w7gEbZrd
bWU3/+VpcdSD3ILPR95ocZqdrQBR0EN0OYTIR7xu7AnWYHTcKj04O1w6cvYk9EdHaRIwc+0oA2HG
XCVZ2e/PFSSxk7AjMXlaDuWHVg6s5IHFqKdNUKy8ncrSt14GSHDQn1omc2NMDslk47RbPHXjx/vM
WTwt3Rx76nzeddf+7MADba7IHjE7t/8HAqs2CtJRBpVpiVKqAl8THvVgi67mAMJAsQfgnXL7aJms
IswjhwixrsZqL98aLMo98HZBgcyvfeyVOmNcRuM3/1EkRFdtEmU6Cy0wU9eNuOWjl3bx2+tGoXEq
FWx2+4lwCiYuTSw54wD/oDdEGaf25KVpcCUhhzzWNBq7M31ZCJD6DbOHhsu1LpeFOSLC2biiX2E5
2Eky+EzvcMTx0LFHVoxzvDcJndlZbxonBMsQUZ3g89Onk9qKlVXV5VxFy724uxy7OYzNmaZPQnkD
82qNliuTgkFjHUvmRice4pXMSusZkYoUQqVrDtGqmj+azVfd9eBlY9tO6v50uxJbw3+pKo10P/gk
NR1rfBWq9BcOG0zgZzgq0vB9Skme42hx8i+IfdrCZYGPq4J6F5zEHK6pycYEyVVsATRDuVy6KYvH
c/eoScsyH6RgUdoegb+5w7xcOtEbhm9m7JVgvHbqXjHrZMXTYN/L+xYqSgvphbdN9922KnNfXKZy
QY6lcC+bQdxymWeNo3HbHKVM7KRwSsStF+swBKZ6gcTp962NAq/9cwSoSohKHndNkinHmqzbCefy
g3FM9xHs57SZtE1mtGvNEV3iP5U8TRa3k4J6DiOK7tlo49XXkvV4EUMvRAU7ckJgvcfePOWhGCF8
P1LzBBZBqd9DgQnHdVJhg64X0eMOya+x30vSOdWWgx8QAjj6kpwqjCp6/D6MIyCWanrEHtZrTUiY
7P7FFLhbTLcGsAi179cP/CzygzmTA8B6ig7kswBthNjaOA0GIZFlrpGONxNJX9/mRv/0Fj6F2UiE
o8Buu9/eZjm5z1YkzAN3arV6Sx6yg+DfQfuEslXP7vuiDlOmCAIPCLMTZRSrw6KkLaqCq8UTAVmL
/fst6mqPs1r1eLg9OoDKEavf+R7BKV4Xhk+NGsnPKyDmXSENrSKHepfwbWX4nDm7SyFdSXHZGcBb
CyWtlDSYPAc9casOxxjOlTVkEFpMUjRuBCqBuzwkG5jE8jcNnNNn3R2wSNgZXrgfosQwIF4JJWkr
xQ7dp/Ut255K8GvVfH5ctbRpwOjMTtAqmBJNAhX/f+JGwA3RVERPlCiinR/tCnYygiG/O8soVKHH
IpU14ibKSxOIjsaCNQnvHM4V5g1IIBEoUMzx1Shh4If//4cxz02sk0hnlKXvLFKpWIHsAzahw69I
ZB24s6bGsXoOsYhj8aY4x6Up3GeW2iEOuNTtrO0yMkkINYD/TxoA38dgHEpTbtXmuXBhjtJ92nWd
Pm1EXN936MKwuaIV6zlvDfypN2quWAToAPns0wnW1QaY0v1eGhPY2uYc277AtlA4aK/YTXqWGMxp
omD5lfB8HRCvowEui1WNfjliRb0MWDPZpdLTxkKbb2KMT2GxDMzRXehEQtgvljgIkA2AHqfLqmcg
1XvzLKbeUGc2xfR+9S31LfQqhWJiiXtNeYKqDq9ND31zkgOHy5joYAShV0qV8gZdu9sxr2V7BbRM
ZQzxXo+EHXvVaRn8d9CZ3ybcVq4YTQ+NfOW3bi7pvj9a5qQzKCKRKWdwqnEjcK+0hq/gBkFp9ipq
eUdRzrnKIrngrDIidXBbJy0Ucd93yNXyX70NPrM+fGgTCuPFG8Tkin/PgSjoW6Nt8DxHbwH+Eb4Z
CCSgq5cyB6//rTlIQZRs7kRia6P5F2ouyLAPjx6/ivqjcMnI2otaMx1lflXCxGhDM2/izATPE092
vFlajwmYsZtYCGU8O/mH7mSapLwF73wmHEjLz9H1R4WMRKHUBl9a5lA9G14rNAeipLLORVWbq1tn
bbbY/Kq9Ec0+EDRSWevMA6DdOft4+QZqNR7mIqDAEWBgfYsACakOKBLG64iv2yysGirz2diFqcYf
utITvU47hZId3+YzAC5jHIf1a0sCtc2wHidwoT5ieV9MqcyoIXFtWzLtl6lGWAuPjMSFc3iJP0KY
tlSVDopcr10JCcIuvAWsEQ7/S0fbuPeHHbgxYgJWckXk/r7vTHBct7GfQqCWx4EMQQvszbZ4xkc2
ZojCoRdIzE+2j0Q8IeTGDlze6Rqnx2AY7eXJenwmh3k915rwnJ8ZTiKT6z69u3OYULD7R303VVAx
5bF25htFxljoQHaiRd6IZv7VMcq5TDSVyOUplebaY+/+nSBd70lrsaJGrNsRBPhhv1IH8csen8rm
AtcLbmm9KF+kGTQoJUwDjw9ww+PTbyiWxm/RmsTRPEEHPqtXStMc0eS4R47yEhdTDAjhOzpfhnUI
hxrgDLqW1kNG4DW9YnH6RFJab38j5S+jvHoPV482hQXt0MXse1nql3P6KlIYDxkmRidas32Ktc1e
Fd6FPKjAtMTBzdEiA1yu4KGYtyWjOgORbu+JZCN3/UeyzcKcPrY5y5IbfJnpRw1KHgkYcR38SYJn
JkMlk52ZiDaulq9L8/kaoeZXyESuqnBHAawcy7HgHMMza05la4GSqxKv94/UNs43cWkg1r9G+T2b
hpmcqFGvw+sxC7WFgmmCH0ChYN87RGgeXwwPR9FIqUUiLNF8P+YZfEXUZ4zxZVq0jFwxdcHmbQ70
rbZdJ6qD1Av75t/dptnHiNc9PMq0DcDb9aPNhNefy5Gjmd6VWTV5qmmJp8lWEOAfpl785JN7tGJC
fm7ImvO+8s5zqOxYEfebVkxe27I5HxBdSfqfyE18xEw2XSoGZCvWQX5GH4/oCelLtaTpRx6kyLMG
oHqWgk+rm6YTusPnBUHGSN+5zIGAnzFeWxDV76lq6H2V6HM8nTT1TgOh6ODgBIXoCKuLNANjLHU5
sKX9/GLd4/5L7pHW4zTeqtIuqPkiUfQ++0kfNTmo41d27aaRWp769X19q+lMpmaqkHTDB5EiRqwD
LCy9smYwOjg4PGk3XXPlQzdJq+3x2mjyhd64pupJ8bsOCqxWXG9EWxdQH7Q5sh7pBtYh5jt+jviI
CnnYANyfuihwp0I9m8XdihKTv1IecLqDlFAUzb0Tm9RNdXr7oJ8bMqHNKL/qPp+UNsUOjzdyF38F
JsDjzUigWz5D7RC5l1Lej3kZddr8HD7irhSL+ltzxhVCAzaAIDu9jSe8VbJ+YdiU4JUPGwTFjPlX
HpjAr2MmmuBYepCJzc8qJMfYVKtFZUVTvEfjU+GN5AjkzCj8WDMWsZA1Qu+gGgvuXY/h8xfmM+4q
upr3d4rS+v8nMlVNgDIXabsgwq97mjLsYPjskRRjvVh2N76HqcfGCVuxRyMyhiJzzaEBDVUMa0jb
lY9h3NiZJQV0s2e6d0Ef1nyNmoWBsexTMgzLecmnj4yAMQeDmqE8dqH66XndKB8ukKG6my9pJ17H
pza0V9YBm74nQv0oIzZFRwykCu9HPJXH5n10GHQa4nm5nRBBLiBEzMLWMuz9u1yHVdoobr9R+Iw+
TEMusmaa0W14wo62t915F8ugQNFPnGjQUZRPD6NpFMfPSK6kYbU6qcSXlQjRILC3SlcuOYlyLs+W
1wYKn/4TPhJ7+/o6j/n2HJe2InxQEb/bp5TgTK7di27Bl/Ss1bY431nAsF6uLfLBm51++aBPi/gD
t1rMCnqUbzNuAFWspLPZi3qkMGbSRN/FXJfNxpeJF2JQHlwC3anW+s0W3hIfo4nAQvqxVHwrrPtX
GaC67BcEkzlD8090g1hrR+RKqF29aOV/kZP4jeLdTh44n/zWgl6TIlQWNamrraxjBwERf+2GTNaY
QzV+i/pGgX+GNZ1nxlcHzvC04cxVNeXS8OpovB2hzIFPXEunWH9FcFeFIeLeheeF4b7KOGRKobxB
0fllv081z7MuntRiwoDizi7TDWiO3EMguxxqKVX+rL1njHrmfX+jNDMF0CBf2O/KzUvYVWNduzF+
bc5cgLy7aak7Lf4wJ3bYPtz+sf5ze2CudkVKC0SFm9H8D7OmF7LDdEgDg/pcmFi6F8aQOoXr8wNc
McLRtUFmkwUCYT7NN61j3YcT9v9705JCMAgwP34PiXEpmAXuuVtyL1FXUmCWiGdSnuvpkZP0EDYc
x8tOZD8TjV69ZhVZZDPUQEdoXq6UxrZ6S+0/PuThZKW9D1xIrbWfwaRGe0B+7JEz0HP7jHgRu6xt
rT0TIK6Wssk8yKTyKfXZefzpjhf0xN0F1ByvlgF6KvbMqkODXk7529JY/dZt9qYE/TZ2SUcfYPtJ
eGGlusiyAdPPlsNgz2BBIy1ofMPD0v49yPpd3LhoA7yi+9Nmh4oO6jah3RFIq0oXR8qQfH5iKNyE
cxFhcpAbMEnJTd3Vv2FlFtTJbwBK8LzWpAP4Tl5Wt4FPQSfjkAp6p1RpMIdbfqIS0KazfFpfeghf
EfRgbxtpfdckX7To4RykLhN+xhPXz01Fe6rJwjcwfqa+AnRkSasa1ybvh1/kjPVM5c8xXndmEb53
or49Z2FTWvpyECu2xI1VBTeUl6rbjCBBTxDqASuFihzamzX92JDNokxB6ckOA+PWHy7V+y00RYa5
WGcFQU0zgDTITiEEaGhCAYnkkAlHUdej5wdblOmG+MpMGaKULOmDf4AWYcLadr6U/iOlw1JG2YzN
aQ6oY7OYKHEbl0t/5bTclF02XKgcJgYcykTIJEifOWKHGU+TGbVBwFiHHonZPTvV+e9RggDlYJuB
xXsW40jjgk2Azs/3H5x78YVmQkdyN+dhh5vPQstQbAgxztEhdbDg1BJYGPlOmbipzEfk3j+qJa/d
TkjH3xopDObLfo0xEjWmSSd8iaNogQULcmJYw/e1LjVgggDKiLiMyWiIUTKqOkmgCrTuRnzgY4ip
3p2PN0TPBlfmG6eGZVzJOClFgl2VYF4wwSbHBLRTONuMc3EzTPmyYI+cOyQi4kV3mE39sLga1h8j
fQIqF1KxoV5hgDo4HSDAFiU/s1fmLJaf5KkoX6QkxusiYrc8c6BGQ/ethYhK7m6OyioRNT/qPviI
Ha+JdvNc/lSPtjtu2BzuHlETwr9W6bczxgFqTaLe3qGpeRxrahIFQECUk/M7HpCpNUtqPc/hnqz7
6gefiXPiLEf9K9xtMcT9L51I5EiP1DaEbZxqhwybO3fkje2C41M4VJewCk0NImtfQ9ORw+IplGDi
bU/auWtT+EKL7JeZgA2myoV1ghg/yIHOuYEpNgk4v6gcxMcDSbB1X6SAd1/W2oneYn8bymPyAowy
49eqHG2Ud1+2O3H26Mf9W2TMidK6DBsoHUzCsOtxf0zjIUvmhqhMXxLaEcW1GkwLLkjy7OTW/lke
lgQy2BXXIFWIxc3Q0g7YVnnSb4XP5sOCbGnht3E+7cTZtHxV848Y/4xuJ4kR6HYfjKCbMag0MTVv
GzP0kpVHO8qye8xQ60dU3Gsr+tGPYc9e7Qs90KG2vZjdlrJK0SjOm/uSf0picBbR5F6u2op3bYD+
tALXo3Nf9TXzbfsNF3KBmFrRI6SXr+qdavGxVrAD98hSK+4bctSbd/qW/3HRHInSCtJ2dVIXpmaB
/oSCGkmsM3LsJAh24neJekiTdXLgkvJmMLafjDZHJ6kKG4ni6L+B2hNHFmf2HY3z8yIgNM4qhgYY
7udgkGmf1oRHikVQjSvYYdFDQJisK7XfuP5bbMGtfKmEEMFNW+Wbq6MQrlYactaz+VXoTHHgjFXw
BnvbgIGXuLF0pZgAwTDQXYCmN/+blVfI3YSb0yfWL3uGLyG3L7lUMcebtbYUoRUCbKM2t09sFROW
yUUWLaVDDmyDfo22A06r9xputtIMf1FvmdrIlM+VN/5eWEi1mUT6g06xVI3XME2FQwg0sRppnzPf
3jU/d7tIAUjQ4jja0vUI9Kx6M8xmqANQwbxk1vy1L1rJcwQ6wPVpflTnzsrENTz9bHbLqY2GdxZP
D3eHgIhvy3VUT+IFVvaXRQ+zExuJziQir7claOkKoXonp4s3pyc7pMv4ygOHUSeBdF3E7BmK8k1p
mjtke1Btb+966nDVjG4reIGVPaisvKeQ1s5vNlpgLbUw8MRtDnYoLAw+wDOIUyu1ZWxf1A4w7dY4
OizkLQ3HefB0f+evFqnqGs7ihBIkJFwkTkPg+mqlQX8zWFt2MJCwGc6Hu0f32A/bmxS1UXcppzXL
N1glo/NRmzTUHoPi3F5XqrbvsVoA+HED1fdoXgRe1JJfHqNTerVqFQODtF9Zx/bbNAEZYZcGkf+S
ScuWg7Cs0RLfD9Fxq7v5TrJJvsHzuIayH9+PBIN7I6MrUiR6f5bWxvPHuOnJsAUgmGCgNzNon858
BvlW5YbG594tlbLbaWCkoeeEtKGIzy4HBl2XNc1fEWE9Zp8oRsCv7YUV/L/HC1WlrCSV7rLxnNx5
O7x31Iaq5Q5uz1XKlpPbqKCTGk9EczZ4pK99NAngTtkqiaOjK2Ys8bF+xrhBoL7WdlvXWYSOkllW
SoCOe8VcN79Ls1ajs2en13HKi7UBwBxFGeojNajgxvZZN1eJK+ZGZvT32tLP+OmxJNzhQCabFEVW
d+ifpClWqVeSJCQSOHBwOr3XDMz0glZfSgKd7sZ2UbPOJbPwvrITIyd3IhUg161rttp4wLfxrqtG
bvirB4tP7jLefNv16bhuVzIaTe6RxjG4BFXlhr3X12y3vLyBk6CoWFdhp8LOX2Zx85DrfL4bNJKT
27YrwE39Dqb43D+WD6v5WTbLCmThpol7NEYpsl2TPI//lmX5PqPkTzTY1sbK5VqqgamZ185S4Bib
J5zNxqqPBk3q6TOikD6jNTLdbYkzbmLnEpBbsSI+i6uJxZePt3qBfUz3pflxH0TotrEHPukLMmZy
P56HNrYWT2UC6CuhULSqPV3k1Ju4HvoNPTLzN0SU5om3LQ0bEN5lTvq8KrSHTsoymQvLW4sygNdo
zG1EdpFV1/4KIZoxcP3BgtYPb4NoAibpuuyIR5J0BN+B5UtFAwoX8TWv10Ipp12clZJXT1S+1aqo
lIPx9PQ6Frhlq5GQ5rB+S4bbQ7ExodiucDoWof/dtCIEHnkvIZEQAmOTrOm5sshc40CD6Y15ZjT0
RLDsPM2gg1WkadOwwmpcwM3OOK0qn8B48ivc5Urqql3hvuHdwO6LuaWOpf1nEWLi12i/SicUfupS
QifCkMdwXK4oYNuIdFFyplPHpzU+BQROCO8QJQRD9jrZ9F1ivTQMbB/3yDVHCB6OtYYZvBZg7nIY
WgFR34m1Eq0JUjk61mvo9a/bNLrPhktpQhSg8KFPF75JgWnsR5/8cWeO1qnTGNlwj9IFBAfyzxcM
zedIxYyFMO/UX7GhLSKaKWuO/D61ZttTTqbb+zv+XihCbnt+WxPaGPugFymBlOh7DvLnlzyuwgrp
lgUKulKAAsohxDGqXrmzDR7qcWlh/evB1xKJwA/lymmAty4TS1GFXkGNq0llTYG8wX92cm3Ti0IP
t8YhQauss9Tmf+HmiShF/CFEQWnut7yZDgU49SyTUL9RKlHpEyLW8OdrxUFh06XKiamS3J5IlkFj
q3a8jfuET8yNC21oVR2IL7/X+WE/fCi9oZSN8ZfB0PEfrPMu0R6rFpNvZHZQIfTtEelHKaL7/V4/
MHcMJ66o0a0uBpUgPlQjfmzKtvSNcL0kNDUbBYs2fNIqbxg72+qQ6DfFFp32gjLWB7AcRw8EVHzP
GCmeYecJihOqrodR6tFPcl63438fyCy6mfMG0NxdSE8Ln7lOdU6prTldkAuFOfTvps3tHqHwTLzf
KQ1gNSW869Uw3TZlFgwahikWtzJIcw63YNHdb/+Kft0V4Bsvt7aTUD6xGnnOBGX7lXQZ2BF0t2+r
ckg0qkzBybKs3brtVckLWxU6xXRoSx77A5RSFQJvDpPzbC1i4SoNslycq4NCv7MAdXpZTpWxoZZE
fGx0P7sTSY/jkUhXwWiiI4w0ydV9AULYm6xaYbLV4dDrwtoIubqHd0A2+OW07j7TYqMrevqV0N3i
yPE5F3u9CN9mX3JCUzPxP6eo2W707feX0VdbkC7nC7CPKCNv/inVCu3Qy76cnUnZef+0UC78q+T6
WJHO9j8ZlBfSp2uMKJgLrVNrW/6gIWPmKtcPhRYCV2n8JXJpamabKoyt/ogU8KHy1CrbA93fkAty
cDAeQ7y2/utSu6gwPK+drKTOpztYkXpr83JAwMJtv8NAbsiomLy4ZlL6t0XXkcHoakiCGOSznPPb
kV1dq8ojsXG16WCKvOGvEvXR2BKITYpHu3oyTc+TRXEPW3f1uwZUwdRcVqDMzcnllkhU3eG65+sV
bVFENv2hK/IuBMj++DQSKgA2QSDPACiNjWbxeS554s4fkXag/sozrNoD2WHHQ8VVUhGQU+Yf8L7+
yYg4zgVpW7Bo6Glbu4I9n737EDf5ZPde7gYi3DsaMPGDHjToCaWBE300ggPo6a5V5qaN2t4FrFs1
NApYCTVQnGyHnbs1YJ8eDaNfUdkB/QLU3OW8oSQ0a0FHKl7iUCNnl+MSR2Nm/j1MyQmLj81UYbub
VJ8LKv+WjdLs3vFIY1E7+hqHFOhL/HDQdV6Rh2DkM/rC0Cg2eEg+GvHPQqF6I0Nvbekc0dILBIqb
I5DNBW+46L3DqZJbbHeWDXbIVdrsZBhjMiPoBhSfBnRWeEpuuSxMyQ1Xv4QRy7JM5AvkcJEMvWqo
/IyLjgAo4FDao/WHNAdRcI/HVsRUntQMzeLna8whASo9QgA09RSd6ZWcceQL1TWgwKymI9I2adGa
nk2gEGTvkDO9K7a9c3PkP42rOnVxmH6uXf8En4LOZTBWeFMhytq5weZHqz4t8i5/QIFE3pUm+Co0
kwwL2fHuW+yWbC1t2hIWgtqUzqzduETRWe5JlK7OEh6OVQD7xp14wolHtpmJv6dWH/SIrP/kuXNf
dFDYzXSEhRkhY9mmmgHhxoEXEhfhmABysx5FB9qropWHp1klzO0VCA3scwxX4nDLi5Uv0ogOOClB
8GNxfXh7y9Oqkdn+F3kdCc7gWOO2UV5b+c7Wlp1FAxo+V+oQYgXCFak0B806JQkhMpXg75o5yp71
fivthEqYvc9cho9z6GbNZX0V+dKw7krtYyhTDfYLaoJTGtH/wlt867LeeaRdbWhMeuSt4eRYsnno
Vvac2/eLCimBgWNKadz5T2SUYzJ0Urw1ysjDVgsikBfnXoAmV4tPBIe8Mavfu9KuY+0ylIra2qwa
uneS4PsBsjMqxnVc87NKvyzWnqkLtlfUXRTPGVqSaj4337ZirqthASJ4zSMw/tHUWtdcIaSX8e9H
yyetG7VR+yVgFk1X6hNz5ylR3tG1aemjA3dOBb6IVrjkZ91Y+/x5nuc7U8zF/DZgwsxCJASsJTNA
obwC201vx4RxVIkMAwQDbW2MyJM9Gdr8E2U4gyzi0GFW6ITv4osPJI0KZugl6CLrsVj7Ztr3X93r
9GhO0lGgMbmUlJ/MfMjFHS3Jsn3nBvZBYYqpZ0zdq2jzAscWbSBB66/goSO6CeL73f5Hy9UuA5JX
eM61lj5EWAmPDe3k5CZll/cs0F4HLnEIZn8ptdQp402e7IFZ2wSgpbHU/YHsfRnKOSfrELW8xo7C
KtbF6NeSXiYCgljfmF6pYi76Gg0sPYEh1xdbZSGNRf8aYEgyn7tqwwvepIgMk71yjB0RiceoE86w
nyW4lcNjvhRXDz2eajxfVkJMVQ8EiwTnv0310QNXYCW9WCrK42ELaBQZIin7vr3fJftseqNeQAgW
eBgnRQdqpNCiFKsCh4QM6SMMjAtDEpI94UaiAG7+TjnTzWIOl5yKD/29HLRtEotVsne/wyAPu0xR
04qg6NgOeK5oPnEpICg7Fsi5fCObRZbhCN1LOVcYN1QqBweQtVerNNl2tkYGYw3zN5rESkrUKfsK
UUZlVC5SbJkL9O0hFYB3GCedr/tWDeW5IuoTwniSqKmlY0086vqlVdtO+1Rva5H5nvw/mHF2aE9r
3uLlG0qbwJELC/G6hNzkorcjj8sS49VKuZ+osGG8EH36OtVLL0UKcQPePoh7X5DgDcnNQ/lC+KdV
6oilSzzZ2DLdDibyXrF4r9d33WLiwLI9cCiP5U7+AfjIX6qCoDSYt8Cd7QjxBJM4YmvePa+5g4K2
gifNqHdEjlBIkEP2nE740m2Bq0Mgl6BZm/gnuUekQCr+7pg85uUvA9eKNsMTG4mcD6Mj+C+jboVf
XQo5CY1fBtuYAq3c3upJcidjhLXB2rBbORWSQl8AnDbLWw806uHgs1rVot5p2PrxZaK7bKmOyeSO
/4rWKRvt/DAEU00iheRy4D8WfDfjtvb7e4Fml0mEKdPwvVuPxqVPbRq60J+vnJBEJb2IuI2nFZcs
y/2noaJ6tp4y4zwCVD5Rwmr8/vvisehNYgJllbB1L1gNKyiwr/Fgp/Du5OQgGTuBtbtr8a7bvNtl
NfwT0rhCMEsHX8hXkvcxa2FYgRRIp1K5U30EslaI90nhIcKipES6INzdNT4b1KK8jO1DjTohCw+u
uldhMi/03AUp2R8bkrgumvhjFfk1mQGeoUaVFA1DzZbvQ29712cFhBsPi2IRlvDRbjbcd/Q3uxTi
j1Nxz3WBJOJ5/vz6XGIUBGMxINVYDAmbGAtT2z4CTK3/EaA6xmNTbzHTlCGq3nealiO1G/LNbQ1y
iYvJ07Z8e+xrtLlieGzwBbYQeYs/CWk1BNcOVc8/3CtlM4DmaVahHx4X9Ru4Y4Yg9MT16AIKFsWq
dBe7XfzXTZepnpdWmlRcy8eXrBgrkoGb9PeSluTiGCXUCnRAxssFt2YB+CTh9MGLp5Xj9DFZQpS7
GPIDPodIUDvwWfk2ZPesQa1XyQcXpyDPNr+IUHh1vObc4RiBmTCVL9VvR10h3yUQ4qTvFBFLX//S
YRKst5gFsBOYcYYtVRG/Om+VbCGMKGIq9XZvK+/kJ3kf4mjiXES7PHcsOWAUpuAu9kJKWAKJ+Jq+
YlOYcie1kX/O56caLTuyGK3oj86mQCaZ8BzEn2Mf6PfJbgdaRpl2XZnxXxHYCCOT0STK528wmlAl
YXM51BORs2om60q8SSq6YrDc6JpnF5VGwBb9V3zOGlaEhb19M/d+jNHTtJim7Wg6Eka60pdz7mJm
fh6JkbvNvPhVXsVj+cQ27GJlMT6hUbix7F9olb6YpdamMRAz8aqHNcUYw22uw0ojIAj4JNIoiqZ3
16tz+fONtR0IhVL9tVwvtqZSQJnh7v5SeFusTR33HPgT8D7tQgkjiy6xe+GmBsEIGH39VXk7qxUW
Twev4VSZjByye2sllblQCbhtkmYjIr5Pn42VrhuJspeRYkU9bdPRl1y/gWAeQfimF0a+mYN7d5om
2N1xxFz4K9JMG2EVVUUrUSs972fpBhfHRmLy9p+0flCYKiteAjXOt753ROqx8Av1zJauurZDYyj5
osB3Au282xjkCaIi3MQ3trVQbWLYS6NiuXNxMDdlWl8rK7e6dkQJOK/adRuTlbevjWu2w4M9dSyt
BPhM8AJ68/nWoemu+k0QWWHeW1T+ep+NELlNL6rP290bJxzW1xwSrDlzCG1onLFpmOwcn20y2+Ih
ERv2TDPt2KYD96yq1m0K8pXn+El/iqVgJAHj6sdchGmfhsaAakF3CKzOtfWkJvV4gz17LFeZuL9Y
hVnxp6xecku5FBWIXA6xuNInXT70Y95hlyQMss8InxFh4+SdyuaU6LOfx9flF6TE4QODet73XB8S
RIUrPUp6QzpKkrjGIDpfgotHf9+kMAQhA3kWOH4GnxLVHcInaNeGT5UkGCeAVDD6VbOi3qNVSpKA
Y++Ev254eBVVrqWi4oYUGJm70yZDdLKBN0IAWd2N1IhQV+S4m/1rwxuwpZl1csYB+bZRoUKhNrJZ
nWRGDF8A7eNyXjLI4D6p2Qq6Sad4gwVlC1QPwPPJJi/K98BwBEruEOk6D2yElISkXwDuYYrJD3bH
rueATNOMw61JX4rdwoiQ1IrBIWGHzbP+9u1fhxoopdBmcF71YDCii8NRAJlPapl49iO+1iajOREk
qdw/X3+WX/PWt+f2FAmNB/FOy1vtoAY3u1kq6qh9nFKkKK83Z6/v1TlbcSWTwPtK7eonPR552XSq
xvDeT0ogpTS3ub/ZiDEU1xWPvZc632wx0+VyEtl5uI/93iX5UiRYyCQkoYzRQHRJPyqI9RaLA9vz
AwqaktYkG/F8FHTM9mETb8GO3fBtGzAX4um3Ak64qNGL/Ki7qaZ6CSPb4H5M6kMtqeRZU7RXtMr+
ALGlzi0YByLrZzbM9aVPnL0GxkD0Uju6INzFsSiLveyQ976SlLM2+SYIDkBSTT+fFcmY+Rl5z1TZ
wPsraz5nuC37Dg64DYQOUkOwmlRCpcXbnb2AdJ4DpTSdp8+c7+f0XZqEWIR+a0AQMrrPsJeKlk2/
mOMefSMb5OJja+LnZwKiIq8tI9WrRl9scZ1+w7W061BGnxR56Scv3hUUDHlHeIbrOy17L0NiWQXt
bQXC3R2OfGow4P0SVr97AZXgceRopOxSnn84BxWX0Tlvtz9j4JR04ykQoNNy0ECRw9fICoBQ7sNd
G9cbzSE8oin5H8y9Zkn5IOKXcYPYT3pHaVLFcQMfwFoooSFdcJZI4gLqyQaPPcz/rXfwdrkYdt8m
+OmMQvdd3+/vyCHRVjxV+lcBkw+ZqNJZe5xv6EwrNaSpu68FuCYBnnBQY/Y23vuF3PkBxTZfQLU8
TpNQOfU7lB4TuwR12H1VdIxTS5jeSvkoERgQqURknnHkLrHVx14iEU81S+5igpLcXyqMsA8NXFIR
5yH+ZuSaTqWTmQYkQk90Hkqnf/uSZgDmz1JtOnOS09GZLmPxw1fO20D6aKDdXhyUMnvROwENwIb4
S6dwJQQzucJMBIoZlO75K+lq9zIZUcZFT1AxKtVozIR238Dy6ctSKsgRS6ADLO7qJzdThRLgJMDQ
MdSKMtkx2YHBf2HcLk60gPI4hD0SkfyMUBQ9Z+cV7kT1VNEutH6LUt3iwd+fp9s40q3MNKD+vRiN
IL0EQDaUgdRBQ6uI+bOTC2L4IAeT5b1Sz55AAdNv1/Y1EF/sE4AcZzpRW3f7VxWLkPHU18hrzwb+
t4qDaMPaCRWGgeoJw885TY8Jb1q1miprEq7vSrGYvkDWlhcGI4HOgzsSL8axY6xgEO4TTYLyGl5J
7vra60RLvXuCnSxUf1YkWHrrwnR+jN6W6tpJDsSf3V/d6K4OKLf6fsI7ph1MFgFZUBDMrPs62Z8Z
lDQM74EGA1EapvNpEXNunLOI89mvvExuNwwc1tAjv17nN/FtuyTAvZuxD6rDUk+hZbPTZ2XjM/PA
vpc9EPq36WFtT5bZj444U7h4CLMi1D51Q4pZ/vCKJKm/gWA3XubKMmM4JHnRK6Cc5+Yd14N804U6
VQCrgHlfH01XnQqH+stAOv/v2Y+YS8LIZ1KIbrRA2YzlkY398DywIzyiNOORNXzEncpY3E4N6Xra
fgSEwIFljy57JN++JauRUIRgYhFvDgfyx7YFCUCpjYpCVCH+BAtFS2Mf1JGxEWYtGApaBxzcWiK2
NJ0EaPFGYmN//Sls/4zWey7ktBhDhRW8I0QRVdW16791fmdwaaWHEv2eG3znr3NwBeQk2WW7usgH
efZbD++9z4F4dvSxTC0zevhfSDPis7U5ZkGx+Gwd/tD6RYBb5VvjC1OVR/xfeeRr9whba9+Gm0rS
296BP9Cr3s827M038mfXUp1j8cJpQzVUdPb8cLtjZ49FVUj2jvejcT2Ty4gMhAATpo3O6FC1kZCn
qvEgYSku3g/FHatW0nGfsusQQVVaHoAvn+peI/3tRS3kvorC3mg+HWtnb6Ht6Q3kB8IGBoqv5wgy
xM6LDfYvFyfS01oSnJTAAuvTzgWzzSNeqOdqxEL/4V/nX+biunmUHVxxx8jrteSx88+N1zSYMhj8
tHj417k7xLDCoKf0TWvWasvGwx341SRRtltCJWsBtQLLKcHzP4h0onIYQCcpDjGY2iu8nQBkQ7A0
K2GIdIxdiR8QNFIbfWxnVeiLKVLfLfDdU7pjCQLle2WVxRwlE5tMoP4yuc36V9jVqMi+fRYUMe8o
dCUc3fNGuuDpk5k/qYWDkD/ibMmJj8PconDbyYXj2aWMoQnfIS+PAwP6BPA93GPN94VPQRnUTTP5
JsuS2CAz++EjomwW77yUEFzJPXpG0kMlbYy5WuVlaGr/6zm5CnfrugLJxiWW4vgB6WtcBf8TspLs
dYj8o6kYT6S/7Q3K/Oht/p1jYGxiet5cseK7hrmZ+DH+nW8meUXZUMIMqAU9Kz8Wgq4KHE8FOkuR
ynclB5fCOCgilQVEePfLuVCxD0V82ULK1tVffJ2uIkYGM9CgMoJwxpWFtK9GaSoGOR+bIjt/6mNB
8eFLAtossZ0Fy4FE0t07pbvZTwKA2jvJ8skiKBOQdw+Wnd+f1QzaFd/RzaROeqhgKxBNQZPJYoKz
W2yy4zxB47oav0RSTndneQrpl6FASXHduIVAQrrTlDbtlaI3N9K0qsddgdEIqCgifaDyg+2Ah446
WbXYyhg/MAs0gokB7KQSaNz81ApTkULuc8p2xyvFqAYLyFdnt0eTfOUQwD3r3Gpoz6K3nFngGsy8
lvr8++wUlY5LhFrwgMUW2GganmbASC1VGT58dD5ZvPtRug9xGklZzP2dGv1pdVk81I4ajJ6U+20M
W6FEym2y1Ae8NUA9GtIg9X0Dci2yUhQxIkJXMDZq7iSJcsK+EX6SrL5OUYWqLyejHPuJ/HaZi3Z2
1s/w4tJx1qLuK418WcgbTLCzV6UvjNA/9GLJwx0A/6Q0OXpccEhaDQ1IiF7gJ+EspeI31dNxVZ2h
bgFH3fnnPOSxcrdj2eiwXE9eXpOoZ9UZr9P1UbUX9PcgXqiIYR+NLPUEWB7yhBudWIOjISfzrGwT
qibyVLMnHvQbjfI63aEWjJGOmptzGo6HZCx2F45WtiN5nui1m8AmTFHBapYHnl+JQQuRaiSCy8Y0
tvWi9iAvwctZeqBhfUbQAyN+GBMZ0vrjiL4UFRwHEpY2OsQV13CSRSTtgnijXCUQAJcJ/Q0a7kcc
yViLTv7gG0/Cj1k0hLkhXTplg6UvSZbo9J7Yg1rs1YPMdQo+UI2SGYMffpBmZ7lOrJFIgU/Vkh3R
MjzUMlDfGltujWbEeJ+hCXaySSY0/bYs8qXRYxhE42Og+W9eWR5ivIZSzhGUS91iUYhzWn/n8DC+
eN4UUVs1Yvg9Hpy9SzNfHIcwkG3aTFNwhu1ZR7fF01hW3yyReMF5CdNKrdVm7mu6bN/BfeY6sYTh
6nWWu8kQgNlrhzyWlJ2Dt/k9cogLC+9U5vFzMsbGxfoyNcnGLtA3OkgG0bt7XnANgi20TUTFKkMY
CYd7pLu7Ic7mTcyvSMkHJUbpd4X0dzdNspdAmJ9wke1avsl58igaXrx2+6Z6zUJwdHTZD0xmv63l
YeJ3vbHYpMtf18LaSVgzTg/pFjSmt4gbmd6mBZ6x7+8fLtxSACyAeopFKflLLHo68+jthMwTVuPm
jHh377EXCia/dgnYFpaYdlk5Ks996iRoox83FCqYOMlCFrGOc39gifjEIVNWzJrXIQTPMRRG31L3
zBz77d6cxVAj7Ul0f8HVuJwtzTw4dRf9so3vWs64w0KqVfn9kE2y7yUMenBJ94WIFpNpMO0FcPOU
pIyZfbOmuhUazbk+GmJN26cHcQ+rcWCmy0DRSo8OZjhHRKjTasu3wojZX0jIKpeOHYGp4wiFtKg4
9Kum0LKBah9dOw8WJSJV4fOAgHErQsfS6aX2CeZ39goXvhNy6NlX1FutRBgOsFNU4EFMkG0afD3+
j4YYNNTIaBSdD82tA0V9I63xJVCevUb9vxrozvZoiu0ULqmGEdPBUS20KfMhXowpUf1zCPnfdWqf
cYtb1esIThPoHmcJDuVTWTMCQfvtUOkO/iZS1bYgU4ysKFiZR/6QYZABRpyphDooOqIgHJ8hjE6t
dUO/C1XPGADySj6Mt2f068lkOnFCaJGEzuPFeYCL4TcZHj5V3G5BRZaKk2K/tMN938FZcZ1DpT0u
j7Ec2A9u6L9Tx+dBM0IbnW9StwGGqlR2LANEBWoVFpdqaX8TjPXvCEHYljAAMGz50QFAlqK4XuLD
9jBeONu/2xW1Ky6ScmstzxgVNCUOeKyKx0Xrcl3JDOEqXkZHgwWxxFtDoirqnqKGd2sZ1HuaJ579
8417zAXC/NCfkfN9eQdFpoUbmU0UmYIOENMLLHUL42p7stAaJoHzjitSpEwuHRanWm2w3Jtv3+vj
9uv6+Qd/5btKMIDDM0ygAWPAP3rndGjSllzvtmZIkCWfWcgZfvEqxB8hwOIDMsssNx6ps3evqUSR
Gq0ZDxyFEd7nd3/APpABn3GJrQQKuDq/A8D9TDOWb0jmnpdGthCdYVwTcoLklaWo+WdsTFT041ui
b+I0sAgPeIDr1w8kV/d/nzcsNti2Umn/AnHoQfpjJyrIlHIyy7PxGcCU5RDo1d416T7ca2WklE9J
PGv6liIK51Gx5VH/v+kDYxmjJXolPXvuhXgV6vx1nGJ3tq5yw+OV8bSfo6U2mmwNdIYtDgvh8quK
1YDdc3nz+7HBszQW1CTIwsUhlJTWoRwyEwq9FtpW4jwfHV3oSEo3jLG+z+uoqucPDKCplnExNJbE
9ECr5xkk1yPpxNII7oXK2jI1t89AxjHwREWIN7ezs3BCvBh9lrPC7Rf+V9IC0TyAIV2h4fGhu4bT
+wZbdAX1Ev2exuL/VlG5dge0dmqO1fMjxpYvF6feIJ2AtzjfZFf//uozJ2hcoQ4aRG1ekybYQyH1
E3FTG0w/PYBf/sNS/rkEEaFjLP9pCINpr0TbvjZVDF7RVuPwwKNZfqRwq2OA6CI0eVQteSxLIhPw
i87feJdpUgrWN3GecibVSCsuOOADFsOXpg46jJ0XbhmbrsvKtJ1he9bTJlAxtIHRZzK1QT1JisYE
w40mL2wsi1mz1i7aaewp4+w9fCu4QUFu3PgqJzk2aV047yuc79mhRmJ+1iBtejccjpZqTB9pczDE
fi+B4K30qkAysVREuEa4uPvXiK53AD++LtuQRKXevjaQCIsF+1i+1VKxbHu+3MoojLk2mkf7eZ1y
bARkNpcMwGGOBKoewrZctC25G2fu8530VxssLFLTN0dvtZ1PrhHERp5z4yjrIXe1YtyZgnEAOgPU
FJAXvtZCOdXHIu9laGTEUnV8NOHIZQM86o0IVAChlB/Q8McmdGntusMElWXeh55nlJucQcF80lCP
g0RwIOrwLp1KYtMRO9o5h570B/hlofWfD4zMjSwUzju2NjmdtcVOrwPi4vToIDqJLT0OaAE4Pm4+
MMnjmIUo/SFWAn5QNaN722nw9fqyVctbGjrXKV4XGFQALQbG8j7Q/MvVn1LqOiIycvrYBKNwIUPT
2Tkyaarryv4eXuIK3gyY1BJtHyhVUGalYXxBNP+2BD1e/mL+CwIt59DmC7A9s6j1M3xjp/c5SgLj
6mV6laA+XHigjYWSoR6DP7mioAqVj80JWEkijvuwYDQX5na+50iSMgwbiaqVTsVf8riW//kGfM1K
vjv9YOIq++4kYqyPs65YnSA6fjlDgT7a5EtsX6N+1If6pARbfInxKdaj2DuhMDkueBshW9YOaRhJ
Hj/vNRts4J7so2et4sl7dfwCL1ivMoMmNfoKk0nfHTn5DCVDC1mLNXTwaZBvJ/Xh5xDnAEaCTDE0
3m4Gg8LuNBHCF8oXJFb5nigWkWm/g/b9CDOuDT4/bO2cGwLXmXMp/54172ebV0zRKGoH161v4/wt
jNcjR7NdN2YQ+wGIPywZ4OaO/roCsAglzhabefvnYA3l7h5kx4Ka5rUiPsd6dS0De6XDdh/4nHWX
mDL7Vc7snZ4kZVyBiHmWzFgdE+mNf2c8vuh40cSIdVdTkOff0jbNrgJ3QQ1dubD2BfUvr7609Su3
UjG6Xi/WSEmRKgoXgleQk0Qz2N0tpY6oTLHjmmXsdfTn2+FEIgYZGO6UAKP/s7nVHf0UZi8ysp4F
YsQYIu4zGnxuCXP9KPEDeCPLWiQmKRGuCl4M4r1RRpAQLuH1Qr12FpQuduP6sa0tsbSpOzjG2UVy
uWHqDK7uLEd8gsz/GJarTz/6Vnln0u0IVndjYuc9/ga+w/NFV5204Iv5SItQLCGiIIUUMCEI72PF
VcWZrUr/nH7fGioC3ycV1JJDuaMR4IZ78RGDjy6aMuSECBvwj82w7xbFufK/tnkB8ygm4iOktb7t
3fHP21woJkRhLhYyq4X+GCi7rFWjtFNgAeuskNKBAk8xX5ewBx5Hnq+dlokjzeA7hXH+yCbMB2ds
b+FwpSCZuKnWHc+Dd3gAfC4jAMcX13KnzpdzJ6159NXVwXJV4paweBlXyQhIvSqDjeCO3V/H2uWJ
shOGP6FahwiftGlofqNsfQ3p3IYej8bHnLkHCOU3FFxe0Lg4pghhFXwevvb36XDvCnujkoHEXeZK
6RPwn2oBHJzHtN4vXH9T5CyPtsYMu3zIhimKEoPYjMYRppobrD/1YGqhzDRUoFQNWW63jejBc2la
/7TEek/V1ojXU4B1sYrjStyU7JWgtBAyibThoqcTIZTpWtiMJGDpK4syKAlADO/LlAxVixqX1JS3
fVFCxuHxHS7gjFYonggBcH4rmPvUCDKeltvGwVz2y9nUZDUldZcCV54WEWha7l0r4Pg6Oe6QWIiD
DpDZoZo0fFmsuxaPP2e0SW8w91NUflp9CQAFHtMlNxl0lYN9YeE3dyOUMy6Dd8i7nGYfPXBYlVH6
aXoitAEwrgim29alnGJINIO1zuNO+k+nYpnCtctFBg9soRYHrtmDvrp9QytOatSPnnYGC2wt+LGf
67KyXsjgHTN4A8YeGJu1+kBTijzCAvW7rRWfcNwT2Gz31RhqKenvPHc/yEVCFBQbuHkcfr3gwahv
QKMGMvlndq2kiT0X5feN5pcL02OiH2EZ3ewkIyDLjBrdAn9mlW+ZvL7Ft3vPZzL03vyoaVrnP8N4
qjmaAbdzikOhv2TI0Jh8YpwEFtiDIf+B2cYVZyQrVz58lBu15vKB6r2gzey1+Kf4JUY8xjsTs44E
3mSQxfu2QMpTnODdeW8L2SiN35xUfnxN4kb+lLE8KxNowHcsPYfkHdBqPiUIU7XvOGmYF56p82dV
k3v/PaK0OXQoLVivhgiXJ4oKKWAtp5fuQIq0t5laf++quu2nYhqbttng4uJoWTTBscWb/uW63zm9
S9cExMZZGM54zFJGuNUHS6j4TF9UvgDfUz41esn6dnWBNDC78UKRd4YwU3jZXem04qTD7zvMMC4f
du2buQ5ThfsxkGjtg0MkjxuSvjtA3Tn4wM5L/AtDBPRbL0CMPQEWZ18AsC7ZMgLVz//IOBKvgr9/
elaFPOOuaqwKS+vuqxjsvTQLlydKvr5sqnzbvH09JBhq4FjpaNnQiuRe5aEqVhsVvZRqRxF1G2oe
NKpyJ/ShqLm9GcwRTiBof9hNyh/g5PHOd0sVaoVNlNx5lk1oA4fzasml5zmlvvDmatJuiwN/Ikhl
5pjXaVud9ADTawps2rfFCM2slrF6DWQqOsG7Sxgj5VlZ20chHpyzXE76Qw5tDDK/e44Pd2t9LGbZ
UD6xmY+0yOyExhS3trafJXBYRzyXX4y1pGDWPgENOow+4zVrBKc9a562OXQO6Z3Bubgl7RjmpGnL
vm1eLhVhyQWmmQ6m6k+Wd21gP+Po3ajI90sMP6E2SQPpCpAdH/sIb9uFyXAN+pqmpRk6ncGqZY1y
PlI0oT9kBn+MEEWqyXRpOi6fD46dUfxZglT6tNZRIafjKy95hNOFmIT9LQD9zo7vmhPOOBihgC7P
tSfKlA1bBaV6s1qP/4oVW8OzjtgxMYUcU3MDJXC5mLMWBW+GlRSsJEsKCBt6FTP8xjEnZh1PZ2vB
ppqRVjQaPpkUlpVpnuK6rufMZAyZSNCdVTjpP76U7W7TVVLzvRCxEi5J0yYpyYmzuwNtZkBUF5lX
5Pj+nzFEFjrkXT2V6Zgezrkxzz3Bir2ZJW0UGuP4OzGVQdyjCTmLTeFGhE5VxFtv7pUDAHAw5Ap8
QvG4AtN5LTgYlOeJEvTHU+Zjv8tI8VgZakaRrGdPdYQrHWumulVFgxsFRc5qTk4H0w+36vQyTPiI
dGCLqXsb6BOo+IwQut1Xz7XoGZWoIXwuicixDKZVbDTE88Y4NcSp/LTfDn2wcflGYy/YRaCvjAdv
h9JRZD4Kn0wmJNt515L8CGAbJG10FjKnoNCwiDNuYgzCW7o2l64qCrf/7L+Lvt4wGrOcVhj23TLO
4K3Xk0WmdW7BYZZIQKYVSzA4JEBr5QeQnG6STSSUdejYhN/HfuYE90+gpEAI9UIo6l5fiimN+fqj
PY6soOISAG5uC4+TsS/+c9Zuf2JKKA/9UbEB3KkQoUnC1zPMevSeM8Y2B6azCUv2icyRWankw+RF
WAnWsu4kSEceh6XWnf9Gh7FUvQ93IcXAR6+TkxwQkngzHH3zlijGRvZVRgzhoWoJcpMTvROXMj/K
KjMXJequPdOwF4AN8WrJLumQAdZPNhpqhZ49/IOObaWU98mv/HOvdjkVu7y/tQTq0DDYjApdr2mH
Di3zNJkwek9WQCT4jTWiwPCZtpJbEVUh5B18w6K/6YyrqD0SmMFEiHAI72LoQvRpTzUIPl2NKSqe
qrntHVaAJevhG9OYG8lnAKCYrk4o4bvriHM+U/jhmoXiPV4gIZrs+xZtACBEQn+07VrjfevsTVmf
DjzRj1JehwwLsqu0WdbpYNbCbX0VtQd0oAeQDqln16XAc6T9tplc4+260apJeWx7t80Flwmy6Yw+
JzxFonDzIF315CyXp1G12AfYdeUhNN2bqJ70u1Mhf/zz+exvTnVyb08xb6tnaTFQDNlcE2vCnqq5
2UiHGTM/ilmvhm4uQCqe9MsrMe0+9MJUvhW45NyOxbeRIapuvFSVOJJUhiEN+0CSh/GmTeVd0u8Y
5qq28pb27BYqQSKqgGUoLLL8JXrGAuZCuWQgYTzTTTygretR7bIDUDqyMFSpDchpu3wC3rPhn237
o/8CSP+6724wIRIX4HQIvqU1obZ/g7hEtB9igNdm/sgtAg8i7TxfIExMPtLcThcp3/zBdXbdm+cy
yel1+uSbVe7TyyyP/U9ypwC0vd8UU7HM+sZXW40pho1H4GP5tzs4BQ3pVOAq1++TANZqbWkSp3UD
ABFHbxEzyOqlo4H7d+rCCAQMeQGUE6RwgVzJ8wrbxeOVSjkm/niZunAkIQK1ySS876+k/swQDLF9
1/rbBKSUN/G2DCyMGVDuAzrlG465TH5X9yKzF9nsyY12rYpTCCkAuCx1AhD1MQgtmCzv70PDmT69
5UmJg1iUaZkTSXxVtR6kfPbvqN3PvB0b/HoWttrfUiJu15mFEQseGb+vss3XqtC7hSaWZMwimSUo
oVAq/PhRyqRpeXbPOu1KdD0dm8oPxkB7osXVfSZiB2CNYv3KVT2KBiLcNStKrG9m7o5YDyNu7hy2
28aSndXBbE3aRI3tZmV98taEvRvmS57onSur+p00BjHdCsPpEmvZSgJrJ7b0NgpKii/LV2Jj31A4
SNC/yK9USAJ4YsiD3IcvJK8cmLCSVOhV0cZ583m73+R5oaGGclj9wzGMlNMoSAiQSyU9iADPmvuD
gR4szUq0KH71kigaGqI78O3DOtBkmUZpCfYqD24N1jVKpH/i+iWa6r5Irs9mJbhTZxsysmUgW3Pk
fL3N9YST1JYy0P9O3pRpC+nbCm5AEWmCWBZs5cyK2emmoiTy/Bec4QAibdumqOKxPX30U2gynr5f
d+Z+9QJrTtSFOUaCthAZ4TQWumgoO14NACl11Thotju6kJCorAhJc4OlhmtnXe4QO/CMOF6oBsko
dBINwVjDRgAnt5mo0FRfFj6AUmOor6jI9zKvFd7Ewd6WyN8vSit63f8pKv1Vd1Lj+X9W+fWlkTo8
HhbAMtTyRIbKH80XPcVaYHCVYzqvKxkpmB5DPIsGASqP4SMxUby4A252u8OR8YEEr9QIC/YOoAF9
KfQqDvX/B6hJVJXSKFzEA+oQDXX31ULqdgosKfLSMtQ5dVyNJYUXhCom285X5gWH2RCTCxxlP2rO
Lr2xvymCg4PfNjp+Iw8XXBtvnBDPatG+G7qeCOaSTKTOR/qu5PYeX6l3x97rZgLKhmIHcjVxzlRl
x4RM0u0JUFeNe+5W/8dXSM90dxyTW1oZUmLRe44idgpDoWCPe42p//ZucZlG0MZowLHhFPIXB8/z
qzy7rkHWLsSQMM60sfIP1uIMrEhGDrwK4hyEK8BTQXoBRerWp1hHpjE7HKDHzPNeeRmWp6bHqjz9
x0+9+P4bxhVfoKVD6wOqnjYWpec3kOdLMLIjaxcI9AmOCqxmA5gQYVmV0tvQ0Dpr2rgltqwK5dlc
gYTyAvoRb1/NQP52mYLbUo/mtMeU30ELbvnv2azkFUuts6JikKAIT2xnq6/45oHCl58jpX0uCurr
2Z7UR85cxkePrwqHfd2I7i0KOYpDZ07EK4LFrqFlMP+ybqUtcpuSGdiNG45uCr5IiP/+SFY2GmKu
cn5tWEwiXTtVx3TnRQdVYajqX24LKzTWBQgMce+9ThpwJfJUzkcLTHqEkxXyvKPK6ca4ytckaHvB
r7aloEJMJ3czUaYtQY/KpdQbxW7Hv0uOgepsBSjL2KTKoYWpJxGNeaB/Qc4EwKqtepxd1p6C3C5a
/+S5VWtkYgP2GmbKV3ahDRbCN7WBtuPgYs0oePmAh49lfBKdqk7QNKMLgOvuAsIttRYQTYuWd+uR
DiD1/JtT6iWN3RHeQ3V2DEv0pFE/ChisYeMIZeM57d0yocM4E4/n5Kl1hJCqVWMSlU5Arw+rX4VN
41531+atHUuxlTKgWzUEeoQ0lP7AkYqwUhsj09DGY2iYe66qBhM5Nl+Uv6cgUw/N0kLJ1gz+NbzO
SnG1p/OIeTyW3lkvd+voE+4bMLpZo6NM0yshiLeEZy8e2UnNClhOrRuVu6DyyndVOslTbohiuaXv
lFwCIHn8/G7sRkFxpGq0fEQHLh574Lv31YiG2PybELJ0a8aon//VH60MRpbMbQFIDRx48CxP2kZY
cj58EJnN4uJuQI6wpFZajdo1geRk3pRPzFJgCzs/QkqKu+szgHqnx9CfLQVQUtmJBJLQQuWvb6eD
ihxAc242L3KZDR8BOMhO+sD7mszvD9BdEsjB2LhWbVqaiemKX3exf1zl+QjmA+O6vLmEjqT0KwnV
aRR5EJJu5JmaMmv+s4/uG/6ijT7bDetr87rdsRx8e0JWYEFNYnmktnQ71m+DwttG745dGRjYIWt8
eSuqtIzbY9+TkJ3WPrU8qawFHbsBhu4rBjjM9jbLI95oXvU7/1v+22haFvjpPP1ABjy1pQaIKvwj
WIGKtZ3j0khmekscCVZLgcRIqDrO47GmnD4wS8sWSQGo3X+2U8zVAIEmTvkxPuA+WlITCvO5bdo2
U0/dU8KKHZJN9h+/AR7CFUedZZ70dK/IiQTVv1hixpZp+jQn3OiHojrwOlYvAUYSRQl9ttM8SyzB
yuxy/rHi5mvWsKFrTcDgJF/vOBl+Iq18kynKyMsh82R1SzONQoFwvwr4Lxntztl+5rcGmDqpnlmG
a5zwSPP5sUqJxXLT0/rievXZsz5nKcS6VRYUZmHNCaTQr/1o9t4SP9chOadCQYCRTBYeZh3S4I5w
HVSJa+CxmTuzc+6wZh03SpI428ODr2IB/y1LXJNrIXdbFYsTaOC/f/sdtd68BVNPKw3cL+brmZus
uk9z2PzhXeTFPdl7gculMOQV3iBEvilhe1wmJu9xSZUmvJt5bpw0T/lAkzeYQlQi8HG/7BBxzeVM
l4OnMK8p360vO26gSLbEIzv5+pZQnz6szf77VIhJbvTslM2aIAX3ef3q/TNIJ+MQaO34qiwF9Ot3
KDV2dFOz9Klp0E0m1gW8rAEbJ4J6M6t3cdA0Og3ohRcRK9eQVnFswl0Qip534E1defSZGygP67Lb
a+vGX+PVOojbbrdKVaHpIuYr16HGXEMxwnDyUnJbnw/JMU7wfnCsvEnU87QoT1W8qOsjwQGXIWzu
oweamjL7h5Q8QvtpTTWPw0cvazetb276mx5qylJ7lzIkkEhXtCXdm7GLK9NZWyZZK5ScVN6GAAHr
eu2DvonSKs2WZYcOpC0AEtBN5bjKFnlz+rzrYFqYq6vPTHfdKrYjGGWM9tLXZIdDpRMw1kqa59LJ
rW7j2SCayoNwPIruIObuWmaC0Npi0yFwESJh6+8EiW1YoxYA03Atm/9U1OQpkjeJE3A1/Eqn7MDF
RMJ4Hn6EQ2z+xbikla9+sV6/jaAJAQt5n6pHiwEiwojxBEcF5tc5Hjpdc1wfNLnKOeU5IBqXp9le
4axDzUO84ZJ8YQQA1Q1s74vl8WqEd5IXxW99A6AjMGLSF/jArx7HKN7DMJSOOnHmpfCIfR9ZXq2B
5m61Ky5Q9mZgsc5RSz+prjn8hUDGkIajzLktdXdSyTxehRhLhXqgzd+l2f64MLtVtW899XxRk2qE
aOo8XJ+M7Ux5BnWQoDJ8pWvGLYqUzO5wKhyDO8S1MDEAuFz3z4cB2XYST5v5iqx6rP2uqnEWcn0u
+fRkijnZhiPqC19FL9eAuv+J4wH1AKEGx0kafwuRzYFPmoh9+8CfTTCyt/FFl4AJHAEl7MoTNW8g
0HikX6wFy0cM1k6ELR9oWdTwizoK5RXkrI5KMTtTu2bjx0bCYrYn6wnM3poF0xa0/53UnH7q/7Dx
iGROT0jTfJxwubKmkal/q0/4WeeHbPL1IqWFDXkvaL4SIqWV1ECDCGNChGWa0IacbFhLx8RoN9Og
fV3PIlY9qtYWkU9CLIZrV9ISmYROzxVeNksMNCOhesUjtf8WWgSAAdH5jnb46ERJ/96g7lFhWMX5
ZlrP5/W8kH9JGY1v0+qh0ClQodTpfncGVvZaWN9S7LXB7DehEppvzggaNnuJ6O1Xrj6j7tmvMxO7
5Okj7LbQK0KneEWLNllBK25RZ3ZC11YebTnhBiU/3NpFs+5JWaTX6wSI9tD+msLL+cTFKZnHoGJy
2wQO2wUKEBlpHExFDW4t0joiumtzE27+iORVTJKQw1BQ8TsDRTIPP/Ujh2YQLu7QdadnToltXvy2
aQFhLUunKs9XXmKBOm1llt+E4r5yGFtLatoEoNH86ZYv5/3jLC2jRKEFswOyvqmftbJDO7Chgept
il6aFhkzt0cbXEiRwdtrEa2Nwuye0wr5REhnSbgzKaWWfgC9RSmudfI6iP+23aemgoXBMDsAMATC
iEowUR/or0ZvIXc76f5H6kBOOHT+5eWGo+iL/D1u4x0AC+3OEXO1fxM7M2tZXy2dDWPA5YSxRZpF
b0r7hrzASQetxQ/eI2XVin2kI5DaLBPAPssmQttF8e0NvjlyCap12FRWUdHSvhlkp1ViAnpM6fsS
FyINinPdU+uOJkFZoiS0jd7HhX7/9Wl5PCsfNX/utGeMIVooPlmBj6Yg1de8uviw3zw4w6Kcr+Mv
OxM6NznxcWCdu7rP5eTXaKtNctJokBRaBHpMkxg4tJv3iFWqNqSUkIShv96p8s3I/k37hUnjeWAK
j8bVESeDN1vArHSSDgYXkD8iz0jqsyjMQJP/RZzXiMzVpr4xYBtXdlZGOfA2RC7pVnS4Ay59ZEEX
I9Nf+Y9c948+zYLJJH8oUM3bhdn0zTVOUHHBAdkGS9hp5ummAwNxS6v/dnpw4a9wx/38l2ADOlfl
O72MFq5pnn75H+zJWoJJJfojK4YvnHttq6FnoiP9uS6Mwt5r0FvJeKIdn9ohCP9/ifqKG8PgbsAa
DbLdgM69yA2fLaGDHRXJuZ5Yrl8PiwqzqlDLD9KC2be0IyWXwo9h0Or6Cw5nzMk9ATHhUFTmCra1
W0SrTEpgD715ut+5M0gbPkqxRqERfTK2JDiAuEGIjmwF/ZUBPK6F5Ut/OpUkp3nuQlvsLghxmZN6
fiia+zNOIUnOoZQnDiGp/ZUh3yYUH/W1DfEaYJHSvvKgA9xUj1bcYNfAEAwIdaVLkIIt2EmxJTin
gf8ycEln4GQ32mc4EqQgwuC0WYzlzN1+gxQzdB/roqCdMtzyBMEOHEvc6+TgI5K5VaHb+ln+VFjI
LVz+4oZPuGJYQJ+rMgOndtr3HTzWm+4CtCSJEVcnwMO2g5oTuOY3/Ys4IopjWYSdfT2iI5Y3+wCD
BR+gdKzMjhlTsBY/us4p55r5fO1s2xSIGjvaSEwZocAgXG9OgThBh9wo2sJg97VE/tqvGVnJUH38
B7ACuqYq13eRWbEcNesSU2cQ+Iq5DSy69SCUOKtFVOUYEE3Ij41LcoiK73SW+jf1BWn4lW1fASMQ
03gnvgATz/ELMtW22nUmz7aFUgtM/tGQNmo/V6daU+7rpD50eRHql83m49gq7qKNXfq/e/2MSU7U
e6iZeSDQVLX4a5x7l7RDinEHdcPa220fOsXlIJuKEycZv+ymlGTMiqL1xn47ouG6gF/IxflQwZhm
yL4qFhaCvx32vlQsK2AS1S5xRnemBy60qrP2JA1/suaHMI5H/Wyrpat/tdxH75IiYeeLh8NoK7Fl
VABkcz5Gd8RraMxs8djiX9Z09ShITjEsmyeaRaZnMnF5XZIuOckxvOBc2QKrAIGFe2Ch9Hc0Fbyf
NrY97tyPh6tb1kzTHBJkag4ghZIo6k6BFdKC/TScOK5+bvUzxm2qqObJE+sJHvtqWjSp2BoOlsUr
KO4YHPG+y90UJxbYSHFvRF4b39o/nqYnH6bPGsbyUz6YqTGSl8V2tJk68/6ykt93bY5dW/SVztwn
o22R2AMtCBa0JW8kyxhOlhnVgckeC3HvQH7JD0PJAXkwHP+dF1XOi13+ZEM5AGlM0Cgv+RLKKf83
F+/Mqd4o49jUihGOfF2IsWCgZlo12UpB8bRP1AAGgGqzbwJkHhYt/hnLlm0CXoYT6k8JaZ308Fra
uqSEzxVuId8D5BdmWTOGq9TMnZoyYomXNhVTnHVf5GzPLtteZ1/U3yn6fAXgTyB7QZHkw5QjSqNp
j7CaRvRIhLdWCmhGcr0aRqd7GwYZvjhBjVxo6VyO+kGpA1iEY5Yw8/ry6VWF72fjDuwBalRy+lA1
f0jWVbC2Hz/0Ykp1sWu7x/eHQeDcAhhVXip6b0KVBbQcG8PlbQjW4gGH00ctJE9Qjr0YDIrQcNsw
9hJY6rfvHHDMzhhL5P1wq2oh5ILwj7RvMDFzdavpf5KGIup+egi8w7ZEw4BPc0N7CreUSPWdD0Ue
Pr4Q6Ou5au/1ZPL7l6B4K2zKUDXc1fEH26JAfuHzA8rmyzlbOXMttzmWaK3uFUYAEkItPxAMTzRe
HC0Waqrto0UIfjhUZ5jq6gpykMsgS8V/+sC3PZKWTcPyKf8nHN8S/Blgp2gFEbbyTx+MbyQYSLbS
RyOLQJCbADXq5A48gS4OJRbU3lEUnzrqpRzZ/AnBr7zblEVBcFIL3cNgmRWEGPh/gwoVp2MskpmS
RACru+quCLS/yOiamkWbSIgwd+OX6gYxcfNPpTqRoLnq/bBX7kf385KBnEr8W4doxbxS1LP35MXi
kG1nU4rCqjb9jbZZdvXQuqipppA9i8RfJINMNEbE/SylHyA6nzjnTIZjbe/etiqws5JCyGPTb8vK
/R4gWJOT6HoB5kt7c863vx21K5Uo7GCfyZQWktmx5opXpv8rLLV+U0JSnUp6gjQCcBd8AbqmeJ/P
3TX+uWZ9rtdSvrPce1CXrBqOWc6cuOGsIqoXqQofdlbYjVe5eynnr7Xyk612acgKPDXwSSLzsxAG
Cz0GmoqjOsXke5pGNo4DTpoQ0/Evbojwq6HhiL7PqqArBJDQDV9Pm4dqDhOsrtbKXeZZL6+f4ONq
Gap1Ct7EmnvQtawI7ENx5qZmzyw+lJYAPjCuPwEwflm4a6NmM+zFfMvKtgKT2/C8Xg7eE0Z5CHK3
/v48fB0DSIF2Lkq6bBcSnq3xVlGgN1CDrlVaF4f9I7lAWP+k7Fm2qkCNDRE5RZ36Miy/8V30klKL
vNS7M1VfUZJ/e+TqxxgwnAYDWM6ylvwbx1e1AC+PqesRxaxTDhjyPglpf8myJo1SmI6Epu0eWb6Q
hwuwz9ERXTU1C2XuPyWToQ+GbKT+1tdyXf6CewO9u+Cc0I0/XvfDUhSnali9UpNt7QCos2pyXCbW
Dsgx/8vg1+dxbqZiNjLHsRbpS3T3tbstQpiHJPUJmpRnnEZ8uBRdn0hOefTTbI8DeR1rcnO5DnnI
HkH0LdvtVnDj6KILolRK8TvANIiT+cUDhgZlPzJ+3kN7ck+g4Zy8hyiC50vle1q026uLMcIbp2lT
sF0fDLZS9EBJdiljszoHhg8uHSM8GB1MGmIy8+NYq5UHlsZKJ/fvOAwEbDIZbUDQTL0dAeCDQxvF
+POUoHndALiGROMb16pN0eopbF0+HD7pnffqXmZH7kwulp2dyx5jkP2ulbu2zs1XF+b6Jt/VouS/
NAF5oSST1VisR0fL9NpEKvLlUfi1ARInhr/l4g+mNY5pIxFBxASMuf3bv3Bp7Rhj9i+uCAzEaVoa
C2NbwHMAET2N3ZSqhmFHvJ6Qo6gXxEl4XOyva+P6QU4zyc5WCjdapUeoi5ZkZmOz6dO0g4FOM5xr
mWKgNv2QuhB0Eo1aG/bfXIYExu7jyZXj5F3uFgLFpn6tQNoeatOcoshxymYeAvbG/tgJ+/0z7i9E
jdeXXq+Idbn58u+y4qXx8Gkke0rBAf/q6CXILCCkTM5kF2XVGTYwIANnNAKGbsdVn1T//5OZjOn6
WFx3mtQXEek98zknq4F6Ge4lr4sYgcEBFl/NQobksjiEGFG2f+lDbiZGAiloOPG5r0hWmOqPt/rF
0YVK8MPYf83ULksqIj62u9jWerk8qXumfLXnVZfOZQiwP/zmd5Hm9r2yeo6j5U+G2zNFB4nw+cSz
clX0bhHg4NtmJfkkzKV0/dJArxxLA+D0Z4/26TkmbgWpd/a4hfCWPkcwgz1C/EBeFWWM1WmVK7bZ
T0jc5xetFKoKLB6hMRtfL1reu6RuTK6W3WvnOcUTdSNf7cgroU9B8iaYFc9eOqwewXFmX5Kn8jc5
BdP67FCJZdS+kQlI7SgR07tkTU5YRuWgoPoSBTwm4BXdYSV/IMSb6HrqdXsXfxKX0BPHvwMNHOpq
XOTKg7KO/nJck2KclT/MS+DjIrVeCuVOtxdR+JvGNrASaMOtbS9Koyuo2wNlTctE0BZoKBKQ0pGG
OK1d6NpAU5kn1yJyucU8qOC/k651WhEbeuFS1WQYvsQF+xMXKnj4NwbYmEBbnHwNwM6UNT5C7i4G
Napklni6TcjbQ5p8UrsJQ5tzuyTf5wIehkmeChjmAehYRwJn/jH3SOEeOiQrcLoBAVX2+35FSZEo
Nkpn96vWQxWU6mtnjHo3R/uvvrmrIYezzPg9jngqWRCb8pISgC/vTEm/P53qrZwt+EXCiLa+zvZd
uv1LAjhyRFahWExckzEiCLFoDBwMSIUZ4ZoBx0MFhfGjTHzDsTZDfopWOax7U4q+Wlmq8vG8deu4
U6Y8R1YZo0EScu8FLR/8H/w1MgpK25ArdJ/3Dvtc4bWsUFTVDplGqpPAEwDrRyZeshjoBpZgb8cN
kGtFNPXtFf3S7P/Jhri0uqwJKlqX2z8RMLDnlqbP3S6PVOG/BLKyyOn4JIw7xgJSnmxen1YtKyNa
MtKdx0CWuGcg/lA8uwgBA6Uq1BlnDQUFa0VlTLTImFmdFPYTauPPYeYKAxYqOwkhl2cfwR6lo84n
eTcvE5Bmx4bqVsHjLmH+Vq+5x+nEhmkByArsV10Dv16DbhbzpHI3Cirb95szO++QUcMxncBQorcv
JxLApYdzi57bMjgPijDLuxyL+jtp6z/ereYJicQISiRSkK6SmP2Iwzb0ExUKEHb+Yv4/QjAQ10Ok
CuGezmmeaxb2fUku+29SiVHepSnrzryTJKkIhWHMvLBuJEngEYXqos9Qjgt1l1pX/2UwbpEpSbzi
np/vlCbtV5oTYWG1RSbH8t72ZsKzuE5/lKMQhrCDgHKe464EF+njsOegNemvF79tiVhYAHpg5iIp
ZpQeXeqTNnETMkw8hZ3itr6iTsz1Vsv2fIcQPcFPMRioxY3vr2APA0JEUk73s4sdOIxct1aXrW8m
VucBVrEuEuU7DtYQDD2qJ6Km9cmzGYef4u/yM2Nmoio5Mmb+GZzAhWmv8V9dlWy3F8UKHtU8y4Dd
bIcxFMEu6hqE7JGK+xbH22JnMrxNu+W22NlDphXWtoudGGvV27Mcd8q5OvMeLUo3igvjVxybAs6t
ygQW7dTindC/EVzmpN0PHKm41Z8hUmpZJfnkS6csFBHM6m7q6jjzjQW5RAWtViBduThCG0jBoYuc
8qclu/oulJbLtqyo4ZQXFqx/yhwtaJPvD+JievdNSb9ubijgUxdrh2hcEJnIeBXQ+pXB6EcfxSpc
te6zojOfLrcTFE0cBLfrM9RUOIznQSA+4QEX2y3EIBQQc0A1yOsGiwtAEzNeL0yzm0gGmFxZ16Sw
8hdbnc3ivJzYv7EdFvXvqSq+YYld5FN0Bz730ZWakurSExOLhfqZ40P26JzkDwqzVUrAp7hrdsN8
xbP4Hkp8gR+RYN4VyOR1pRge8uDzkC8e9zUD3Py/JFehjMdjdUNF7hii9GOhN9JuU1IvMj7f38X3
0oR9JZIxMHDyjcnZLrooUAHUF0UIIlv0KhbRTZ7+LNBgfiutZZ3N2ipnlT4m0+kghezViPU4LF14
iGkSrPgEEDaQ3aKU53UrJ/rqq5CS0uXqXfi/RKOG73RZGbQtphktdUy0lBEprsLcMPrtuQcq3kqI
equsKdVLio3RXTvBl67cVCizNyB5XxtEpjTLyPVVH4C9baD5//s4H8+VWgxOpRuMagENphSoMsc7
Ff4yFQ1X1prsGPyJk65nUECnRqnv//MtT0yXFFJNCtqwwH84IchzQVcZgvvmcy9SwiXS6pqvd0fv
qI7hBjvs5InXAl35PdecSmy1JyWDoGXkA9P4UnPeyxGN77oHVW6nQvrJYqS3bymepGMyeNvIkF1j
uM1URE90fGzS0+W0K844NRfqcCAjuIo7Sq5BFVpEMzsE3uT8EEe1Mhqu4oqKiCzaUldBs6m0AEbK
MM/WpAQllLQUOSDp1BJUVwe0RGVaDo+Ch9TNhmKqSaMXv2Sh6blPuYUrSXcFMsWUc3t8/oN+vXL2
V0fajVxUQKHf+skQH0Ph+NWiu//FWR4a50b2EIa6NE/n2sB2eakepXYO/HaSKTgZUff/rJeeEZzl
6S/d/HKBgRLng7Z2glvNmrcZ3j+awr3Nkwi1iB3kq1ou+fN2g2T9guUfJJEhBojcyb7pfevkxIxi
Wjoic/y579lbPp8qw/OC662L4TOOkRl/XYEonWsM8Rt0wRK6cCzTwqRro7En5xAfOTEE1hR3A6iE
arjq2+sRZiv7FKYeWK5TjgNnGG8+33FSURmmg31CQv6dJup9KXgSy/vlW5ipjityJCKD/lvgicLn
MWQriZi9yTNWak/1idrAwtTApf6CFGgkfMeZpKpIS/6c25BlCvJOC+XHQ67vxOTWjQJ2s3Rv3mCL
20G6FDr8prjmvPkETknoI2fGkyrgE4kwXqlLQWFc3ok3Ew4m2R9Rr/VEGudouKlULhLbSN+TIH5j
aHanvncwItRHI9C9tDjzDadqH3RiqlxZ99uKrsTeuWNlwYc+qfucnM814xZVN3x/iydVqi77BDEO
cbwIFYtMv8JAqn6drRa7D+FYgwt2fpxFrESZR1UbzMf7r7/T+jJSi3LJ9uanAjhmaFblJm+zf9Qr
Qi3vCCPBpQYiwBTMKs1onTCsYEGseAaFlHTxanPAwRoWm/CdFcmxKD8cCet+vNw6/Yxod4MtZ5sf
5S4Zbr44cI2AADpiywafBc++iuSY+I0HZhMI0xZ3zpzyqiBLkCK+pjrbUJY8xRL+cW2QFn4cZhuX
Xp9jIsaQ2LZffthox4puhm2qF9mMmGmgldPoFkzdnI6M1ytl/UmUVBS4yBL4WJNfGjX7ZvdfVzjU
+4v9+CCZb86v6kBELWdgypidsB5k27YuWHEnExs8+GQ/oaf5LasJ0WDF+qvgMbwCBwsVQRzzCO93
um1Tnrfk0chCi5TTRMc2EnbLPw+DUlbK+eidP8X1rgYKIXEo5QymcjMD4zma32q7zY2oCe+MP1v6
OEk2WenUY1j96adIDnTmLGY2VHTvDtW0LUxXSzdeMi7dGhHklyvGGvrwWubfVMEdp36uYKT+iTut
bfmSyCTbncdp84jMvxVbnSvWGGHNK+7yB4M2sjOwK8LshM5HVjUXqDKn51wKLEZlAD5Cpwyqzt+1
87aYhp2FkL/HWNo8XjUfW+aet9OmtJwGI/Ian1VsloJJHJwDdzamYVgHWHpWNz827G6CDJoA7jhB
AAtSKVy7p7ahCUKRdlIBiM8m+hNSAQD8hrRj3RD8lYQtThAJ+e/sW3Y8L26ewPI/+Yn6Jf89YoS6
yARlfJSqUMl9MlsrZBL7INYS8TtdOhCLMmpQdoDe85I7F/vP6nlhoQZNasc1oYB+nduqPr9eAvvm
LZkKLhYFNgTSvFMs1j0Jkn3+z1+QoTFZn+rioZFj2BqbzYG39F3Pxe+uLDPbsi/5RigQGVLH7S1n
fWUskX24HBMhFx11Odcs2nk7rE4jibfkH5rSFtoeqGe30j2XhdT/n18dXJvuQ+vzwaggGvjYQrtP
AwG7Bjy0/OzfwiCzUsYIRI7GDBw7139nS0Bn+YwK7pcRSmiWNt5/pkMwN/ro3+xepPHH4waENndB
2pw8xcmxQjNJlxDye7IXGI9woeNanfKgRcRrZ7EPIt21/I7yCQvmOziOOY2mc77Ng0oYeTLXYG+m
GsdRIixW/aKX6yEwB9NLvqxEBPEQCCxIKfL2jjHIN1hIIuU+GuTj4TPahz3vg8fJJxzDznDT8RGH
eBWUApjIZwaU885wf7ODTbpMbQmY+72EwtzqKqZMlQxzbtTM1ughFLT3DUhzdjYuCOSS6nL4eQ3g
s1limNmF3Rxn41ap/MTJyrJ6Zge4KQZAozvata8MzZZDNxDd8r2i0U7zxY94kitdekxf341rTe0e
KrOJbyU0rf/ptInA10XtpDKBJxcBp+or0Df2bB+MR7ghtmi0Q6i0YC/GoC+n89e1xFsszqu0K7qG
3VA7AXTS5JqiESVNprlxItmE75a15yz+w2ZvEtmA0BLXZlk2DvIGh+khhUVZ1nELs45dRIP2F1rG
pvMyplRfFx8zGhGkELqgrD71BJC6ie1ASt5CQun2qC8EGieaA/QBW53UwoPqLsEvGmh9fNEErwT0
MRDvqXhg8QWSM3GJHTrl5L5dvFkcKmbImb2vt6u3wtx83lGqgqhxjzpNrpIDf+ETnKPazx7bmuWf
wMmT+ysT03kG+LNnvEcWKjkSYlpm4cRPtg4Cjt1i3wf4J1+RtSb+lpVfMAb9iLr/DUwYicrV/+Vl
cdxE2o3zd55hLJdnXckV2NNaZezSgT2csDBycxIkKIOsPexJc0elHjg7doIaJ0KAgp1CKH3SLVeA
h1teC2v0MouDby54Mga3a8QuLPpNlcYx6CQjxU2KEEJfKW8PSAlxEHLvcv49pemLHdtd/S2wofZh
J7Jx0RQFqWLZMxHVNtF1nhhYu2ysuySVFzi1Ppa2MUKregBqxwl5yWbN7GqDV3Git5qvnPZ99Jnr
MNWptcmXzciqs1lB1LENL+PmxDaz9fAJkFKAwd99cDP73tOV2Lodxow42OtLgcKXNJgiHcuXU8Ls
rn7tQ+WToVYjxIZPre0k5dhsJ5H45Op7AeccN3pFcFYPI9z0GKR8rwGEy0s/qWXhRgSswYXYiywY
6bRWnOegyv/FU2H1jUofeeV9A9UxzyXSxCdz/eYa0yVffZubux96cMooT+4w5UIpuyHPitTswMIb
6LXSI1un7VvHDwRsMksHU8f60fLr1/51dzX8l5z0kbSGFIZJHz8Dl7DxJgEV2IU7HWuHMewiyTxA
o58+T30pdUAfO+onkWhp1QS+5aK9N+U+hY6SUHZK64U1A1oJG/Z6g5YQdZkQWNWD7W7oHoptKsUS
hRW5ctotN9VEGLbuCIhcsGQMej1JnuBuBu49D0m7VQySyiACxnCa8eZKNN+QgqdM7SzjYWJ+0CGn
ya+koJOY9MXYu79o3ODjMovVEd80AgC9mhSRpq5qzRipIpxBNE4o+XBxau8d0xfR+ap785bigLcu
up4wNxsdwOJrSWONIDXVJMtUhupDDmeQcqrcX5rx5VpTVT6WhNuGkRyJs/lz60LuInhWBnA8bdm8
XGX6MyPDaokfeFZ4t126ru5ePF1LReEPhlU1nkGqrORNTIP8U/nytOSrQC+4Mlm7J8+q3QC6rbEs
TNI+XXZ26GGLEF9Cm0488z4Irwo0u31oakBJJPyEKBkjwykY0bi+PBrZma8hEBSaQFUICpu31geC
3siYO+B9nko108CaFptmHtj664M2T6rdq9vdkdZcXclBXwZSmNUeeW4NnMtyniDZXByrbDKQuJ4W
Ri8yKHt7nfjz8F0HjIQI+UNiFZ9bH2YY4l3MIYdMOW1yX3kxwFfAjlG7IV5zKLl7+/OYww8PWkxy
5e9PDHoVaHVFKTASZ2yBagiVyMzprfoFFdEDVE3JwaV4R4TcBdjWqxFo2czlbBl6/rAS5CmtFn9q
iqlA5G7W4LLFxxPRbhvfZ0C6C6Ir3SisNDrJzyWjURghm6OB1SfuAn5YNn0qMhesWl2r/AeLP9/w
u9DcO985EtOs0ju46f1f/gseXg6MqaZg+VvsmhqFfSOIKw/4WkKCCsazQDA9By3h8fgIhzfXjAt1
nAjDCkI66/ucA+//Vpmv1u0LlH03rKODHM4+glz1+9Xixyp/wIkSDqRmiScuu8wzcKYX6bRjXjr2
7+16+q+9cDq+lhdJbG8Y6TW6cfIqAK7wywUsERGYqvhcZVwAxQV3d9biXI+uKO4i/c4vJDjW7lfU
rmUVnCJBKUUppNBXhOF8aZ69VlKNVondR54k6IgRKcO6WWW+5k98tjaPczmDk7qUIktKMXbtv/YP
nbP3K7XsK6bWwfPkYfvaRl1kjMgPzSHU8jn8fj+u14cE/62PuNITTOfGPejzHKFTjAnI1oIkC3y8
7jTYKiBjel++RsspjwNE8yFHum6sLh8t9wU0imgQko0jbEhf51x165fXrZdCowkEZEpsmCouEVfl
lEbiW48EOsu7u/NF6tiyM1mcKB0oKtCk102UxveCeXbvw5h/dJhPLJyQwRRKoRG6W3Dly39/BYBu
YcvKegT7j4o3HlHgvm+vhAqFv8aCeNWSXsaAB77pM9/9v2yXbaPTt6dmoXOrOVtUNnKKDtlb8buO
Nudpd9YFpe+1QVCxlyaaY8VLPY1fgO07aHiz+rOYQzDVmPpiQHqT6xJiX2Xm/dsDi402y/e2itPa
FKz+kmApCEPGp1WaExAyEamwWFbEHTiiBcEHtpFO4PQaqXf7wnQy0b5nW7xTAz2g4ZjmUeYIxxxj
IcHRusI++Wh9GdZjlSzLHEbk2ezP+U3PL33uTTz2wlUrOB7g8MtDlPYYw2PH5qHyLaEYl3ra4l7u
IkOGLNzhMEXedUw48o6Ila0PI9e762Nt79q4y3ab01t7V8yfUtU5Gcgl16mZt2y2bniQbEK0QpIk
8n/DfErE8ToSs7k3JXElCKhVx1uTBMs/OvxeEUXAxAxRp7wl4uNmAtv7gjk3cFA3EOk3VewUYnGr
XcwyjqJF7/OgJRe9JhRAH0GebXZ4qspDprp/75SZEyr4UUch2NGy/GjmKAHf2l31QL6O2OksyWN5
v4AQ1apXkq8Ao6YiaFLAQ+BvT5Ir86Hj5HVmt/frgbgotzPXsSMOqWuVa+wFgVEkymkqKM5VuJLv
boPHOoFO6zSoXkZkphRbtkA6WsecDiGBXd6FyNh+O5DyK4+xV+TR1W6lcR3USImX04VIZtrV4f5N
8z0GgL+QfHbF2t1Xo9Uq9V3uyGvExz+N2QbQStW9PHZ06ldhrpLwopWl84dx8TYoiEiDFidyLjks
tL0bai1l0ocrGyLB/BY259Nb5ZHTl3ussN+SzehX1lUrSW9ra+ST/UMtr58MPI1GjYq2OgfoVfb4
31C2dK9E3iW2y4qw8TA+k2kNzt8f+48UCSwJfEO5+Kwpo1QaRIpkFV71zjzgvhAepe8LGYEexjwr
VM1tdoB87tJ03AEVQaFN7/qi5ArvoFiWjxVzUb2qwslw10hODTI48J4uYGNbxHRi8kbjBdcUjrE+
dobrV3l5UhLG+K7TT3bpdSFdTb9V/+qr4gn7O8te4KLdUaMwqrobo3TaU+wbl8I72mcPm7+x6L2F
vc0e3EOIYNhYm4CLodQvj5PD+P9TpuwN3EXQxN2dMT3FIvtZmvrqsA+XJ9X8s9ns2bQYEcSnVBjt
KaijCjnMnZu6eJ+8nvhXzjOLNYGPGIQz/CLcwRb5UKL3/NZFA3DlxMXJ4cFSosDVVpwKMec8r9m3
oeuTcZc05ZmXDPtMCADwYRxC8GqUcGbL+GEcwYgGfFdNXdheYdDUmf9LEaqIqb4nIqdefdwrDfjW
tgsKdz6wQH9vE8oU+sfzRHRMbO/cqsQ9+XMiSJPmF7kS0icopYse7SAclLGkOz3OZCp9+9tLKVH4
2QGttqmTfwaU5SMXNyyO7uhfAKpzAZv5kPP4MZFjYtVdoHVWw4BQQvroI9Djn4AbFqhjZ9jHE8Yy
IDRF445dytUb+D+pKy2IdBhTLF2YZTR6SzryWmipfZydbihMDR2mRVkaDJ6bCbs28lVzOa7pqAXJ
ylwV6InoEoA8SfopWtrOfdTDhYi5TdgJOjTfzHp1NbiyTCw/BRCLZH6Q415bfgdRJAxqrvV5X8TP
AFl2wbneelT5d0Vbwx6Noopc8TKc8y6g/hNdlxUYRIMCJxOH5pOlhuPtVG4YF2+TSMfPQzQKbQdR
IMVKk+0v9edENRBrFATg67AQE80r5n45NBaa4y7kniEzvTRzUEJ2OiH0Je7Pv9uBiFwdN4wLMLD7
raDki/cFZWKS3S0v+9Js+TRXJ8KeNhDhCZLKJGeEbq6jXKgkWQGGIS4f1pRjfRFIYCmdHIWwit64
sB7WYd0UfX1XiI2+qkpjBmpEkmAbPdBm/ZL7WdJSZ5fyrvb09YfExnxXOVm8D4+pN8b31m3otIci
ZFh2gCHRrC+5joLg86cqMXQ++aLQo3vakLqpMZWMzf2NYTnQbjL9fXYYBHfnUM90WUL7NB2ZKyJw
i2EFqWGZT6OTh7G3wA16uqL/+tInGmtgK8BgfUorNh3cX7EMyU09cQgPAda/meAIWp2CKXhGTcRg
tKcYvEloThAEB6983eXi7urebA3FgdgkHXmWQxWLBrG+qmL6OTV76RBJEqt/k+DqzY0QiZrXzDNj
pGtsdXeQgf/60krOuc4lq4y+LY8/69icucSnfnudnNvPSSHcbpqoA+5lnnxtqEQBl0//lY34Vg6n
hLCP9oDZthu08++NYfJCLPGold9/Pp/WcBl0Ohth8OJB7RVxGy8SuxDxTb7SDSywvgO09jwaSAT+
sR286hFt2Jrxn0N0V0RHaOU9cy+biPM5lUGgrScbZV+6FUidEYGWpNNHmlnJk3rxXE1EcU2VtVN0
+QGGnZmNCY6E4pPq3Xn+/pPkBuZvd0pEqwMqt/T6cb/sn7ZGwOCywm1gYSU+TZf8yavoYNfreoSz
vmCpE9lGkLsg02UkcpTHynW0DEleop1v5EbE/7QnUkMZoZc7HJB/rpTa7UFdmSCSFcLSIrO29pwI
WSvMjsoIWESR0PwvRCHrzaAMlCR9utfBU9TEN60p+7G6/+98GkP+MjBMNxHm3uFbNCmHA9jC87UL
w6JeGh+q7jo22WsECFYH96tgmyBaoH5GgTa8z7XRTF+LKbFNySbi9W9lAz1J0OJQ3b0Fhp41A5ye
atvuXyIfSQHl32gzi7zvNfMK1Te2FjI4x3bfUIx5pYvWVDfGzPQNN9EnNZyqqugCIaYxQSdnKtUY
Fqc8VsS1L94x8fr0JR7defSRCYmkqutZKCe+/FzeKWRTCoph5/l5oJ4yjeBxEYDBcekN5Lwkqlgw
zvAtce47NEJCPC0yDyz5Ajp5qubvE2oR2Bzc1kP9y7KPVHIgwuI+Ogb/BVKL5qqbha+S1TUpWmfE
0a799WYVNi5r/UI9jv5QZuXrrFSk4A/q05xAqRvg79yMLhwttDzh/ET9/lQcDoulUX/zIVfYYQgk
ugLC0foYUwUi8zjFyckk2N+wmye+auqJ+yW0XY5qX7Av97IdQX2lu8JbxPti6DT7vH/fLgPu2MzD
yn26EltDNjLAy38vx0RGJ7cLUQS3iIy2+F/25UJ8IFRUR2lx6jPrOWVezrpL90sIgTaYWfcdSvYP
NiyTcKeRDivqeRgw2RKv2VnIsF5+qTDiwjzZD1YSEc0axvhWRkGP6Mz8yn2HZJD/uVBZRSBdKUPb
3Onc7u0rhQlvmpkYgyj7RWI5C1JJ4V1CFbnSIJ9J0LprPg7ORDqfWg22co3J9BUdR0XjmGYmh8pJ
y/QZb7OMkXIQ6AlxNV2lXR9WBso6kbURuzP0jYusFjmpezuYYZnXfonZhFDGMqNKS0+ul4Fvjb+k
HW5iEDOVkpzB9mJnl81xHsH8+wCLvRnMrGAGWEeIjG5eK4bmaF6gn2d8hud5K8TEX8tsxjDND7iP
twdTut1O8FGBVMnDbc0DtuS2ZiCaJzhquRh0qhHWY5KudKH85XNIdHddQVsDf8S4y8lB53r4u9sm
T1sxXN1PbSjFiYI7e74pC8AMO7tTVYtILeqEMIpqZRlM6SEkGmD2/Z06EiMbNJw2uvlgCJFUQlmu
DygFLqwR9yKuUdemUxTCuvnlPO6gBOw8eYrq3vpl+YLesHr8kQE0F4KdxWm7V94R/8FaJGr1XyN2
tpEJ+QgJm7dIyivrq2F28hwZ1fuynVNPm4O6cxhtppSGHlfV1Y1Zq2yfslAkw9VrEYN0KVL60Vss
3o6MBN7qThbpOKiD5mG5RFVU247L/eofoZSIuOo10mGtfz1H+fYc8tUU+A2cHnp+l/aVS0LUvp9y
CodPsybbhi1RimaD75Jr1aXnOjWl80GRM6h3PhJlZLG3UCt1sjbD80G88oWYxwuehhsfLt8wxdW1
kUEkGV1o+BQvsJyaKRa2yOYmQf+wELi5GgnSzjE3/OIdAbhahIMMXcU1xsMRMDsQsSvNqtgaLQyw
Flh8++8bSBTuNeik4dfWQxdrNrPgpxizThi5DhBVw5wQf52MLIPfDQRZlz20tDDeIDSYx9nvsbMe
ibV1OlHD89CZoxx0sJ0gFDuWKijO6YDyHsjt7WRdhTlkvn4SZHdZ6JXHs8qDQQD8og9FG0yWENBk
fIcP7Rr+eaxiHuNsrNXVFhwqDAb+ivrDro4JkutZDaT1cGGzSSLnIbgYOCjvqVDLuPOyQmkeHJ9z
4SnT43cw3bAj+5Jy6fgLRPFJ0MtYU00gTnwtORF9gEKvl1g1QhJ8d9YDb8SeAIMMkzxPAywUF819
wztR6vNHAxe6AJ96+ja3pPFaMXUKVSDazWSRcQ3+pwP6oPfuRgs0dGvmFfnYa69D/XZBpZPpi0NS
Ttz6mZleVbA+Fyv9Rsas6qhMp8JZBEv2Wt7p6mFN1iGTFtK8UTRB5J0EEmhoybQJ04W/AueePTJd
b3o9psBGwrNHvHXDjSPYKkc0YrKGxMVsVqaXR3KA1hXRxGAX4vUu2yhkTzdWufOqdETXjMSO0RX7
7t/l3kwS0F+GGf0Mgic4pGTUQVjGajsdZDhtcbxjRG55eH+8Xpz/wjnSeODcbAAHCUB5N59oG/10
vv1TEJTkj91jMK5HNAO5YIFyAtkBxSJeaAt3Er11xNUkHaAjgrkXBWVSZo3l+TDGOM3uz7w/LqQM
jh/ygsFVvG+v2kKFtDa8iQ2tZ5wIYMd/ilS80otXEwwwZ7FyroNUpJKiD04ENI0g+y00u46VuFrG
3q3cOGHzCjIYA9EZaZLCICP8G0MOcO2Cr7oe+g9A+4IBSgUll0jYXwAygTm4AQGM9KZvdJORCa9D
ypDkBMa6VwT+QoveM+TkRvGuLOWLol3pzuLBLYwc2LNx9Cc8yHji+Oxr2XpM+Q5pLwfmNrMC6urS
LcJ2hrSmXQNyrLsYbQPNy9n7w0wb467Ey7B7mOAXW+4ueOBmpqhtsJn98cFoMjNh6ywR0RmZbn+d
j/eYA90jycgI2EC/9JMPUr6rSr2+3ArbKDHR14mkIIqOTi95Q4Qpv4+KSBNMur7D61B8vcPU+iB3
uNGXJYPFLRdJUR1OfEF0/O6iUvN2ZhVI/7zhyZ5FTb11Ql6dbh4bXM2ltMqaMaAj+agvvRqS+ka9
Pxv5rTY89qNY2Q9kW4KpuahyAkBrkfEC96JVvlVF2hjtCxyrhSEgpwTagfUICi1AN0wXcBlukEk5
rjCUTkZF7f1jVbwZdPeNMJwgSBd7vxD0JAzpIJcOmknCLGwktGfi/NGQgl8qfVzn62XDK/KV8GnQ
CBqa8dRoWlcGdXfMd3rl+BAJS8zdSjrV54ptSfZ/P9f7je6hIvGGB/v+/i6jyYxiZS4FDPV4uuMF
T5EnfNysfr/XQLJJMWDjtU3cwk1V8eKZ3gPPbtWaqJL7qjz+LnRNViRkF7giJT/iWwiZGrV9gcpj
AzlI7cZJ6d4B/AiQwwEvWdn0L5h0zRueuzOMZRvjoa6datTUUnrUdaeM1vsAKX2xrj7wrbcJdYRl
EeAm/n9Os5BM9INV3LP3aW3bA957kpTX7Boju4xQUSlAjwLAQWBNZLtyFdIqRmC0921S5kxMfBPp
5TGsDV0+j00Cc2c2Zp71fTQnfqG5GagEoCg6Rmv0+cnkTuqKbBPonnihPeP6vzbACNsIY7Kfhnkr
P6SWuyoXlxAyvqyXUjXYOw5ZfGD7I7Nt5FeWY4+UwDXSk7lCZmnKXi8nmpBxoqvP78EtpL/5HC5j
hFOyyjoZh60FDaGOCtxXkfIKYBJcB5b1gVW/VgBymWdjGthuKY8m9EdCSqEQ3MR51XEhYx5j+eTO
duTPDnEhZY7ItWw3ItTz0mLJN28A+7m4WkEQEZJT0qzoQa2UW8QR0JCHt4t1dqshp7NnjBwdTdCj
1noiBHYFXm/i4rJf43Nq7vEf8iFFZ5mpcftgOog85odm+K754NoOEYwYPlufDHdxMJdNjAbn8DnM
3e+frepGNvLm/du+OcKo8NBcdCXEHR5YWzHRAU+D96sbdoPLGVhBCWr2IUAvbfzvoCsO2JbHKAzB
XnR+4gGBeCJT3bE+9LtlboNZFtlmvRj8D3xBeB/YJojHz0efFmrHPAyBCsHIhZl9qEAXLZrYMd5M
xfdtQvUT4MditIXB/ItjD4Ccx0tk8pQwXSGxFs0e/uXl1n5rUJLeEgX5qDQmEVmXFr9vbFcFwPGP
Jk4VIPiD7yRhPyqUVvsgQZ2bHys/HrZrFjBKL+UUL1W/wQUANYO8B0gPBb35r/tsJyFL2M9suuNu
VnsKXMhRSbsrWzpUQhyCJ/yVGaiHF2pceTK0vN7sG8jkf+geM6OAjHKbn5wI/83o7AqbRmeA3kmX
cB6fwf3Wa/6vUUxdbQ+u9kjnDNOjAUXMfjhavUiXnyGn/eujg8oSnAz5Ukc61CPE+tx9ipnyPKRm
24vwTxpW5wgPMt3WfoBJazzECwFl9DjQZMuEaAAXZFPvCoHz8l8m0mNW34/x3fJebutUhpiogNlP
g8DLmF1aqFr0YtQYzedVsuHdCQBplmZwVniNHqWh9UzHm5fFgbk9TRbzIg6a+EJ0ES5ufT6dbvt9
BRLEfRwVDbNLxYXekm8t8xe58Y2M2uVqcyaIN9GcA98IFSNzIEBcRRjAha5JWXR4EyyKSqFHVDOI
AP9Rka7Pf3vUqXuzsPzXEhyAo+Vo+zVmL4XjmyWvefF/GYpAGebzfAlwbr6kWlWfX2emZkJmbsi+
oQUxFmjsdxjsq/uUWvN40eKeSyV6RbJW5BQ3Rxae3FXVvf/aNpwZkmGptEw118jH5JaMzPDHgt7D
in620T/hh791Xpuovol9tzz5n4TEAhZrh4/VtGX5zNquddbSFe3S/zCeon8IKmrtM3+6toigIAAN
oYEEOPH29tlPMCrCntbHbkdv5+C7airc36aex0j6Tdfck1k8K4wBxh+9NswFiUt3Y3pkXXQs4FH7
kZnx8bPXLTE8GBFp5+d030rU7AbrffK51p2zlDdltSrB88oVks/ZwjualwLEfmDM4xv3IE6caPQD
ZjLm0TbXpGpwQWgVcc3p9ggDq8mmhCxksGVF5HDyoadw6sMLFqqlWY8BboQg9LtHD+v2XWRUXKXD
cXvKilHaY/3KsvjK8p399+yUBCm4y3ui07ehkwNHAGUOHFxd++iJz8nalOg42lyQ5Gv7PdhVFrzA
UfYUpQ++7xV27T/sYMUEOvjuThLF6GhY6t1WEo09y8vOsm8QBtE9MbazhtP7AwJiZYJUDLTcPh22
hcPU1LgC0uq1fimk6mLbA7Bcrn92Sds677Jp7QOKOSzabpOf20Pg+ul6W3LhiIuDy4Vba0GCluk9
ZGTVEEc9HYEtu25Qh1UXQeMnYQZN3S3l84VuSsCZ7XoCH0H036AWKfcFYxSVUnS2V1CPdNUD594z
+c5Yo9oNOpXI8JCpx/3XpFTb0O+edazrAKQobPTl+LwHmSqI/l9/IF9/6Lbk94tDEs84UkdKEXvn
LYotdYo53swUdhlcdKH4JUGt0T2nCI7J0gwyxdLbkl8wjZ/jmOR/LpbVNod392grVNarMPpFGcSb
Y2cxIc9J+q+f5bzLihBGjsJ/Z1tzcAg/VqfgZYx1ApNHs+NEYxc/paTnuwJk7GZf4lB/x45kloVV
JMrt6q6fhxqp6OwghSI6Vrn2YaCkixxEExZfE9fH4Ybtxr8dekrMj5xfcUHLAu/8OrnAHedzMsWD
yKezn0Gnnbc/Sy2cm1rTaVeFDNWjqEAztLc3FAmnvbfNFLZZCK4pQ0MTuXvbhqoJkQfOSvFbi4Xx
5EJpXXFr/T2olSUyKrKxlsbT6jgSmt82JwOFK1iD0mzWkuMzfHsqQH1OZgsby+vHWr9b3t5Yt1IO
9L8SS+O8iBQrnOWE/Ulw6U5yHIDyqSSobhXCRsVjXGOIq4adHc0r2jEsFBg3SqizVDhujVa/iwAS
zzWa3DMU2toEZm6s2PTNQ0goAe3PIzkLToWZkfP2nbpyXz5P8V/tHV7BMxC1zeKrJVVXfCY5Z5bM
bRQypF6U0gGxrlRX63wQcBll3kfvZ8Lfpsh4p6jVAZmF54pWnBDrpEmz4cFCzORngJTxxzh6Quf5
aBvh59lDHm6MaxBlwYSwJBSBZLBgadhxlikxcpCZyISrCv79zUy+AIGHdu7w4VflU5iAB+5NxE+p
QwiJMq0ESZ4AMpklWM8xccpWDBGKsEza2ytHIenEIWexNSPp89vSwdYk+9/pb5C4ZZdc4eZJNuxW
1XmdSgOi6fsowPNBDBQxMflyGgkfLx4FjQMcmy1+CsVvKehXg5qHxM2VWsQnp7q0T4iPd870uQ9S
w51zfgXVMy+tMzdWn6p9hqUxZHBR3mgknSBHUq0iK+mjYJOa8oLZ1d4uoVFXwDBHS9ECRLRtCqXh
U0ec37yhjqH5JEZQpePwf4vrnRHOfYn/ErpvoV7DU3W0QVMLqnYObZZ8qJzxFOR2EvqjFUrc1ogD
Qby1qUCT3PkddyxBYr7TIoclzhCNnR+WuCOrY6rLulTCdZOYcjLF3mavbr7Sijz/Qo2cP/8AiOXy
WcufPq991NkeZAY34krOIIWC93BirlGHgzg4Xgxm/28SJTTtcZ5xgWDkCpuyhS90YVWnIRf+DBgf
uGnPQAEw097VCk23kj+co4zAZrNWsH4iD0P46HHamynu+PVCyCC5pgekJrOimvbo8hNEiph3uxxb
OXGCk9JZHEqRQWlGpLhSQk+sQ/ySvwmDoW64t9uZ6rNTV+6CDw38W8MrtYsYqvww6L0YV/1PL8EJ
kOnveYaqgvNabP4k/mut9bOblvHJRWvHuOdNVRkIPXE7y5MhXh8i8cH+KB1Ep2YGUXILm4tXkGLn
Gq4JVYpwjESzRYBav+T2qzFX+SzrcJwzVFYCToyOW4KK08PuzIu1uh4j0TaAAVBx/BKqQDdtNzyG
1Q6Z8UKJJTxNKi9kvCLxwKOVNF37zfDHQVx31+sZX6alRZ1U0uHPmUNdpSozPcJAar32kKn5APkI
6ulm0TNusmlU1KeXhbIXfq4an3u57MUb+v8AiJqHjcMJkWc6YrB97Cz11bJUlZ7KjCNwXh0mMSxv
GChoVhSz31fOn6TiraxUONMtmc9z/YSrZYSYNzy1J3UYsoCfeT+2/IChajrEP5li9OgGkJC480Rd
QV1KpiwBMs92nLBo3EYW9f+pp670aqbUdvvn/AymYtg+GUrZUdvlab8HhTqFcQhEKbWyCzU/l3U0
PteTeat07VamAC6q5yLih3OgIOUMGcq00APxkF6gIuOrnm3CQRkw3xpzcOu1p1EbWLKFMv0t+Ren
TB8fqwv6Dp2PrMOaSnt/Pho5naiKEgdaWB5y2O0uBOMKDRTn1Dgl6FkDDST/L95QOzQm1whmogLL
p6ETnupHLikhCbasYdmRWYFZJU/TYInlKtqWmFocLeRJZk99BYvKCeewe9yTKk1TKPt9LADeESQX
PiNLr1nrVdGKDhsY+PPBQw+kJWZJ9pW26UwlBzvfq1ZdkAnEyboNSM9iNch14RTSB41WWiqy2nNA
FzzVaXHLSIchHCIAPjIol7gGLzmae4AwUPEroSdgr59b0nUpgkdaaAAFqjljZJ+6ciRmjRShEzxE
GYgFI7M1G69fLgJdu1vyQD4QZgn5u/xeszUeTihQWCI3GGiviSQIvJp3im6kRHq+fLrXw17m5Yr4
ncYHWYWTIUSRAfw74o2qRIvuNBVrd53x5U4B3BtUxrWuqSVsHr3DlCkxfEu+1f3Eljoxl1Wbvg8M
shBVhIabqa5ta4jPXr0Ll/Q/z4ILlY45W1LdD3FGsX53THAkbiSIxcb3BLhtJFD86H5maA3CtWX/
CfdkfsTzD645qVGSFej20G4ZiveewoYNO/8jM49r8qQtsdlr7CK8tUze1GocK41tNAQ+F/Hivb+Y
bQa67BPDlZrH/RRcjUgDCD/lfs6ZIA3NwKsqKpwXRwRSSTVpcal7gyMsP7qqLE0nnChSD12Z3e7G
kVIntt1qEVtW1e6jEERhVlv3ePnSLIodFtjwJlcZtX5dr53Zm//iz5lCRuhLfRpjV+iX54slr0kw
57HS8NWV3VBeWX7jtY2giZN12xIZWZIHkyrMeP+ogmfjglLxtYVza1mSTpV5FyMdICqpjGjFysaS
jeZzxE7qG5cH3FCkauC6ng3Kz2+kAFJqmFUSChXeqQrrwviguHpBBOTBZAy/7tSuGWnYVbZKzHJR
tguY52ZmaMgBRNa9qkd65rZbSTRIZkwSEx9bTdTyrX81jyy+aimZWrxXkbbxajtL6TH0lE6iSji4
ZEFi93ev5kvsXG6GmCYtfHWhh5Z2GXEwcYU3DEz4xy0nlNAH+UAY0KinbMY5+xgXoR8UP0H2LmzO
Ef8C3zGLX11SmhXWytkPRh7mu8t6n+8Rr0DPp8Ku9S5ckNy0PXGhHdnzXWrvpb0pMTnX/oOWrmAy
xgMNLXoC4pDAgSwtmXlN4M3Idq8Erm6yFnvj3+t7MTv5wc2Ho66TE7u25ArqPX0Oq+vrhdC0QCCz
9PEEAOweuX55lDhrFEZq3U+MMiXvpSdgmhaowFwEtlQjG1yuPgAJGGckhLIWOmR4iPQCoexk8aDf
NgXjCWEySz1k8rJOWlrDuLY9fX+9DiJHNyt1L0jf5neXDxTE5f1yt1J5sQRwLliL4+jHKDlYn7i4
dCDoWgTbDA+f81nJ6rj/u974jU1hEoh4XBnq37TryOs7nt0FxsE26On8hwGJeaurT776ov/UHmTR
GvzR7MA2h4TasWTqRQasJz3ERbnGId9R33ZAmD5ooiVJ/UTGngyRbZ/2Hl6Y+uT30R4T3qTyK2gx
af85qB4qF5PuIwWk4KwcYxSGEN6OPmoiMs2k6yOuK4ca2aWC59s1Dx3o/xsbXLDGDh+mwDWhVj9z
Rdonn+TMgluPxDP+DWhhMp4dmnuQfstHtT+ucZGUhqVQ4bnrZlWSHyszlsK0G4TBH2okU7NmHkME
hpx64c1BDNCXhVJbKLWrpRFmnSowVSvQCog/I1vivZsdPRTIlWiYEr0xctrS6ReSmi9bYY/SFKPp
sFINMbptODbaDn5WS7aDnJNlWeFrHMj6FqlMhPYhcst+DkSPVnB8/X7JUGtjlqtPnD1dgMWMSexJ
e/8z86v6yEJIn3FlQq2ycH2kFzGP6S9Hr9DycHUUtJooY8vSGcelEGk68zNh0sOCjhfJ+wJdhc9p
lzJWlqPrONq7FqxAHU9zaJgwvp1ujUSTLMIDD4UMHEwFJHtBLHBkFm/YWul8kYu90nOzcvII4Dbi
FAVDQYG+AicHtwaeEMub9RIXg+iTUofzEbIxawa2D/izcjhtdal2Y4mMjSCB3XIVKuVQeTaZ9oZX
6w0YC4A+BRLwU4QW/lh1uvROU98STwK6GQ9dGwg/14VdW75PCGPyb5cxnZStuC+yl6brYllWnwfI
fiYP1ywLFCrSbbghiW7TVgAVHBfccTuAEczoZXfMWnt3boID1o8YXjfLI2JUEOD34Yw4jKtjITaj
IlUWg5iq1/rWBbPKjt1jC1kf7WMbruInXNjo40737FwouZEsoFJIj5913amG79IDBiHqZsKcA/B8
WlnDyZzHWCFXrs1tFIjOPKLH5tcKz9HAFvRJCG6Z3XymZNJ5B1jptwSu765PDP5nWAUUDcPeSCZV
Rj2WWSeGa9Fi/oTP2K9uTHfsESiEYx1Jr7fUAiVTsZDzB1+64wLP7WeMVq8DahLR/H1Y6CEqmFlP
YLbk6ONN7NK9UP/0tcl7LJqmhM8hqZB4TAduZnc9VPjdqx92zUzaxZltIbi/RTLKNgW6sA+hjV9m
jD39abalA65Zl8VY5nkkSE/D7PzYgTNuMQJ04XmCbhheh3Bzn9quFiMsHqICM3lAeHTuqzE4jyoS
Fa202p3wTqphtdtEZIsMXIJJYVMRM6YaAFzKokxo/1H5Bh7sYHGHtWjUk5RgJQh9K4ItB7ccw+sz
Ikd6RC00c18ngLqYo58y4gcILyQwTwBUR/ibV+px1ZoTHGctU5xqdhGQnQyIFhURHvNt6dAdiIcC
Zxo4KQlFc7bEuP0TX+twhv9JuRt+ANduSB4MMX3ONdr7OEcY+TXH5afiWkDgyoviygStaOhgbmMx
R+m/HXHgcS4iAOka2y9UDEHjom7vIEaosSqztEzrXSeVAg2Xz+WOMBXNiRBq+1uIo1a5/XBOODSa
8/VNGVbtfceP1TAO3Ov249fn5HEGk8OvB9hS2n5n60bi+/BxOK1ACRzO668o+OeB6njk4+830DnG
DUeT3WzGxTAqEbqJ/IMQpUSVz4ajwlN6jMmHFGrq7GTF9JMWHVa03uIaX2tizI1GMqQv+pkIe3Sm
53jogAWqf8PHmMnq1D3dRrpxvuUG/QJ6IJwDrqBvgmBbgaGFCH671fue8jJB7vrKG4mhVITUnJO+
u+3kbN+3g1X6jojBDEcgdszBBKDrZiO1gOBdeXMQYla8Fb2jVs/adpGHLb5OmBRw9VKqF2pBtAIT
zgB1YhPIzB0doj8kcf/iYvCy2j+c1/3bJaFz//qOlv5FNJe3jjkhcTN1ar+dK5oeHQkN6irjoERT
UfsuY3g53TaadFZ65EnF94N1fU47kaKIJcVUTvXpMQlks1bTue3rYF94W/rNf2smB/6MDpgGWppa
0sigQwVYihh9W1YrmxPlSB7bVpOMr5+s5Uiak5/sQXW7onB4Bw+Z4fxuQpyuHdhXCRbnELvHljgP
eE//HvX0OwvHN2EzIM0V5td7BVSklywS5yKHIeBGSTGS5TJWt9lr+Xm3v3RiW3rlRlY95VDbt3x2
hOsbMqvkYuBlG7ZhvlZzqbwvbaJID+piiE9cdrmvlVmNPrP6lUijq3ZHePJnax7IFZaotvIZn9SC
JoarOaqBebMvENpX0CUGbn7aYcNo5WonqINGu88zpG1mKcdP0zmm0X17tvbJfzY35h1mYrIkPSQl
dk8NUo8l+l0eFSyKm0eBpwNKSSWrEEjkRk5HzBhgi0kGo4v6PM318sGGYnJaGZ//3LiOGSU9Ztp3
xsQbidA6Y/o/ykSht3Lq8I0StMw2CKdbmVYf9dAjv8BjPmtSQIM4g0lZ3t/vFZqYP+w8cgW1mbfH
zW6IQ3TaccsLbYVFR0wI6aOlhxtC6nZw9x1C5OfVLFXUFzEVyMCY5ib9B8t0jhAI0rQVZvxE9Y/7
h9+1q5kwYTrQGWWXsubqiWy/6u0wS1t4owHufYl8dcggl5mozYekm61BNiZ2WQCDdfx/B3mdR5eq
b9WW3yFTvgPxr4Vq8Z4WgjA64+Aa+b1/XKpvHzGlZM+iar/SKtKbt0AnI6awPVdDsqrW6iN7eRLI
GMA2d76z19uKHieHmApQeUXEFEJpNLsFXYYGqqwwQWj5vJUKKzPyBoQi0fn83fDNtHssCoPgDArM
aEQCp/pa+zY/BF7xev6jMXnlIi+YPpPbLv4g2So9suBfpVNHjFvwVtEua3jGVm3He8aBN8lREoDb
bpYT7hHUsDoIOFs350pJ8BAWaJEFrMsaJ+hgSDLU3lLQBLCdSOWYNErJOOz6YYJHW5tpi2WbMnxz
F/JgxriZcJ2Ynr1BbdARGlG/iUPb82OwhIrAZLsMytiRpxt5ErH1TiMDqhkkCe7631lqQ4BGeSYD
s8Uz6/HXMKS3UmGp+WTf3IXgHxXKFfZNw1r3PFkEX4uFaE6JSxlf60crxM5kSGJxJPDmTr3appKu
9ZmjHVnEqXJRX5TOmk3OISJjrGQqKXhnh0SSAYqsMiACSiHOJmf0f5cJlKcfhIVNsP4MU/ydhpUD
MYdZMNg7D3b6CuJzjoXNHRejRSX3JqLe+emi1J2DcnrO7QD5m6DQKdqMnW7Vw4r/Mb/91IjI79J/
RX3qDlSiP5siLlg0qmqQ9uAc55Qm6yPzk+gBA88KGrlw/E9FSH6tHBE7KPKiyos8YwjAlkJlyjgr
pXVSwPNmqi2ZrIxmgqSS01ZtFwspTx6/txOb2RiL5ulEEEwAXPNESvk3DUKtgyh69YyHMFwJrnj3
Lpb6hFdr4MXZ1Ii2MX0uG0OSDt1hXAn8UacRgse38BVGqOn9xYw8ufC9x6jVmz8HR8YvapP/e07M
yFHDkgdUSDiwJJbuwbIbKE0vxD5VIx/bWqHy3BVRs53tL3cMfqizQKNla1VX0z/UKsbu3tNdLL0f
+ARbHGCOmQWLyjAVoTUmGsgQbmPaxDkGA9pbCXXnLBqRi1UE2KMwuiO7fiauLplZyYPWNVM04WkR
E9k3gPtWr4DKdlpwY2lPO8t/FBGV+Znc/r9v7iYjI+AVTKP93Wsp+NjkivQZFy6cNrHrNTWa4etI
EDte85QfSlQm9kGPrcDpAM6Pm/60w+J9L9KKCeBvNM5mYY6wfVzonMUocTtg+6E5n+IR/Yh9glMB
NGr7JHnfSa95PAfsXSZbiz6oejDfe0dShuALWHmP8+KsMee+MW+HPIg1pm3Qrbf+Ezbr5t73quSZ
T3SPljH9LkFchBFD6zn5Fd38sAaiVspIF0ZPaJa9t6+aYQ5s1l2QUJY4Rs9STjZNCreJaFmDi8di
8CYh/UHRL0bX+sLNyoUu/+kl8+IEdhDUIcr6gGsbeJykGjHN24ShU/K4IWX/kUVKZaedIdq5yB99
aAq8L+A7iycx1xCx3uiPxuEjbNL7oit9yelYDyMU3R5Nh1upOWNvxKGlabIU8MsYNSy+OVdsDZUh
86PTvI5TXcaTNmDo5pbu/PCn6koHrv2dqNKiU1sk0aJkjpzkCrNiyYyRFFX/gJ55TNuQO31gE0pN
qOXVDs/eG1KkZPGyeIrXWqJDC2H53dyOVHOGJO4k5ONIDoniNe9sqYFGg3H5mVRa1yJQow56PBgK
Q2QEWtqA76ytos5fqGnKrIHe5yugHTQyBtyKBwbgICBZ8ga/PqAPKdMiuN9vyXWjGnL0R2V0afbB
V6q7HycyzTcrXm7ugB5kqJsjPtsvYrS825wBaKblni/VTk1KlSz9Rhio3wOPh5+8yhX9FOl3baXq
6Vz1pWl/OgxaKlPCegARX5qCv6eEDwA/5w14wS7bYwXVgn2LwRH5Au7nPNylaWBc+fuYTARBnfRX
uqQcb/HILJfVMH/bqaHfWFWQEZWYWUHdsF5V25EDZr0TX7dJfmApbCm7SVa4TBNbYfLwgIdWNyXl
fdzW2EY9TUZx1LTt+ClZVgf051PXswvlhtpSx7zow7KCfbEs44zRGosfkRdWh8pwvu+Bvv6yOZOO
jWalsu6A+5oPila+gsVGjOHuN8vzsE+fsS5/sz0TV17mhqJ060ZZ8R9g5+pJlMezfz/MBUR2InhY
UlCBC5RQSvEmvSX4s8j4L89Eo1CB6UCqKeGvl5+6Gybcj/wOdjJYYttnv5gY+R6cAbUdTXTdkUaJ
SnyUYMj8UxVv7vZ1U9/9ukPT+G28PtknTGcX9t0ABZ7TLg6xocOej2qPEpeQp050dU/Tpmrh91q6
rjAA2H8iy2f3/nAjIHJumroyEBAhy8Uc+q8OJCDiezemi0Etq/JWdWbyrlPcZjn5xouCQ1jTX/mn
humORXBUpkd8I8agYKUSy+u4lT8f3q1EZXy2q3zKzfDl8UtJC+PMeM9JQ3FS93ukV0hrQs7/CKZj
KKGVNDb31kalJtvhK9t7IhypgZy8AF/S0J8BY0cd701IZe2LAUPqWfk7rlWT/aAV17Qur2O7dAzP
5cyuFxMfGgOdN/mzv30QGuTrRjGGEa1Pi4Y0a3yIBRCVHlVjb0c+DYQfr2qQinvORP/p5DP7ftW+
vHBTUf8gXIqVqvbceL5TZ1M2HWPpjqms8NNwXXN6vHsnFRODTcw0ldMIkXUoGJ+G4Bsr0b9XcdKk
Llt3PS7ZLEknOklCl4nctssyJoc8gzM0rjTdUVMBBwjJdGWV0GUTA76bnGE1J0d5xMe9/EGqWOxm
tonuSUlDQKYWQlXys8j8R99bcjXeYmFVhwVUIQwY8btkHuJ8P0R+AJkfqKJC8dbsyb4MMj9ncGR/
xru58GWjda6pWmWoxhedOOCkB71twDzv8z09JK9G0kD+10m5C5A8MMeLOWLWb0sf/4P8yX8uF56Q
5fei9mU4unKPKR26g31XtgKRPT8dQLtwxIw10ewWeJLI0O4ljOmgI0zvizGPkw15OL2VVmc0oQ0e
DVqizkxvVqDKpoDxw95cArx4y7vbuBnLtFhqUaltOxHuKn0d7/X/2r+Omx4enl+NKfvGeIzLa/oP
Wg3FIcv/kVB7Dz1CcGh7SexBTLLeYUmu6F0BZa4AKtvyvXsGNLuH63KrpCa+3qWEFNyWlCEbmUM1
41OYn05afh9wb0i0lGhD4edjl5SLMggZK9u+CtjMyKxa4R7EcpV6wj167Jv2/NA3me43kuf62VGv
FC8SygOIGBQ9KsQ9FSxh9ZRSnV8jUc8diYQMGPtfvkvLU97F8e1viX7z5mKYxEaq99R875lPO3nV
0ps/Z+fTQalo8ozWEkqHB7bmfcOBdrrQXbFocM5sIQPgwX9LgPgDpxfQl/kP3OC5vvsoM+p7K7Jj
LuY2iPtWkWXAXWddtc0A7q/g52K2/23hYU1kLzkK5hF9LHKNXZolwdwcg8HsJfFiojekqpXizWSD
hORt1AGjVzhoOdU8x7/eTWlUbXXHXfGWTmpqzLzyXten3gqsVNnsnmnTPtc8hEChbybeiumaDdfZ
W2g4Wn54skvRTOWgz50zA9tLG0W+hJINbmH9F5IgPnrri3t7BXkBueWygZ0j0bPZSQOAuEAR0v2f
wspRcdKL2tOgK+QgurXACU917u4KoBCQmJzDWxxzUfnwkxFR7WSyCBY+V757ZXOJOF8EtjzlrQXE
7ufO8RSaevFgV3q988G110YNtsetetp+vCRFJ8ZBdA6WaZ9QL1Nvk4HNFiPcltlVn39PicqTikO4
+HT0IK+DRy/cq3Xw8D1lN+Rr+OjfdiJ4WFTeJ3QpcZcynWyCv8/HocIyujA54oinyNpx8ZhPCxc3
DLoakBiG4vBqRZi1jTXBL7ASwQdGcPblWDxAgCt+YciscdojzOClUBLAXL4twlyYZ+1gxgQOMTtE
q8LR+m1wRPmTffRNOBn2awpKTovoLAcToSIWrMpUVamHudh63w3rGySXTqSxNTWg7yFie8+y5Du0
dGzMpOeD8vux+SOfVllip/GrY4H+QNAalMfvgv0eIWtInkkQxS8XoYU2+Nf0UKZV9YllrhOsYiLs
87d0ZcJPxtUt2GrrfWU9oaGz9dj4jgEm7oPC90zYfwUNRTjDvixlNZSEHtqrh8J70n+u7cfekzE3
X/cui2Gs/l7pC8Wk6HP/3gtUQb3c96Ul6JIFbV5u1ZuJB7E4rl3LM32++1xduhE9/CSFjHmHeK98
5mafEUu41argHZDaMtdVJ00F6kewf1iBZBcYcQ5ktF/a1weySrZ744g1JG6jrk+Rg1+uwMY+lSsE
LFHv1JCepmeybXWwZoSVmqLTh7YMs3PkTgsBOGiVBce8LPIXPjkkzIF9YgztfGk02xwr92eEsS3/
vHxQgskWrnH3DhBo/kmaO5a88qBaBQnZ7+mkL/3iEx126mIj9DxK2/LPjZnBzPAvhEuE3zACHKzD
F7X+5eTmHvnb1VGVrtsEANMwxyv4e6r8HootJtGgXk75FcXJ77YiH7CP6F+z0H3nR04fX4nhuzwV
QnzKEzs+6Ig7UIzqa4VEewhuMH9inc4vZw3q4V2Yy2dZX+HmKYB5dfpkj9k4SMuYgKOP04Zn3WXl
1IN1ookDf+AxwvqwcC/0qyxMfPGHdfqlJUGK/h70YxDbB5Bh7Rej99JyuSxR4kwugNsS0d/bflxP
QyKY0zmOr5glAtmc1iL7pQFv6auTVsSaMCrHcBhNigu6QkR9R1uY/UdPHsgARUn/dNFj3jAKbFJY
/vZ5CGKpaYfoQgIbMQEvo45fDwXTb+0LHehOIFZYsIq4v8iQ/bv9xVDszt2fS9O9SaGx2NouJnfr
idX4aJEQFmqbym97bv+673FG8Yrx9JrG5fCfLcbsIvwCMteih7mJ7uuUBskohlx+lPhPRM4fVsjN
hOAuG8ZXDGB1INS8IcFjjhr4w5ZWv7IiN/SGWu6RcGH0ouH9OJkDZtMdwJHh9X94lJRXiRwrb8pq
4tepeFb3v7oYckDCVo4qoBdGL0PagOSQKMtpx7tdVE+CbRkx8kQKunoO0dhmha5yf1ufK2w5BRea
xeNDU6ns/a5yV7C06S1VMb59wyTaPJy0VPjLTwRZa7rIyWEbWlz6WkdcqOBGq+fTyoJRbjBrBiWm
hOudNRyOUVExlyuybd2lkqBZjQnDdMdfW/8GooeRFucTX59IT74gNiZg/C8rRY40SL+pkNHZhOQz
tMhKdYjPw/NXY2S9X7anOJOQS5uiIzfaD7RBAALSDA0qveM3lVBDIn6Wn+3AdHfcL9RJYka99Tuq
u/HANGSWS0oauvg63oDK/iMYRcTyEhvkH/E0+G4AXtpDM3fduSB54X59Won1J7xdJ6sawbNuH0Cz
Zy1OVtKMIAiL4/6RAXW/SCJAScM8fwvZL47D9hWiW/GB4JkHQ1XIBwNWfmIP1N0TpnbzovAiStvg
WrCArC+NvPXeZ5cY5Ve8R2nX70dO8Jp/h1Ud7PnnyOsR8ZRPXqZrUo9U+lC48paDAb1cOVy6fF7l
grrdWjl9zGoxtTWjPRpfSTiGhC3W3W3b9gLm47p2yYVl/NY3nRrOYk50DGMTfvOFA7T4PIdUZ+AR
hxdugGDVV41XP8fv767TzUFkFYibVKwSuWKlQ9Dz/WeAa6l+amaI4hf9zUMhWURPsIyLTGCQCMAv
dKpKKYp+d96fqhHqtQwT/Uv+s2rxhNSDP/NJct2+Nw4oVu1hWf7W4GJAFY1f5RNtRvppGX52Uf8b
sI2Z83GleJeiMZMfi+LSHpL1lV9nNgK2nurNwa+y1U31HnEFQ9gAnV1NcPI/g5pLFFzxMF8GvLtC
2BcD+47PGhgE1CMd9knkwFIqQBRVdII17xMN2NtGn08C/nygyRSRCFDDwXYlxVcMbWkd4zTc4bcN
FRU76dC+4Ra8TRCGFNm/LDMP5vzUWLtoedsas9feJ1EGqGakskTxWgvWJziXb4sjJ3Z7ExIXlKP5
SV79IGMzxajWv/opiADgLkoEzH1I6CO7Rub/1u9lyd5/R7vZYsshZZHnUXS3zT6rQ1X0E7jJtioO
oHKu/SSqpMx6SjEDwhwNBL/BupFCn8vVFQrMF0HpioQNNTFmadovFMo5NKZhdewd7QuP8dXONYm3
yzyd57jqDcWA6UtgqWurvwxs/irXdXvk7tTNXOafByb1cqUs67m8sPBRVclzwWV20rpFk8W4nwJI
MelqHMJMhKxIhl+sHva13fSp/dyVx1xNqONba1KnKYuRVvYKubwXjCQ687rY8uDBvlN29DgtLeoo
oD7uBzRsENdEm4k7nThvc3agjA3DgT7Kroi91ZnYW8iAUmGuRxoky4/q4dP5G4aWuwoE1kS90fPj
qWQM21xI9B/bGOhehhRnexxtgGi/iZlo0dqXdSHHHwdiEANeKTvk0YsvghOy0YTscGtQHNae+aoR
4Ayh76U/rXovaqL2y5XJB37K6t9dO4yy3T3vaFkFXzS1foq5jrVC+rGZShNsVe7hSrLs/R0A6eV7
SjUMj5teQ567N3e4mUvgkAJrPN9W51FsSs0jFbOJLJFQ5tfNTSL875wmMCyXZLlHlHvQkVXKUHMh
f+MscJD3ePpQ7Ca50/Z/OFY+j3U2gkgwssJGtl2xfJKUb66Pxf9jjFhyFS+jN1OoOuw6uUL2AFh5
1DoUdZt3vpeWVWSVtkdYshBO6/URJyTp3Z6K1JrimylcKw7Zed6Eh5FPSIBuHHyTl3s+e2pOYEtg
oK7jdq6Y36P3w2VDBXMFVqZBA5oGnkRFv8akpDOhtYaF9zrZl6DMLHgsp+ntRg7Xxriu2HaVawES
XanzIF6f4/nB56Cl6EdUsdoH+oQZ9hYWtgjg+qcOeCMkYKKwwWJgJsAWl5iJJzSeoIdww703cNpv
ojYyQadmYDZMUVJkrmSk7Uhe43cr/bYSH9R+p0g1q9BycVAYIfPXF5Pe6jFYFjWjX+PxG6DFilh3
89WPNpBNr8qcSNzG7CQxnSA97mILAyA9lNUh+qZ1JtcPG7MC8/adsPziktl3s0oY5TnQmwn5CUHJ
1RRPEF60G8mbuOFXrvZSaqF7oFxO5+ZC+PlRTF1Ubc8eon8IMGrEbkKynIJtHUZ+u/XMdyCjoBDQ
qIJrUYMp7QO9fnOh3MNTs2G5X6pavtn+WwrKKHRE2RekQWgaUQRIV5Vq4m8nocv0JuSwldGryhSc
bdrR1m81/dayGCZLm8R3aQ+K0ZN8yWd4cKfipe4dJnkl9+GHUarMOv5NiDdzSjK5RtJD3lBeTuMX
3RBWnCkOO+G7W0WHx3tSIt9HSrbBWI1u2h477ovB49NNShkuHqpSQ+mR4p63KNRzGweylZacIirt
diOoKNDYVr/bBG9XbkawzhGxC8CptMgJCVOpx46rI3HjYaD9gGJcIqWJHPPfLm0wEBu5SzON5aPI
ZPPmTOcRiBR+O0zxvLoqWHaLhtbH4QREjl4rCWmgUJ94O+XmKtHT72Ezw/YhlHQ7BvxoXjk+UPQL
UgIyGw83jBN43MPd/YI3sxBYinSrE2pdNlJt/Xqcycux4QIlClB5H8KFdOYwhTudTbSoQ/L/y14R
EBYemNpgxl/9zx2UYAOpQWscTv0+xH2G1oaLgPbmrDFLeV71PJpyHCW8qCDgdpkMGvWY5qlXbrh8
2MLabTq3rcPYB3R186H8jacAB+DYaKwNaqmTx5/M3V+6VhagNap1n2MrKuO5YjzKE/f3H/nXxbxH
ed2pCzo44Of65ecg7pXUFjzZFraFv3R6BqhZ2Z6VUlJGabZFXg31GF/qZQTre6ahO1hNJXy5pSkT
PqDnHu3KNM9CfrPcCvEj+gjxxR1Wy3Z+dqH6n8bZxevTi3/LazUcUuJkPe76Zz8lMQ4KdrZVNWNA
/OG4XgO6eZ/oWCHOhFZ7/21PGYPWEGcnEBsVEl0Uji3XVo5JG+mNu1tVvmUymplFuCdbpwfRPidI
Iuug1q9CgvT76I+a5xspQpw1CJbCTaazRNuzly4hx1kUE3BHpGdCZAtV8f/utBT9nlgcU21JqIfj
lebExos+cGa+io9kXwCB8pUrk75aQYTp6t4JU66WMpYrXQgeiPHhuGkqD6qU/NwgNdDnjmoDme80
gLslKnwH/3e+LNTsgI8XjqTXNCcMWFKkjo4ivaPJJ0gpZgMQCyq6owIXSwteyHxSYBQIRNgT9PFn
2OH0D/g1VK6Ns1HdgYQpeqENaElGliR/edOEKD8svWHQA5dq070Qq22CzS6jzNMaycZCh7oalD1t
dHYoJsm7/TIafCu16pKBNRFl212d5AWW5fJO1mgEB670v8VexEHOnlzz0ZVK3NTelFdoWUYDxCis
nrunKhogYaD2m/xk8/Id1qNTRIrukSQIWEGZUUT7vYTB/x5Qlvm+LESm9djmc1nPl4pso7QRCScr
RjT+nAlR3U9KkDJ44oacnpxqPhX941i8AgWp95s66d5gz8TH7OAIx+Y3ViTWX2ngUkwFycUZNiK3
RaemUpIOLu2HmoVNwCClHID1xc6DQXatFsqynpq6S+Oy6iI43WxRcCjN4SLTynt8TFyk5eEKUFLH
NhAzmFTx5yiKXutFGWIHWxXwJZmZQYU9kFlGAF/EcUDooFNH1WtMdOWFQSBfz3KzxupIcjQutllU
WkTHegM8IR0Cmf3W8830YHI6PGC1HmUlfIY5gWc5FCTfI078DwrEzz5Lm9QEel5wHSCYpEfISNwX
DzG8uPET2OUD/UMFMfM9oqHHSkQQrtKFxAuJTHpbzXpimJKlPQjqihWjHwedW8RYQbsVWL57K2MY
DGVJ1Zz1vw4JIdCr/Hg7SDm9PMkYHM6GAHVuGNo49gGA3LgvRrCYBVvjW3wtwzZOhlAamu5co2F6
5pXmBTlVOlifpETl8XBIOatfclTgDFqF8BNCFnsgoeKNHDMXB7ZaGTt+gt1kofecTvanhbklus0d
IzGI0uaTtArwFLaaioQM4aCzZXcrhXC3+Vt+xezy6YuW5TBk/49U7PFoXRpKODggH0WfRk2PVm8L
ecAfRittKioz22tyK4awpsYTD6e+OQ3RRanZOrt2UUH9hnOqqcsTvqVRrt083226izPFFTJdMv5O
33XvNIFIFpO+ATeDuQ+fcbQPkZinEPU0YY9sOPpEKJokza+dgaMNshWbSFxLoOpeX/hvMZEUNsi/
VCLLjGVmCiUMCiMunljOsXdc7CWFEE6jP1U9jWhdb28dnp7hBJHkMlPbPtHjDP94IuwZRWFQEE1Z
CJqs2/dpwNqvsCj/nuGnn0UmQTerL+h8RMnGUiio0If1NaWIbBrDxpToNesb+7Ylpnyhc5rxGF+J
HwrGSHTS/hF8akz7aF4j+wk1QGWI8xDzOEBKemOjZXjyHiP9uJqb7TEv6WaGSETbI0Ox07qvpgUR
5HrKb++HSf1Lrk7+x+8tTrmLVhPMS5Uc4vMs4W6RYxEVJV7f6j4XinGX8yQgqCElLxz87iOWdC59
7O6pIKFGNSX9NqnO9JxkeZUCiiKfBMVLrTrLj+P3as2EP7yRnKZiwl1BSXp5MdoPXM5KofuCRgru
9dTlP778604a/M9bpgUhzQoFZL4lgGCMitvlqAQdTyg9YoFfkk/XpJSMLJf0d1DBwy7gqVoKo1/8
fB/az+DfzDLDoN+3uytdVHwekdjhWxFqInjky2TvrVd/N9/G0DEOwn4AMLiQ/d2+IwhdV9a2Ml/Y
BQ/UEW8JtnULTjwibdUMTcPrpBMCUDpotZfMaAWSxIPpXMLKsqvq78awET/3NCm/CWbF0aQ2iuGG
MYDrlCOR++UhcMfG9Hw5xlw1AcggX6Q/aRzIn+/gnWVqOEVjkg96ea8eLfK5VXPgHb1HcQd5+xHt
ORFJj9nepz9QDw3ITvbIgpYBKoHsyEK2bc9dEhKR6m1j/BNn9c3wb2ClHK1gHf6Ad/7ULAzsQxH8
oetTPLrC1gkYYO2eF7D2hbRq+JYFS5OYtJIOme3a6/NALfBZdR3c2b7JjBIgBb9aqMOWsvdpZ4tL
OWV6FFd2hUgCTFab/aN5g9C1SuAivtQJsOYGMU7fIiB0twzoLbEE2u93WaL61oCtc9fscDzvNm0d
QyTiPzVchwKmLtFDmGk9rgsWaKHx1nECCoASj6QvHAHTK3f39TOpb6PEUU7o2kSM3AGr4OP1I+4E
waO+n/fkeSfQ1znzeBrTomLn7sBxk2SF3VD3Zrj452ar/nTMsL0EL4mwWQtQE/9h4DcgD7KVYyok
QdHSsQD658xs3i813zC91KkbEz2zsI8SAUIZtkG+qHeULvFZhSNpsAzmzcvrT8Amv3nkDuWG2qaP
3oM43rk9ZZ+mX/1ivSUyvS1z+JYvq/CrJYA+flQ1/R221J8YaFkaE9Q10Qui29DS8xopkpvLprQx
D6ukt9DDNLCu2Q+g9ljPrcFhzKN5eZHJTRGiOhZYI19rOwSazFcZZ5AFE6K6fQQbE7Uo/vHjWccO
V7TEsVGXYs7YbkJ1msJtxQvq5ybATYisosqJ/ymfS/bMLukcqcl+L7F4L7268OnLWYyN1ADVDotD
sPXhZ83qJ6cq5/psuE5syuhDEFMyHDG/+dmIVMrsucrjBXtSfmau+MOVIUfbSQQk7TJ0x5P/UNkl
QC1Xgn23To06X3Cl+Bgj/wK7KdIu1Uu3iazLt/e89Ovzug4n8mNCcCu2pIutNqeE+6T7dhbq+8Px
Yb0TAu+KyTB0cxpAuKb2DPmUcQ3dRklJW8b7YnpyOjVfmAwujoKSEXmVzWNv7d6HOe5QztNPg1sj
WF8aRs0NyeAVugDMlAMr2A+JuEpp5PZtooeGmP7uS/ZhPKE6xJkFAbZWiJMHnRlFJZxcN1THVdrv
/A8Mdragqeasawu84laKHmPjbgN8tpiblwn1BZ3LPOmiVQHVJ8WUpXXj+cClnPw3axmI9UNyIful
HWDrfBnUZVYWC7xEI7DzoFUzf7xRUxmUqkgQdCtGb8fzB7H9118t0AxbwZk3PAGKEW32VBhAhhaT
+wsdjAMCNjkPkp/W5SoWCGfLD0Y1GpwmgSf48yU1hlqYZIqd9uPausROCKKDb9Z37LAFE2cFIaxf
Nx21J1c0Cx0W0/EeYTCkDGcLWBjwgiNRGHuZMbUx2b7VtW2SDvKBzXLO4l2Edj6p9I+eM5k4cI+b
Va8jv7OnriXcey6y0QZ3AZMlC27y6echVfHQC6BAx/dkUPkkaugoKQ1zkWe3TnyQ2Zpx1bkYDP1p
qGTwnDA78o/9+pcXSncfr2aQ0xXSFPbefxxaslurE686vP1zsyVIrOm0Swa/xbDLP8jMEwk4c/th
6aDJX67B1PRXAhlNOezB5xEVEbISUTPSW3kDISXJC27SYxXpp/atOcU1Ndy+u233gsqUjM37NpEq
xiBMzEpVqTWFrSeaffXkqWvv//QQ6Nulp3GsXLtoMdZhKRUDc7X0akJvP1bWxibQs/jfSAn3hBuR
KWU0Wr3lXeERWjGl3/v70OZGk2PJ7IvP+Q0R4xKcyjvzaO8ZfwlgY6AkkhUk0YzrPOPcTSNER7VQ
oxBllZJ22mWx8bfM78TbrpTNRBc9WH7ccGq566MsKowSfux7qDkH/uoT6QHudjbnN5JSBj5MCCN3
JNjcaxygGzvypjTKjwYfGzHytuU7jnJknySWjtTSnwAKD/GqNLbTYANWQgkghe4BKS9nsMNzFsU0
obI0zfxsQo/GzkEtnnEoVkmumAIaQ3absOA3pjrqv+YTemSwhh/6TQC60gmGwQPtMKIKIcReMQcg
1dkF8CgTizH6WAYNl0WLdgDGsIAUys1HlGT0q6aOj+GrjbvjmQsPOGy3rBKUv9AP8R6oIBUdfdI2
elhwpbzCDyhfWaOurLJQuqBrM9nB4XdLo8OiNOtQobAp3Ey/0WpLuIDkWUP6+vXsqWYfMp4jW69u
jhAi9Lv/9DHyGee/Z27027o3loVQzIspI1wRPwcItBtGaiTWJDamta92Tb9VZp6bv8sbTuIw4GBy
yWYg8mniVVRuZXG4ybaOgH5TLL9CvQzJPD98EohB3VIsPhRn86yd7C9eOomAsLcXiHjvw/XofYjd
Y94gG+DuKgGT8QBvBzsVEKTYwLUUlkV5v30WTRe3TE4m0R90K9b8g6hJlw7e/JbE134xZlfWlT7j
jYugoc/D6JRKxpSnV2Sg5cwANPQP88pFMGmT7jCFYJp7OlqtFQJ4iLNFkhTOtyV7v4WIe95XlEZE
1FuKoi3ZS/BaTphmtzZTRbCTBB1E4Wtl8IkvVdqHSXK8vxSp+GB91rMEnbozDzox2EVHNP+TgUw+
mSb/Ate1c9YXTZPEPOPigQ2ekQKj4OssR/k1eMHJPWxNzYmHkBcX47xGu8qV9PY68X69F5apT6bb
Uq46aPqredLeBg1RbwNqdO9DBr837qBsQUyzujCAbaA0QwlKnRPah0IZQZbof58kb14cjU4pqKs6
1pztLsTFqT3DoJ35QSRizGfR5nO+9Z0Bqz5vsvNyBZ8YtjDROCk5+H08/6IU03+aot2HZh4h9+SE
OvczWeJa1xbVPaiE0MY2RlaxZTp6hWIWkJtLc+NDgegURk2JBbkXKLn+DM9YWFRi7KwJJUQXRzPG
a46QpgmEsD5B+LekwB13BfeMqb/i2YQ2lf9TNIqIglcHlPKm/3QTXn0p0hLxnH2Rmu4q+mOtas+B
5Kf2Svfow2vgPZDuOmIGxIPF4X0DOG3//wtunNYP195+iXcpRndwigZP0tgaa5V35m/A0yOS2sMA
xXwoLtXUGxBXNOx04hsvoeG8w1XRBWObiJhFjnZGjqWmpww28cJSgk5uxJRU0+1anMYbfo5AWxs4
+OgXMhOONvTy8hmm+LbzBraK6GA/6oOPhj2JWuecjH75MzOrC7A5EV13oiSKX3VzSan0ZUMSnPa2
Ob/rCloOHHDnXT9/FHaTnfMrF3fOvktCAyMZVyj+uQMuA36U7zHcZFFzvhk/ZZdpxZVg5ZnOE41K
Z7icEimR/g1s9g1rk7sgCcX5AiITZtw9g08dOrctPB1avHYxzNhnitrKEt4Jfdh4Dq58sXDwpGxN
ecB15yo8k9K/TUEHLC6Atdw+JI2zqnfFIOmpS5UhVn8qJLyAOTfgdGtjkRO4+9mbugrG3HFTRG/F
63PBXm4Q5lA+2xWvNHhxVkq0g+O8jBF9EBl9SQpQs+dDDw7RSFOrZYWjGZJg4nwjfQLNxDJhef03
f80YNiK8fhq3Gd+KP8gTIIturP1GqgOuxw/YD+kFVHDzb8VDzrB8w9f9h1Uz+/6070uIuXpThVxb
9iaNV7PJKm3AcF0m6zdFuwYvyh23WmrVPkKk0hud2ffZlliiqfZWsoLKFerhvnuERHlEHtzEsxKi
NZL1YTLRJssDsZD/N7nvPAmF+brBeAf6fJNbPhqO9/rNOBk0HZJlGeh/Asdmmwk9uvt0Iuc3KY0m
JmtOYP1zqTKDVJVKGyBBQJFHe0y7IO9ZD57nsG0XU7iepsX5jQwaCN5PXOSJF+QXmkxEITcYgc4n
S9SjPEchSNLwa98RU00SVXlM9lWxbGeL5r637B613Gcb0dX9NzlnMPLo37wxgOyawAtC6PrQAHbk
QC212NDtvEaHmf5JI2tksec++vW0hkp3CUUDLsGQ0sPu+7sXpbIevBPddMvyQyY55gDoKa/QTbql
HYRORyc7cKLtTHnaV5fdfEzCxIRBqXBp/45GyTPVZJ1QNONQnrRBZPOdwAeIqcE3uIaV929/Uigr
F2XaukfJD/aJMcngtju1J3KNJQ8SLtpf5XcwzWkGEfK2ywK3wXJAdaglBOJhk/lyhHtwt17RFHmk
7KAKbiyYz+7dMLUhwwaQiy3sDl1bPmhRtcSjTHtFax4FFkRePJcRh6UUL7Ew1YhUKZCvkCfhk0NK
GNNBVOPEEVtWnkxinlzA6gEsMeSEe4XXWHcYN/dANcEwkP/A+1Iudd5eHxW3iKrcwfWCys2IVOku
6dzcELrsJceJTug0nVMmvZx29YcrLCJdqXZydllOoc/NTazxZHTkKFQjJfZsI2uS8sIrjQNICfuo
+3E4CdcpbrzA4XguIw+z8YX3b33gGQJ/6S8TdO6OkHDrztuv1oO/umCe7huXRg5KJyWqUK9+LZRe
WDf3/EBLByFwfURI8Jdz6o3Izx/VUQANd2mymTWSi4ltUnRuyRONQxke7O2QTrjmnoWz1/3K39rT
0rimY9pco+//lrX8MrOSHvFFj4qE6/ZcDSFXbGh1tYmUkOKrSLp388M/qdlwB1xlOXv/qRxhIom0
S/d0IVCSt2G85Mf2M/jo2pst0r7jVMEEbbg+lwvou9Bpu5jcXhWWfFI4mce1yZXE3bsKjZl871c7
7Rb7YtEWHf8SHiCTw347Owzse2G+qX5j89aSeAk2GWycK7Q2yr2G9gA1YlgpuUooLapHjJOujocz
x7CaqN4CwPzlCnps0XCCfkLTtZTYSwVZVrlmeGHD+USXvqQe1kpGkNWuTIEv+CchAr9TFVz9q8u7
hP0zm8l1mUk68YAYLGDsRwbWDci+YJWE8CMGqA/YVcJ6BVSGjaZtpbRr9pqq3WLwpKLvaDY8u1kg
pkQILbTkJ/oZSd/kcxyvyi0UXiuKk37026UsS9tjU94L9mc2uBFBVQVQoYPfgpaZ6aohm2uuLfot
NiPR0Vkfax5MaKT2rLj7CeL+MPwlWDJ9aCsjtOEEQwxFV56+HAmuEW1UjxuvMBRBVmUBohNZsdEu
9/aX/zBtCtyQKGkcL0erSwpUKV5YG0r4Nhl3MHQWqe9NN9DuNHSost7Ss+nqpiuKx0mXk+iqhxVM
uhf+ORBJ2nGHevIYkGMcdP3cg8R0zpw/1LQZ8w2UbZcTjoZ0qh8TtPOqz0r8xmffViRFvcvZj+PJ
961k3wjwvz3FMsrSXn9JtdvFCQvvibzJQRg/hBp5AFsYh4Py+CizleJu3DDBnygTIro1eeivc9/f
3QIsWgeA6Ba+xY93lST9smNmTYP5hUrhzvWYZ/0G9Jml5oUgJsKXKwYWwP3YnF6U4dsvxVTDxZxo
FIMgqFlEer3BWxuXuoIocgYS46p++jKvLFgx4A/MR6b2kFZcxYfGtLayRotqpGcs9xLVEFQe5ums
W5gvv7BLKnz8GrncpnboZVB7ggYFB6m5kYeqK5j9rquCaSMsj3UuFWA6DOQEewoSwlRuUzQgPpR4
zzbcOQEudi7lTKa2ULDAiNBgiCINqQJz1HOzHn9S0DQ4zTz8leVPv7gI/ui9F8qAkCBt0ITHFh9P
70GUdpxhSoX3701S2gQ6XMnz79cGh8008vxIuhGTj520djyot5dOVlkBOgif/H/S2bSVhIzDwNDI
LR+B5cTfk9YsrK9dhpre8bDLzcKPkEwZJigCh2zOqbcjX/Bo/3S/YHEP2tP1zY0utb5ktInflj7n
cnk+1kjkl2C+CglRllgk7+JwEjt8rdKsZaRtLzUo6a1IPKmpbqJbyLHLTMaxdZoaq2FGdxS8tnZO
ArLb9cVWf3TBhyeociCJTCc4WkgVu9r85Yr1uSu88F7u9AAo9ns7uQvz72Eu9IHNexISbQcTxTZI
j+Fk+QVQxnTKCtzj7slq2vLQzCbyfGdNErP9f78CNAg5hT2GAhde4Vw0VbgUuCGFc67Y211onMUy
GnUVMFrDO+fXoy0WoMQM0FOIRuIuDqx8R4vt0gfUQwnQc/kRUDizrBvsWE1UAndobXVU09Z04Kv8
dR1j+1UyMX4SBCAf9exQdB8cGW9CBz8IF7K777wm7Rhn0aD0+Cb6lyTK7oJs3XarOh+fxaZu0q61
GmMWI8KZ5DYtvl6ObAebTLwLOIOFDWoxir22o9k8sragkCEDe7D+TMM1Fl75TaI+fQEnbg5zJdeq
hq1j3VUeIGHDyGE4i4/eGzDuggPGWzxtQPBcQei2jj0WE3G4yNVxLongNjD5Rd26SA9NjM+V2J+y
xCfNtkBWQizW6Ipbq5uke+IU3YIeltXzp44BoRHtt8neKp/z2IioHMS8mTZ7AEbfuqy44YngUbEY
I3qipHFmaM0PoAANj6PbeMjt/07pxQTwDtbwAYNHBopoz8BKyhuRrBIgDh0tPO3cXAU55dEG4MrD
OS+ZcaMLTkf1IT7EvNg5/U0KVPntckjYZYnBu5J39Og5OtGxlrpViTPI0fr2Hsn9xSuJ4wQHAb4J
N/Nmt/1m3uPhb5H4JavC867ZVrFl7n0DMF97xidjqNFTZ2LSGnxz7ZHtJ7e8hZ3LPjD0MN6HgWSK
sPIooqaWLpn+rb7CSScZxeafvqP3CHkYEsjhfvUGJaG7B9zeP4VJADi/fPmCt94s8q058zaIBvnH
rg9yNbGZzPOPj/74gLmsQXK+k2LkiWQDDO9KJuVhL9tG3tmEPSTAfSpdp51pQqHgG8bGj3eP/zsY
3TsnoqiqccwJLklQmTzY3z9Ud92DlZd445Rb0g4cRQhRURM6mBDzaAOjFklY4sWob6drYMUNEarS
vb+Q3VE8iRevrbhOFHNSLtQz5i2pRcxr9QySLnht22ZJ1BrZ0ZWru+4q+JyK7EtRcgymBrM3iPTh
LrhsWEtfA46Px01njdmFuvijJ+1tj1AFrMOhF37mP7k3gqqq8ZSYnG01K3kP0PduAqA/OcaCKZi8
CjiYy7XlercT6auBwDoRByY9XQW7F5qXjhgray8KRqS9flzBOt81IODEt146aRbqgvhRr3gwnHI4
VGXrx65l/Nw8uqqcVN9i3pMM9nGw4nbeFbDVBU8cFRzMh8cqyPEG6oUoU354yvbIcNEuc703+hky
TDEi5wnDH2xsY4yEr9Am4fjSwuFbbIq7g3QQ19/INyDR1qjMskPBQwF1XPfhbBq4jHJXwVHTaM6G
RGWTkFh5NkgSSLZWFJayfaz1wkoPrk35z4i5e00g9XZD7cjPhcJalm+IduDgZNb6TQJrEtCHcm9g
7l3XGTKzoxbAzwfHsoUFP4OtrJONhWQ17/gpSKLRbgwsI/+m8ptFjwFWdeMq98GHYxkHDMLJWVH9
CWUOc8Pyu4Dpk16nw5NVuHWlQUIbTuvj4ogRFZ5zKjkCb/7/33i7d5KyLkTBFQ3ohB+/YGVjXNY6
BkGxtEeiis4ZaFElH9RaTY0/KmVXUpo79rC4Ml/3inIs7CtB0aMjwJQApo+RQDygZbvClVWBMUqf
5nqte25+TlVN9lpeQg9nc60aICnM27YpGwHUb6vr131aa9VYTzKxUm+tlJijFLS0+bduufSxxoDQ
VBwMA9cO7rg8J45MJ3HG6AgyllKzhSLnIrB3uzHmDKXTyb3/pvGxqZgT4bwkZSaGzgtMZyhDEzMN
FREcOPjgkWoCafyeOnj8Dn9GbBuR6qfuUuu9hgdUI5H6fwJgEZ4v7JcuWuHTG3cg6PiLaZVU/Pg2
S9HmvEJaJSbT11jo4Ie7Kbh60Sihvz/7TFcaXokXpAIN/TF052WVmy1/LEQrSDmD59gqrlp4GG3f
rq+NFlKQk6frHI1o4atUQQU46iazRT6UKn34P79Pssw6us6X1Q7w+7UucNlDWhr0iWQB5uPNAJwu
HBWwqCqdme/NvvGsfL5f1HRYilLpZU3iQJ1opW+sEVddv5YaxtG0OgN44PFqih69RRBT0c4z4lse
uwj5AkhUTpLqQUXWQnQc+pm8QhwTWUowT5cCBmfElcsew36HxBfuz2mNoYKGBrRdZexr+stzduY/
O2MuIfY3o8rOf5XXiTzy5FU2duKf8uPjSzjzBvjtJ1CJOPp9xQMNqcLi9P1Rw2W3K9F2UzNLPKEo
jmvJTzHayYLwvWi/l+QIrp/ZoNR8YvLYtGHm15mTM4t+K5Ny2g237cspQHY0AG8MEjnP11QPbIn+
+8wsf+fvhWH0QBX7R8jFgaY8C1h7o7m10IEv8eHaIk4/YAADyaj70Jt6puYz/+fjlY0GWjkG33ps
gILsMONHNh1DqvKcutzku3gBNndDlnMWxCAeWiy04sTv/wj1wkzC5MyAqyyxqiG+5THPfc7Q93i7
alZOFOoEelzIeU+VwsWvheEhErhK9c0UCjRs8WubW2sq0Sb5ztqoHc8STi5wQ/b6eyZ4q0Q0H+iU
cj70gTejmbLSXvyt6hUL9K6/KZAbESmkq9xA5B+R98tc0QlEcpjIFwZmqrsJuLUCG2Xf0K7+rOwP
N9I5Q0pJ/TfZUbewQ3pNU/h2XIYV4ldjd8EeN9s7WEaXrddOOkL7/CagzkE/uBt5RRHWf6lYhuyR
1CZNgTyOxv7ITBY+/KhLIF286nwoqP7O/8Y3riA7vplOC1LrqJRo7WKQFcIEMTsPr2cTTpMqE6PO
lLupo3eRenofPp7ynLtODRq63pYsy/bnb5CsVi+OrnD58K0rRXdp19NlcnMmgkC6rzl9gUXOrIPY
yDrkoeaCKzJJQqlvolmWCLOC3BxN2vN/QyvJMHYOYfcIu9DQ2h9ZD4mb/hqp22iZL+FmMoKeJSGG
jNGcQtaPZKLmb8e5VvZe/Fb8lbl1EObdDW9UOHc0kyKiopY2/Pl1r6D5qqt/n/19kR3+YvA/Oavy
VR1sQNnSe9TweXJ2sQMGcbRRZRf4o8swGf6qXZH1EyOUlj7RHrPB3NN0cab9yubn4oR5ekme8meg
VBPU6+Wrjr5OxrfDqPKKobOVt4eIHwGnSo7NK8NvnJKvyb/LhAztK/O1QBaSMQeg7IkPfmJMEz6S
7os6sYCHuAoKmabPpqkRJgXCGclG4/Xb1Wqw0mNoxB9ime/4ktvEvXoDwbLBmmV6VEtJZ98QsfPL
1bFPDrnQ36Jg68Brm0GlnHbVM9KLz2Zb16p2smYwL6qPpzX8QiewD+7P634xIZPcdsbCuTVzr2ht
t6b4K/3w62Qj6SklQFGbPVn9Uzq7+acpZ4Kvf1ya3kWtjzygSt2Zv/ium37jUcWNQXnDbOtzwPJw
k5p4rS1+zOv3+xZ/nKwDbwkee2S4VrVmnEJliWk/Y8HYx1NBQqYPPNjjK7vlmct662/M09aEGKY4
CNJZ/LMnh/xEsOcJHNBzfD/497PNPeMoAfwyMaYUQnVsrr0bb8ztzoNkyxPAv+l0fWAKn7j9E/J0
H6xIpDkcpF1Op5M7AqdFwwFLnj9ZbUU0mMz3YYGTA1ll/nPUejOhBydBPlXgoFA8pVvLiVD0dXbH
aBOQvt7STCdOQnstKuZ0SK/ZS5kBggMX/OFck262jF9cl0KdXI7/ynTQh0ydm1bQAkeA34/amkoy
4b2VReExtx77VJ0yFlvehL2d5OJQa/o79GCRFvgWBHwIndIJcJ7BZu7lPTOGxitHwtE/yCsP9oEY
BQm9fMEb7BA6BcYhFvt84+gmigxUIx6HSPooBm2x6GwmHBPlJIrMaKSA5qMZycnsyjb4mm/6jPfp
iGxnIdj9P1jcCPjbhk6fzihtSYbxx6KgWM3F2mEjI3xNEaVXqpRUIR/2xP7w1m/qTJ/PkWczRNDc
ErQWUteAccK8ZeBVRg4uv5IXpWK/xGFp68xDnhU92KHIMMV7ut8/FpsV+JJDDhcGA/2CkcQOFL/k
Ss+TSAEgTmaxcAtVMClL72a4x6/vKXV3vgigePViUJPUTC0MG63JDqk/vVBAs/hXfUSWQbcqIRnV
ddP7fJp+LpjI+HGxCCzxlTTLsjdyZpMPiBLhl4HgMm9xpSLOeaz3BGuwhX51YmNUvO4Oy516Bfxe
Wym8VCJuwqyeOV4WvoR6prVrRD+AFi5DAmL35rcpEsGZDwEseSGuxhMljAp+WXFSA35rdtDun4Mj
ahlYxYwSrsnBLX34OlwNGCgp+q4wAXmKgDkXdunOj+OiXZVulYZxduYKfq6bwhssVLtBWFG/Ejvt
4YdV6Dmdjj/z5wG+dksXQX5UYAZjXYDAgpMwaobHlOS3HFSTMezvoEn/5lh44ZsuveOgck9i8R5D
+D7nFPbXquF7CBfd8yyGB7OTQ4TQQR/ugf2cpZ3wLi+IcWOs3xM0ZEzQTiTFQtVFW+JzPA6W7ggz
pFBnXjnn0r0Y7w0RbW2ktuJ06yiyRGoBTWiQAlcFQtCad/jh0f2Qdv9PEVuVCHjDP1Tx5migI+8h
x33N3I0YFPoUcp8WmuKtABYa+IQJFLRI+n6eW6pblo9NO0d9306Vm0eqUyLNITrDfMX9UMGpTSIM
R+DogbkxPWcrPB6bHcnhuaVRO4Voh0ngMa3vbyuooLhyYOjXgTfqGcPIWyPFLfg8xCK8qwQjujqc
E0Cj9R0E9DVQLPUHNaPUouU3aRuMZfayecV2JOpOEjLw55xLhV2ZncZpsVdTYxBzM+UyIgj780qk
jbL/6Yir0AHlMUbAk8jGH8WooVJ00B5mrzEu05n4CLqQ9ueDY5xufBRe6dx8YkfQjj9JdWc5/l9R
2cRw4z4DWE2zDodWz7V84PcIBYnFRQMDrzLT70FEqIrwO5U8rw0Qro/gj07tsrKPmO+7gVyo2StO
GqZZSChYiCwRWocD7nNvdC9HXWZGErFFdj79E1ZOX2BC1udUrw5MIphD2JZF9U83U8RviHydIDY2
+bwjgp4UD5Q+Bsrr8Jab8VdsRYjVA8ieL+DOj5TEMJaVgzdwJdnmJaz3w5cfUVnIYe69JwcHJbYY
1lVMR7rDDkFv+lD+GTWLtUuwpOenpEUCsgIoWfH4e3bzb6EOdtUNAWUG+Vaa2wWjyqjxsVA5YHrh
HE8s7cwLEx/0fLDy55pzawh40A9plJ/NLjKw95/aO7+DautlYO4StsaVMWrvKYHJcM11AsOPkCyx
cV9YnGOyb9dV3TRBVnLIvkiKuueFzLnp9GkrL485Hsh4iYgUtm6Di/usoLynos25e+p9Zlppx4y4
pwA8fzk/gHOnyZ5m7wUtLSplTqQ4D7fzeFHWH5h4wIM2Vo9mQFZNX7N8QUlT+RpE1xOTSbxWefDS
nqAHLbQRu94KBPb+5VlCGGwq2B/w+tS1ci83DlNgJbvj1tIT7UmNJuxsbQlDh7QrlF+Jo9XDaTzF
PEfQW6k7HUxpI2bJJmBScvtBDX0o5fVfr4tnG4yLVupZ1LcWlNYLvGReZme3ZpHtTxdI6P+DI3zo
YNsAG4vYVIN5mYZKz7u7TrI3nnlriobBB97XLYzVM/rt6C7VFp1egZmcDgESSkPatYHw3fRvXCvu
giTJDVNbVeIy+OdDBwJRSLfNnhuVTDCqqfqC6Wuahj5tber51ONfy/DWRvgFUIeOo47yH3Ax4QkW
0v2QrWPZKI0X4uA/S/wH7f4+I+158Otnd34Z/T1s/NfFtmGs/id9FL5Yy68NKSmU6xBPXv+AfL/9
PoXM0UEQLrjIY029taea50KE8J+1cke7hKWkjug4H+C/XMz8HOeJaqs5Od7fy8R2eSr8IYx7uNQM
izQeG/10Ao9vpJ0EnS2IZjjVc2GjG1W8vndD66PYwupclD1RyxLATsrlDaaDXKaBaUItM2wWQq3F
ZA5UxgPQVL61jm1b3SPP7SPOneQ+Pgws/eFwz+x0w6vGan5ZBLk/IFWfScalb8Fj5yDw0i0/GouX
e6Mt54L8MsiVm080ytWuhE+42jqQnPsv3/V663qnlBnPeHa5+qpAVj9385CH7p2cU6RtSposHChw
7oMujeTXogE27SXpXrtEd6Oip5BKfGQNzNPyliUr4OEPJhVDx6WW3xLG/L5NTzZdEc8k0wJ89cnQ
7O3+w98gApb3OmSBnt1u8reRuHTfTqbtENVyioKDwb/bZmhy09VPEazw7QQof2x5e6X0EzEGZRq0
wGZh3jhynFXYP6Ugu7Njdn9b71cTtoqZiYX5yHwDP9nwVbp9kzLd+obxkYANhYAShKmfgtA4FEmO
VwaxiZ8qmOD0Uh8v8J9AFW6/XoIUqs4yJjK6uRgl/Fw/ikuReanJL/SAGOgLCbcSN2vp7M5DYjYM
iGi7ksZFl8/A8PlGh5uJG/V47LPh2BbfiZwPnnIjHrTj9dq2Tt11rfNWPskT6rLsZFXsskNMw3Hd
UVvsZUPyaZjbAkUjWMZyKA8ceEBpRua4p3O4RvN3ybLKj6h1e3K/i0YDkWsNj0W52D+IX03EFKOF
GT8nk8gCjNflbyguoiV/F9AIuJ1wOuut99C62othgGoEFhtz8mIg1BSz/s+l6Iq6BOlecbx2ZE+o
wgD1O2SUAHcObmRAVplNN8hZHBXJ90NAxFTpHzPG+IcIbZ907l+UaJohxiNaIUb9PzZzzVFNIxlI
C5ouG+4Qj1odMc2VwGJp+swU2/FxtoOaDO6i+0AMcpyqvAjRUZhfO227RFATkMRB/9JAjj8sOIFh
3YzfHHAAS7JqFHAbnFIl1fa6Ap2c3/1HT/1cRHmV4MiBtONLdZcAZBCxhs8O975XsWw8oE9jVJO4
QbD3L1fWv1iJuj/l/TuIKmpBgATvZ4Ivtnz0CJUnWDOZ7rz1mhZUZyewVJOXNHBsIidsrSHWld47
p+eHiix0Qgxm40tl/HQBr+kPlHqD5H/uTkyW1SOMOK/GyR5FYGpyFF/BJTDLF2maZdMwmPpfyTgC
ugaelclPl6d80srVuOHDgnc78OJGQ6OJgUnfAJXM7t/1UUNCj35FEcdxae/pzz9L3SIkGYcKVYR/
G6lTM9KnLpufvuQNTkp0SPKRCixc48QYENe2gXzvkrAljaMmHonmNFKeUmtkO4q/xvgUuforwag0
P+GTemR54wZX6BJYsNB9fcnc2mBlYx1ez6+taaF4wj5i4HGz8VL9u+PSNBbAtpTLbIeXdHNHmRpK
PcEMiB5ZXaN67ndWZkCtPntiNcxeNy0J5mRG32k2F2HgXmnIJqmMsdYEKlBHuHdU/Joc8sm5RTmz
BVgoDQ8pKzzXnDN3EkKAWE7NwuxcVmdxDREHBZxaz1GThei2/cQljWFjNNrCwUgxzolXTxNWPVjT
pDPGFAf05Wg5NyAZlaDrLkamXNbPhCAq0glMzEhZ6e3Iw26LXyAIcL7i6J1j8JYPT8ed52Z7wAg1
cuK8+WpM1h7e7tJ1ulV02BFhDrrwc+j4f/Fl4UxrZKDtjSMXbvfHP5iDECAuqhOMKFyrbdq8igrd
OixHhccuW5wONxPmm5gM9QAz4oOp5PYHfSQP4oPo3DSMzWxUZ9NfM7rOGLAlJZX1qmsFB1PaHJ9p
8P4jSWIMV3MEkJQ9ex5I6k8FrTQp8tFhplTtpDDYgV57u82TEEUnFWDT56KAhAwT4rGTOv5pp8dE
wnqIen7fnn7wgXWvHWAIQzoS2QtgJP9nf3vHPOv7RJEvKPQMjiluBXI6CQitxrL7tJJiUvBI+N4L
q47t2GcIRhqKET3zizsVnhws/oXGGFLUBouRPmv6S5zwWSNSMy00mz8rAybNVeYtT0A7mjpL9B9s
gwDhEZQRwRhJE9HsE8bJaFU76UT7R71CxkL7FHqqyz6uahpfJV3p5/oAGZzo+K+My2rkDOej3GDL
X3w0ZTR90k45nlUyUT6QuK0lIEvdvmwnC7ERQMhvyjqN31CTYZwRcMEg0JfkN62/mKYtIG+gDkEb
LtFrRkx+HhVIIch97kMvv9tzit0M2NCEpU4FIHaZg1hFhWw9PBM9d/E3V2HMAIZnSCZK7GM/s6fC
p7xKZO9/RGUVFSOsvdiedPq6KWENAwLmk3mqOGk8K/+sPNKF2jU9B9YVtl2o6j5Z7SV0fSYfmudS
wta1I/WVMBpfhZFr27CMtSpyUVw0Dk4jY0T4re7XSnWwFkvVk3ZmPerwYwyDQVJZ2J0wog/CbPrE
OD1E++x00liJrc07s+R0J/RAdmVOjYBCDf+p5gFaIP71zuz/piL0X2UZTHVeSRwzNP5LfVKLprEH
XwcPbbV69ck6PEijQvN7Slc6PUQBf6B5SBY9y6nJwwhy20wQ7MZpNQlTWQG4Kf+pJmXHFYpXXQHy
KfuTvFZh2pVYUgS8q5nHIHgCRNyNecjfs0vHHtBLaARTQXNawQO0+z7b3x/sxuVw3o4s3g48CQcY
UU531Vwgh7GcndFHW/NDqd0krlyLjDQcUuKmn8IsITYSfXG4X+QTY3ZLfC3lvoOitDFcfvGO+sVu
U67Zm4V808lYs2dRSY+dL48ZBui5MFrB9pzOHkpi6sH9MrX9qmlpl+SsP7ZFqxa06W5piCtGYQf2
BFADNBXBykCP7jkXWaKkGUXqOeMnTByRibPqBk7298ebihcZmw8Al+Hdo7RsIv9dCIfp0CxTNXrU
xmARPiVgl7mi4164lsykc6oS0eCZzIZZ4+oRMp9z6y7LOAInFxIMRju9mKWm4zW9CulF3Qx8GIcu
ts/MhwPkBdpfyLPxp8NdNqQzymJwFjpK5EOzutOxkN8qX2AY1SeRf25/aP7+TfS97kL/RYVCKbwb
AXfKQnE9oXNZ627Pjxhz+P370bURMqiD7Xtm7y0zLAvu10CT2SS/XPlrBq/tp6J7yn+nbnlrGSb/
guU2E8XDMv8GFEeBfdGtSof3SijAWEMwYun8eNQ3Xp/pt4hRkYfIeUcLG+wpxXYMWzyXO0RD6wFG
uthT36jPx1BNx3k1p+BdhOI4saOOeIoMYVvEnb3qKTMCHiFr17SbrZUXNGZb3iy9zkl7r//v2ajS
qnVH5Audyhb38mZUeEKzVQeivzjFcTw3hLK9ty8zrtXFgw5zsuYrQR/wdzahIfnFDmazlaBv3o/U
JepSnIuCMSI742aI59yu4tUrp7zYRmKnpJlRxQv9lD4yL0udnmWQslpFYAekDVkqPmjU2p3JG4WZ
6coddxZT5yRlAZ8miXB3fhRbG1Ivyau7nmz+iOyezqAAiXOuyFCKxgbJvmHeWyZ6Z8wc+OALcGvr
m6Dn+q6LIQGhdrRyz9XR7NfLZh5O6Toqvy6uvM7eCn3xyRSwMXTc6xvO9eaRHpUC5SSXBkAbVg1/
hNWWjlVXfbUeex4N9LiZ2Pmi3fqfMfAbFAyFGjURE9xAuU7kgryaE84jj54Z2B6L52g2rXUdIHMq
GEVkr3RQ4QEY/3ysZAkPG+ORZZQnlpBlXAsqtH4TNLebIXcRlazVOTGOVzUG55ks9dttzHkUgS+c
D7P8G70M7sE8tRVH8HkKFg7ezu4uCgY2D/s4zy3xR6qII79UEyPp2POqi+N1cCm4MqiAsn6yjW68
SUO3DwTNQ9rtt88uqYzV4bKJJL3eo5aR1r3v+unyVJGdZPKQFO0XpgZzBOTCYMeLwNs35HGxItm2
d4VVWa6W7M7qg5Ywk/+hK3wbJarHCr+BLORDj5NyqcJJcD1uk10d+Zs9yxwEynpSzTJjktxuXmOH
IFY7bEco8nVYJsWZ4IA7AUIxNUKIsR8Pr/udY58bwwcua6d0QGCM62/uKjoEVg9txLUD0/x7SUAc
cbhyjisIzSxRCY9E6IsX+bzozuHoPTHQA1NxEUGMplvYbBxcP7C/sOIPgxecx1r64u3b4/z5BnwU
XtvW/lLbeEF3kcjxO1XKORVz/HhsEmuQpOMU6j8r1XiZ1Gihdz4CGwgIBrSrCR+zgIzMcfCEQ3Nl
hAXJIPxZBrmdVyMSHQbp6tE2oAcMT+rvdKM0/Maf2CgoIfa74Jn9EWOOJEJwZgSwt64bdXGKlAXR
f6IVEJ8BLL+LB2chIyj4d46HW7H2LlbrhuSke8CvItgRTArWDSbt5FJekC6X36xcMJvC5TbFZbj4
l99MH4wODf+ardVW3CBtuCn5d565X30x+CNtDI2m3+aIxB2aK5EVTImtfpxLMZha0chl8ZRWaeUN
boVh1lkQHxNGBymVqrXbgz+2boDk0ugPS4eeKRgFTR9GjphKwzG6fQ36uSzFOSgTlO4T/6bLQK22
F+CrQDJDiwLl3dy6zPt35uOq+ROlr6kUj5iU3tZxxJQTmfPWg15D7DVEuU7A1JlMJcX5QnH79hC2
hpeUebO/rpm2u7M0LseSGfzXa1pNIS5I0CSZEImJGcJPmwgw9UhmpJvmlCYmyCnH2H8DRTW6ZorS
amzy2OOf5yidmoaKPKoyriOSp0/qAURd7jyoeNPpBuX5X2lnzzF8AJgq2WK+jbZ+yH3gF/mnPJnL
t/lhemkbbVHSUZ6yxiHIuQllA/6vZS0fuWtGHR0LuzmHRUlorvmak01pni1x/7picOx59E5qFSeI
v9UI+2g5gKU/rPYiWHL9PxPMDRRAujcv/ztuuiEZYe9SHqLZio22AgxfDwZl432vrJI5L2vF36JL
xGCdJFU3jeHreTzm/OyrkNY8ksfJV3K40p0pXBubqMQwedi1YSFwLTp9iPLDEmJrnh6wPaGC+k1s
/OXBC+W6V3d29Dth5IP6IviNs/dRmIje9OXPwu5FFcrIXwOqhn5lMmTDx7zMoaUUUJV9/sdUCAed
QBz3eARlRE8+vgZq0XaPBzlYOZZiN+q3oOhQLMm3/rjAQxO/B6l7cuvEhrvIjDwiVGai3DmgDOWX
27vAKyDymt9GoNqSj78CBkDEyiIbIVvxzly6sB1ae4WadJGk9SZArEPzGm68x6RFxs4j4n6TWQIS
awLjV4nahd8Um+0lZfk1UD3Jq8MdWa54+pbyEo4O5fcAThJSOS1MdwQB/X7U0jf5814YpUan8o8d
lILf6oxoYxOoRp8YNXgfehvooqFXVgcJHXmn6eBY0uykFFc9M4HlepOHuSRqz3Cyh+LFbSn/Px88
PL2flhlDfrGnYYAmMWCjogSTCYKXVTRGKUUaA8bRB5dFY0q0hBv2OVbbhVnxCximxksJBMvqrwB4
Xj6rM/yUxCmo9lxa7sdI+nUHaUinTyLWdNCvpVklj/n/A5Pqw3kwTeM5t0UpI544LWThfkn55g9w
KZi6qBU3ncs1668yttTBUs11TcigbREc+GHJjWMiqyAfx0c3H9z5IeXKqbjNi9rYoCQHJGdY/m+r
9sJ6hQVVBqBbTvkZ8LjIZQFoVvwyZUujVP5ALK3IgI7YoJuGz7rks76/+dFGe6Xrqh2LdV4hpK2/
YMOhsXW7cbeyPVN8IIh087i+zP6Fmnhefax1KLo/sLTi5FvxZ43IIBCMJi4Bf03sHXuE5Rb4pVDm
PJE58yNNlGV7ea3OraIogS8djE9EC1aouGuE1weyDVevMHBq8t/FKZaCd2P3bdpQo1nnbq4O8I4z
ryn/Z6W7oxMwP8AAr+mccYlzWiRYpHKjE3wdvaDYkTFSFlWAOjo6Gl7iifjoXXJXFFJqzhuHgdpp
KxaJZUmW1cIRp6YnJb6MRBlgAgK/s/5I+eL2LokzsYDxI7edaCsOZeVyLA+zbslpd3Fu23RpXUqQ
lGvT+ucAbppwkKAn9Max+vIjw0TA2Z+BWKjrn0ItQnY84H1Nh4wgIqrrkXXQMOWe2z6kqtI0foNX
ElGPvhOwF+rHLH0pUUgnP3xXO3b30zl+FDHzoyymttg+AkAiluWVBriUkTqW5JhWG1h2UgJMueP7
1WHRh9D7cyT03vdHiHKlTZCMTB2aiPWOwfhkOMm6Q/wnEJtEhnl0RBdxGTCy1alBRoRmOjGzcs/3
6lwa0gerPYdt6FtKEykBFYLRgNIZLOwCiGBCY5kTHFrduIrc8XwSTe3cTUStlnIJ38p9lZEujNMP
h1hhYy1KRKsyuxSBD0EOjGlnKE7TBIIWjTeUd9M2I1tCwtzUFaT/FQWrYA+QOu01jBDy6XYVdX6O
CDXQB5aHW0hp8XVt/fAifEsSzQhvKRyl9KukitMAVTXgUV9KS7LfsWDzjWtqvip9/y6HXCpEkTMT
oPZWYu0hOVQKZC5o+iEj4RNOdacUtrDaxu5aBpRgFIdVGZiSjCOo0+MetFlMZOR/vOsqE/NSe8Yk
qhE+IJGiIX9Nz7iu6PTUrZ+VyMr38IaAVyZx4/uAQpa5P+9DIf+2Dclb2Lz8gsCqupQYUXzFSqrf
dpmMSr79ruN0JpF5nKbgX0/gto335i85fL5FQwH+p5pGJlVSvWUEyGO5LfjHXcT/oHjj4vCGjNBd
9AClwNLfnY8eidKDHnGTEeeQt2LRBTTGuRBz1prKcqcXFjfW/gR4HouuNdNdH2MmG/gujmT2uTyU
xBWkIQqN/4FbATQLNIf6D9lBu3zVSdxYX/6Pi8pvhF5y8vWhazw27y1Qqn86GD4qjJ+ORb/dxnbL
cPRkozJ+vRGK6qeYRLAGi0GbcsC7GH8NkKJhdE1Ch/pWR7f5sV7fYtBIztzC7SAoOVWDE/QypLZx
tB7pWMc+HrxW5zMYaCxIvhvalw6krS0SivjQiz8J6Inc3bt4qHaSlNJ9icQEy2N3T0hYt/X9Vc1c
O4pLtQDtdKa3o8MGVspopJ5db/cQEo0fI6QkVU+q6MM+Smj7MScVN99ig2fxQboBRzdO1BBcYgB9
r5wbsvXFkytxLO+Ir2ue0DpsFMg5oVqG0+O/RFxN6POw8WTlL8jub3V6LLSusI5uRC7pqYSlbQpD
R5Je4LtxNMPtHmcMk1DSRhM9+io7/8HyPEjNc0SzbnXt/beTisEDq/7BRG+lkrZRsO9PsHA3I+JT
Q9nL0LBi/UGDy+oCymbyPWUKGVgaA25pAnGotK+g0YgVfrhafx8ElJwR8In1J8ywCIJ7Ur0WpRmP
aWtLc2/9MrAiSZ/lTxap5htPlzaWNFfP+63z0X8yJAWVcvROx2StBE3v8IjNwa9Zw9eDJFmKgpd+
BofTR9eJ+is99g1EWbMyOMMYyvWCyhMxdSUfu0ql5PSCOUGEb4Eq38A0fdD3ZZlb3rpi6ROmo/ST
tNO5XecT44GK8BJvHTRpzNiDOGN580B2NWfBaJRJaCWNQtFlUbdPOQ9OA9vU1rWsMVoiz4+e6qUW
/gDPZn16jPTJaIl7LRLbWc8n+40cwcGlAyuSCZ5qJGhtH7z0k4dGKt9D9YuMBvxuv3NrktBcZlah
GTNs+fY3WOnw8OvmF2wp0KKHkWboM/6ENyt7naYAFy3z+3nzptQIb8C40F+ji2Zns30YrbgEy0pq
hVYARsLNa/D3DEMqhC0175vj/l/3xteLIyLr644L6UhL51jfrRw/QCjIwjDh7jP3cNIRVekAq/Vl
Rq4WtYu2x4egEJME+ADmmMhSd9xg/ZMbAmEC22vRqBSiJpPdprbOc0YPg41o8h7zZapaQtKDWyJm
sesBs5SMF6Qb5rtfWO3547TvSyn+k96mLYRFRWIXRlmf4hsChLxnIHBzbgYzEjNlPXiCSO6mLrHr
5InU5FNfi9OBQXl0UCkyh2yAl7vdSF7BPhFoSCjd0OeTxdnYJ+jqtn8ptYvoI1XcoJLwDqitU8KN
EJ8E/NzXGacwTltykGwpJUHK8ndxQ9fqT9uNppBfpnEm03IRFLOAqVAk+X0tSEOOJ6NJ3ZbZLOWM
lDxX8wVyPvOkXoFSu0YgcVv87fvB5EWOdNHddkzjMkUE4jM0iDBCqkv/SxGHndhmFKTfnaeK/975
CDrgexFzHVTafm2nYG7V8hY0VXAPHoknGGyD6r3e14Z+bosGX1mrsHP6fKGctbIWBsqurbNQvWm2
BnAeqA/yYouKuo7kGCzUIIAYzscgWR5HaNytAHMMIskYYuC/ZyGFo3JOMAZDBEHfL2i/sqql0s8T
SW/krMKBIJf9Ta4DLsiTOskL6E4rCObZwmITRyNXZUhKLWKKkTPm9eVUY/440VCN12g34JDvEZez
Ul5ecZhNe41NWADyFEZ2QURkUqhmjUs9vU6avRw/2ku+2BwQ764nuXCklT3s0lrb7/r0fuS18GTG
xRjkS+W5ahX1UzwZ5aLDU9WJqulNv+63QXMH3BNGxt4W3GC4CoJm0Y1mc9h27BKZg/0osmQGeFqd
NCWlZJj4H4Pm7xxc6o5vwj3CMSsk/WnM1lUkhJg7Rm4LP6qKSELNW4Aqa42ePylMwB5WXRxilI6w
zJrIaRtNr7lnsI6Ez4qJ+ZeNTJUSTb6Koq0zZ0tCIgFSNyXjSpUkSdO3jmxxN5GK68ZVpoC8SkNp
gy8oRmBdKEQUNwsKixxScm+NvmV3gGqMQk2MRH6RzD5Ml3uxHnby9pcaqIs6y3huyfT7TjEkMPTh
YlKRPkpTh2X9s6sJn4mk4BwWjOpNwnqu3lk0B/Le0fyMSYSJaKfwXCO93hmwrlcjKqGYKEIeDYiy
OCtRBuLkES6/6H6O41lOwnE5IG4NpoSDYenRrPqeejPLsKri+96gz53SKejXU1P4CcP1A8f9k/WJ
Mwqzb2ORjRJG8QRsRPeWYyxCU4qEucoOE2YwlCOr8KJDeFW5cdm2FLizzgEwkpBzU3LQbOOj5qV+
sKqxdvJZJ/4sCFPWdlLjHgRtKA2RXy+NK+Bvqoj8lYAz7G+q+x6dCPZo2VSoJl86Rx4j2tDVS5W5
3pbLiahqtAvkks4Xk+6xQVPWGFemwsqPnqdRmApo+sAIRaetOOR7C5JZL7hrXZcojXC7FKG0d9Aq
Aua4ivxP/g47AYakJtFyFVmp6T+UBk14uzaaZGk6DlYgMLY33F3ZRLDt5uM+tWuuZG8rlTfc1LWj
Bg45Tken1LBIq908xsxkaKPDbrE6L5PxNvYrt5jqUVKG8shhkjRtAyjH+/SweSOsvXaA4AjiwtVs
scgGkAKis44hcV8yGS7yU/x4THz8g1PTxmD0lrJhRHO9tm5sxQbGXC23LFQSxk3aBlH97aFtzuJR
VYtE4K+Jxwn+0wKwaf4+G7FJqQ/MMA7fN9eTPk0+tai7zXlRx9OsfPfUrgh176RcD5/HwEylmCO/
kmFsWnlQngQ/2ukxSvKyAw0ePEeC9yuCY7LrD/OTrNu1yVL+EGIAtWINUxW7/Cm6pG2lunq6ZoQQ
q0kftWPbNqGiMxOunS8IwKK1Y8+TUghWQ7z/VDgEvionGfInv1oDk+HEpHsHidPFxGd2eHsw9pfC
UmQFN6FuIt6Iu84zrGCo19xW2AW/poT/AweoqRzVgtsUAWal5f16ykGxpjr3NtKSDIIONIVhRTRR
fqEgO5t9s26GRSPkLz3bXPMqMzNl22FXW2HdJBowUMbg6HUs4S2UZ9jXzRrTrdG4V7d8c8x87c5Q
4GlPhPc5blZiaQw4fL80cXn9XIbQ473Rz+YMm9eK8Oot4j4SVB7qmdjtt54ERqhnbiZoH0S/fqaR
qWzilBM25340ABJEqXlw+x+v8xfYt5bebAtyeuCqr1VlJYTd8C69hnKPOuZ93Gdwgw6vh9lqfIzr
EnDs3s5QjKC/IhlqRgeAzOtyRV8Hd+GCT/SM89ubxCwJm0jG8h7hd8d/+msABxBGv7KE/FdFV1oE
0CjZijh7LiHkzOXNyq5zSCznEOfMe81OSUvbyWXTxDUW3etRo4Z/NylS0LBltJPnaY0ZhdQBrDMU
5BTZgHfXvhGaHQrVrMUVqT0Qs5Qs8raNIJf9vd1PAvLUMnyCMqiG2gV11VDW5hMBL7hwOq9KOKpu
Y67VlnA1GGcmV+PWDTbJuo6LJWWLK5E7gkIDc6HC/BYWbslxrunvh17C1QnOzEm5xWFQGJm7RDp4
uCJOCDAk62CAxvTgTiDH6wE1IcF+OPMf3kpekhJ2y8XqACGWid8ZQmJ9HISo4bYUHFJ9NSRRctTE
38I7rVxvEWdVjKU5Ux+zJdnYkALAduuRiwx1C2jz2eL+oBZt8/80d+fS1rof2bvcfMq1q5KwL5Y9
0DAoYeSNVv6CQDOZtc0bTvKzuczuEOOMhM/cDDjK7XJsY4KJwoG+mEEYtq8LNsyxQW2oCu+X9aql
VvlbSuN3uqRi1A7p+ty1Q03YLJwO9Yk7vd4aWiJUQQ69WHJidQvJlRqNaej7hmFN8IAAdTj6yDkc
Axep/NiUrZgoCnI5/EQTKn5CQugecKu0p0JlD2FJ6pp236EDblPEKOucCwVtPCLtY86inH1rrd7A
Es9LCWPOEwhu8hB0II+sk6+t67E2bOm8LBomRd7ag5sCg/+eRerwTHJe07Tw0W/Mt/QiHq/wxT9R
Ks5t06fr7Y5jXNUY4pBxbzVujCusL3RwZ3Cc0QrYBZHBNyyOP7w6VByJSInzG4H7RvdNlLHI7wYP
Q9gbwge191O9XUiKfwy7lvpzvS0U7fNWG2/Ii/YbEt72ozqW8WNi5jXjnoSWaQ7c6vJ/Ul2Dre50
iuvO2dIgN9shbJ8qsULuYynR7M+wuLAqWnYPID/eHA3RUigqY4WWIojJ7+zF0PQHyln27l4bARR8
yJYHc+NBHEiJejg/aDQmSV+iaK5SjFvuSl6wUz9waMyyPzRHgOiwV+11KgQhuWcarKfnLXVnN4UE
tSuQ3NSCYGSgrYdFZyNNWPdDa/4BNzbPepRFyYfPoH5Y7HgsYWcQLJkM1ftpr8UwAMLTEU1ryp6u
teMqFQ8TH+td+PKQiN9nToKorO18LDzMvhjeLMXaAYngJ76bvxASNmOUnXyp6ukXngIVaja1kNEm
EHsi5cJGE1ybVlIqC0Oh5agX4R1AiezLn5LgIEnGPZynm12pPRblbwSKeg32J8MDn5oKtRvXXkMT
uU7vN7OIbXwt2yuTR3KgadsDpz60ynUCWW6/LEZ+qC30bbUQY+lmt01gQPgVtHZWYEjtPT2azPP9
cdUe7bb3IcIiZai5kSN8A2Pb3TgkRhprYDecYBVBedb8zdVncrikpjoruFW7wPDgugz1sCgNWJae
yC8SknPueIyy6UyWSmVD9HGqCwwcKcJYrKzKW+VlK+712ak+d0Bab67oSyMq3e2ToCuoF9kzRaed
T2ufJ27YRXd18wGXFl6ML+m3IpjHrmKE0JLFm3yXeDU44PNuD17uwL2paRUbBSwOWD5w0A71rQdm
0y2qJfYoMU69CvYEVbT3a3LZRh0IA9dSz9XRw7bbhwNuQS+G6KuzSIZgqrB8pV7BliVvdq9FDuVo
9hKnTU91qqoY3bNyTyvRL+6zx9Si13L8slnqE0FCkUgTiR2izYqQiDn+qSWu+hRsQjYNFM3YDSjS
KnbD6Rwii/bU6B5vAnJ317DMRuVCn3riVQCsT/CIJ61UXEm7t9+MWf1dqmudLCYrcEJ3zaVIXmei
otHjK8n9SwwY3ztk4Br1fNPrcNl/4wTsTkR8vG5pbYr+6dIUQiGstoDDk0u/9QqU6kWZC7C2glqJ
1ROBHNBLQTzlCvdhAqyw7FVAIqh1MzVjNaJHS8eUDaG3L57qD8i0IdFtMjdt6Vqdxsj+pEs4Qwtq
KUE3DS3ob6UB8QgXkM3RWenh5JyPi0Wa1hlXaCczL7kqoAAS3n6SEbCjhbVj3CNI5A8Rq/xqZAWn
3ImcGSl+b6VII6XXPhDxaQKv+j1uuPoXab+jnceTCi8pDvtwftX8OsONo0TLwmRpV0MhRjTfT7SL
+RtnpUOaSFfSKm9UFWcQfVEhpfL+yiWgIq+K6JDTtglHgFO5EpovwGk1YGKWBlHdN0gzBufeadZt
3omKeoqTw32ZE1m9cyD7mtPPMxPYyl2rGoue7/w4TW4vOuDXZqnZBh1f3FPnRgSFypDzCk4/Tu91
SjozARn8S2SmKx67JDJzcUPTtgXdQozcpi/h9/MaIyKUNpVMlGY0BZh0fnicPzEYVRVQ8MUAJuFu
YlTLz6HeZHJVsogouj6QM6UeINQ0bqNJN+hDnLBXXNhQA1hklQQ4qj9tp0Doj64vpp2xWRLeKJO8
xXBuiJXwTmg2uM1zF7iYw6bqDQE83GzzUbBH2sPM/vHdANHi+gIxjRyYlW+P8IANMm2mzaBKV0R5
pvsYOU4SRnFfRRToUPv5FL1iTEzXRNAOI4swwV5NKajcKMQiQGaL4gtuBXU3YUYOZtGl4iIbTGNP
wjYRNpODPc3O31NyaDNrDGTmEoTMImANJZI7O/bOJcUjxpd2RTFtvIbrWEaZlDKNZ/Du22i8x08I
3DF/1afChaneMMjVTTEqK8uNRaEIrZDPifB05BiL/uBHgYCtQg04YhNynbI08ld68xTVP/eG4ve9
ZIfp7Uo7wV5XNtiAj99QBfDpphepj5dcSOK1xutYcI5Z8oyPZcpnDwLaS/P0J6HC2TF5QXeFxLQW
ZFA1eORkxJGH8opIfd7ewKrM6ywIXDql/9ziQR8N6e7yl5L5QIQss6jwxYx7Osprw0u0h+9pyROa
dOaLv1YsFBmUFUPWwZiUi8IG6P/VJS/C/TJDGP7fpv//FW4jwrWE4MlusqLnL/EaC56leT2+aY0U
sckC03Ho2QKp3ipfz8TBo0gvibmkhOdIAQkIVlmbnAip3nQJIUpjpih7ApCq4TbgX13PpPvY+SoW
+vEEUT9MHv+BYMgXHLPI6vsiGVX3pQ7+RPDWNw931C8eGpMuBHyfgLpSBLz4giBo7VISXC98PmDe
IgF6UYCETlUnn05zxfhSMbYdz1dlxQDyhnjZiGiZ5GebfTfSd+aix9iMtLS5fyZvsiTKfdOUTK1b
t6qZ0+mET9us14GwE2Ru250HlcBTAzqEuSa+PgZ4cIITOwnoFTmiq7iT07w/IbjkHl7Tc3EeR4c/
ho1+XaULFcntoV3sLqDjjn76gkhs2iy9RbaEqdjmHpHoIyZiio/83HnF/afsWsHMMSbiBdXlNDSJ
GCDrIl+je280x+gL9Yt3Mi3gOtMxeQuWFHWw6P2brIeSGtxd2LFGf6FiM2XJcXQ4hx0qpwRVmeUU
WMvaiseN8oYCMs+if23U3fP340zUPkpLu5b8fdmS2FmIXhFLomR+WxcWjvRKP7B7n8UcXYTZpAQH
S3KaAVlItaDr5Kh0SnXSQSFKOuuYkPVvhgbNvXnE6BTrP5E3LDMKtduqTg+W6xQvF7YSyJ5nh7Hf
6Yuto/fkJPMx+YguInXGmNe97BINBpicgE9G12DF+6rQgcfWRKg0O60wzDsUn/RGF/qxR/dia6C9
6qhd8+vnqlqKJ2QhIo6tJwD2xqzqQRYxaViX3Q09Y5m27fdZK8iAg3NTDsGFngai4ojF4M7exHPW
MxUlCcp+JnOJnF+23fRTZG4h8PlNn0GYpXdiz9rgBPa0zQLrTkxMgRRFtSwqMYuebd9cd/bImMzh
/lKenaVl2gQWvDCGF+2frowK2SX9Uqhg0mIOqAIJIpMS2rIEptxMkjw9I0zU27F8meNO7c0NEmNv
7bflU/JbQ/jq//C3BA6s7Qwa8QqzRTMsFFpDHjz8XA0RRD7Hp6wkVXKLKRbvYiBboDyz17LV3w98
Q9CzZDOXHfYwSRgX/mijzQZvH1AHCg8sfh9iIsKmwENTApOe+z+6LGzjbznvJs2+71bdnrYGDnrD
yy53tzTpuAeB9TJNLOIRKEl8dvRXMFWg1CrRcK/mX1NDGjUYAlMKZAmPNKe0HpbWZWReQl+VaRn0
0l34JYlDerZS2TtdbAcSWwtYXI4cMEwzhv/AtRwcbMd4x2gS1q882rerqvS4WYiL9QQk74peuyKw
Q5PwEI3xhQVkD5S+T1g63pmOUfCfJuA2vkK6v8jcaorAE92hMoxQYc19IBhtXY/VllV87ISziqDo
4kBs8PWVKBY42j/iPCOPDwr+QSybtuNOrD32RcWFUK/u1/1IHuVwZkWPNhZSmMuNFTYN3jV0Y5ly
nVo2A3w4zpKqg/DeHEMhqst422ASG6OhxFMhPJdIG6ylDR4eMyY258A0uXXAjUbt5p1tYt4e1OVS
UvFwdsBnJpI3cW1oiBzI+MH+g8dsgtrIN9F8FpN7uu2G978QARvyEK4mzI2K/56rZRA8U/FD6CY9
1DvIpuUDc3HNCyi5ycg+ehRbrYubt0zO3q6b30SjjvfJe35FS9GNW+m+kySR+0eUe7cvZrXlddJq
/k6zCVRCeNvH+Yx5GrlTBO4RBz+ONQlZ4dQU4YM2K6L8qScP6surgQ8XEDGvzx0J1D3kJcgcT5Vo
7Iltc7O4sJlLF2LDimdifOZHdFsIsUWd3SZw9qBTYyaYQY58pSvoDOF0xYArMVbqohFM6Pord/V6
TDvz/t2dieonnUnSJw7O84feIaoWkyFRezpKtCRNVVuAJ0OVBZ8jfO5wcHAnp+tyKEyog93XPMDK
7t0j+sQRMkGlk7vrqR6ZRkV5WmPihun0KiHV0EBP5ksVIZX3tF3h+nwu1/B+BZtokau7YD4MsUef
r4l7HaYsGNXlELdVb3ZZMPnMGcNQeLi7Jq21WnsK+3zqc3n8RnvVu5xGGBsN41WxO+dXCv6xIK8i
LcJ0gDKVp8Kr0sBaIalzKZ7ROaA8OILRgWYXfFFlxWBX3VmjbY0Yk1jGKXtLePDUh4BgnPbmlcj6
WThvNQ59+o5Gel3uUcRNBTYc6ey5yzSV5uJRo1TTWB0qEsu0Frc/3sxHnuhwjA5jOOvVP89+ibMT
kv79Hb4XQdpN7/KZBMAdr+f8mK3BbXvC2rU7HTUD9eypd+asZ6yxu1EvISCypnBJwq9GENnS9joJ
kyBUsM1qivGV82JMJKKqmNS6QgnQC75EeFuirK/5BJ79raJD/2C848hP3QW/+och9ZX8cpShTMTK
VmGpcHfGQONmrfvvtmE56ZjB4oB1RZwhmFTf34TS1W0JFbG5LAMwumPPvNE+Venkpu/flUcrP6i6
BRmbeyzT1UJnThFWL5wyQmORTmH2C1ivcfWMCG6roLnRXxemUniwu8ZZZW79lUTJrJjxSv8KQV4u
EFNHbNydY/W4YmSwegz1tt7yHYxR7YVKiQEZ0QXcA5TB31YMhX7pJnYJI2lAI0TevlqTYnSpadGL
jvoGuun9yLZ0htvgl+YrIyAR8UdVb6ryPQnjNVRuDNo9Zazt5Lys7bFQExV8b8LELvFo0Crz79wD
87StU2POiClqbDAIgMRZ31eI0Cj+ElObfVel6rrI1YGYFoRDqUO1sUpdVGdwlsns2U3ddE5mLe0L
Thvb8qroJGfetLt9jex+2uXRa5pHswQyP2f3flkkR2txvVtAiUK1Kaa9P9G+R3noSq3m9rNXR3O/
jJyiIhm9mZh1tZxw0Npxea234JzRXb0/btqjEOLMtk6NJ8uPBqD2wtdmUIDRnYXzPoOwCz+D4/Hu
NMveBhWAmdnsBSJty4bS+v5d6Oah7rpKzROfSpNJ6wkMx/enpLesQ6hULgk6ufeBVqOGnPb6XYmT
CTXlMWNQf9J91jEi2laMDV3EoP0YnGhDrcyj+OpHLmViiUeWSbtnYrczp9nZHruOsTHqg8DIV6QE
4V8M1iTjQjArju9J/xSKaji0gD86VIWgiu0kqscsQqqAdHxvU90exXHtWN2HI6ex0H8ewsE6tk5x
4u0T1oLf6EATDWRB/gwMDJHqTO/Q74GiFPSpV5alj1d5HhQjNhx6iRxIf5dHffg9vVN/VDxMTSum
YLzQA9La36YIrh7z8UHgczW/uptjFf4DA65ru+9DyQEpGSN7IRjWj7Ax3OY2ZWd2ILqyzRQFaAtQ
xLfVDA2dll42eOzJlHhLN68al++j7TkJkY190ZR+YhXQoQ35raJBA0e/qKUxATMcTlU3omNfZ7MT
UpTeNlq3PrgfMbxvkfkvWC2Q8Dn2ZnzXMmOID9Yyr72sjenz1arQXyFBk6xT3Vp0dc5w0AGaXHi0
2Zu6jFto6cMiQeZC3CQrM08zVK2X/bZNMYuAVhnuyh2BhlZTjFleoUOnZt/ND9ZA1GdWe8k6aHwi
+vhWk9qTzu6Qztu34AKrQDaBMWUase8uQB/p3aq3pYWgA6FYeCtUErXmOCHS1g/8i2TS6UM1FYgk
zkvlFacP69ECCjqtG74mBHq6MAZQ5BIVmHUIdZHUw5yupitaguFLwJYxSvul8Uvu2evbO3Bvxrs9
xFJyLeHNMOQJPDKvahMRgWQQ2a1OI73eLKPd9GzF2Rcq3PfKnLfFUUjB/T8NK46gi20ffOv6cqF3
1Mxniks0yciyBoZ66cTeNruBWVDRubt79etFpONl2AP1zY5c6I4YniYOym9+H6HCLCSLl3nvPDJ3
uNI2YDP+G+LJBaCneA1KdSu8eXUc1+u3vEJlnTl1j1egZCdO6MeNfUfP/FIs/gPC9QxyiQP05Sqs
QLcqkuUhqTdwlYxPBgQwjid8EEjGLPauaxJ4lidAfT1CMyVHVI3fFlwpjMW7J9iQMOdrL/PDLzNk
TrzR2ieRQuogX84630exYKL3Da7PyEva2Y5KSipHocjIJY0rSFw/dZ65q4Bm/fOdoys7zBKXXlMc
nUJ916mqkrW2WOCEXGfn3zbowkpIB/xPAwuolEh7IpFs2grKyqu7S3UEA46vYqTIiRaJBqZW37dB
5ZeBrEFbHlDJP6H22/fAKKKcSQ+1d6LOpzRFnj5Ukq5q+oY5mAkAR7THCMBzWyPCraxxCDWIbITH
Qu/GPmgRntg7xocJmo1nbb27feFWt07yMEbol4pBVvr13P3WTAt3esnREAUUdE4Qo3BaMXqfqF3Z
TpoEwc4l40TNd7n1klGxyS4XrZcOPOPkr+4F6E00QYKNeThsh3w6q41HWMuuGGFbg+hBENhVLl8B
T9wvHrL2xCxu1vz/3R0NzNUSHNSstux0kJGmIXxjDHu5jjlxPESW+kViYA3qz3Y/kdQtAxCb6E9l
NdcV5YlGT5VhIZeOsFhZXXwVYPdrA2kdPJOeo1oWNz8jKb6Bf8ET1eSYN6/2SuS68/O30L6cF+LS
bAWlpygi9rt11f4OnnCQC3MeXVvZvvo4R62uzgzogUfI45jSpBWHCvh/RUCG8UJr8UoKXYswHpRf
5UZAJTQFBAdz4mOL3XCu4m0d9vp9ZdDiPMoexHyQcYHiEJHOM5oC91oIixa9NIXD+Soj/9VAKpJs
KrhKBrfDd1Nb5tCMEXurWyr/B8PZ4gR/Dow5dh9M6N/ljRQj+qfAmA1QhBYzbgE82IvHAI3K7BXp
KcZtk90M5dMQ/iW9QHtFM/sTmGGajMHpRpmORhKb7QtpeGjZd78MRU14t882fVZDuvllr+jLjxyr
rp/9LG7e7vhd9juVpyWphtOX5T19GB0odleCwzuXmhMC3P4/+bs0PyBESjT39V5PKr1rB0v8yier
WityUAqO9bypsT/NfiTEQksNaSAzAXUWFpSDSN6NLiJaptibc3ZnnHZjsl7TfVPrGd98PRKhxzKQ
EMUvPjyUyn/gxaj8keRKk0mno+sp9PMMUMqauIIzlYuYd3tyUZMbbsxrD3KI7ZknzFGSEf+gmiLv
BgKU3Ms4FV8Hh5y+w3oEdmlr7vk/VEQ4vG+RcK5/gcjWGbkN4LJDEYSlk088OA+ujPBimXDFJ9QE
K+rTptdlTsb+tTsRf/sWK3dHgmC5ohxKHR08VLciKBXhRz3cSkYDvXRY1MRvP3dkJiy8ZfEEDiWK
Zeg1JxytnIu3vwpnz/QPpfrOF9yh2P74JXOhQpvLdqDq0FptHJdZD76DRGoap7iUBBHeb8o5e/af
xPPCT57zfu0MvzgZ9tHBz2hwf0YrakfOZzqCXUX16rnKeww9f3K8YDF9wVvZDzzg8O4zrGDbzdg8
y1SZDmHG8yG96az6sLuM9BcvhP1xHVIHlvy1ikuLtxwjvXnRwgnX1D7KBiaTGI+yrfPqcIA0LqoZ
k97cQM5/QRNw0vgsHDFKTBQ+dEPrN3lcsTfiS+7OZbiBzpkl4PgIvMink+Bh6PjlQvAgqIO7YHGw
cHwFiN3juZXJARR1vFyj98UQeHlvfmObN/x2sHQ1JshwWQsG6G0hwn/SchC1Ksz7lniaNzWmzOSn
Aesabjj00zcrzHnoAsFqVg/zNFRxUaV0Jn5HgeVnhXOYr2CKpPmCWGhP1CdXfkw+Lf9fvNoNyKUv
jsVNOZoWbo4QTzoS0ew+AW/mUSAZIB5bHDAJvpjHXO60jUAXFHVe2CTW4PdqcMNt2S6W++vbTJ8L
VZrJ2/nlPOSmolXk6EU0CS09Yx09TlWcfNVGRXayoubNpNWENoq2MsBbD8x2Y/fEUsOykakHkNeY
9t+Fg6DEYJ1Zibuc3NSBeLPyGLfUKwRBIEykz5CZJ++Q/wRFZiw5C2hPNQ0fNZTGz0MOPO9qfTIB
WiFTPIU3a76KS5bdCIABrgG80eG6Bv1tg/0XsfKr1oBN0SntCqjFcbNMx9VBDJ4/gGbP+9yyw/FR
Zm6yKyjdXbBbKw+UI4v8bUnO2JDZ1yx+3fNj259/VSyfJlWqSLtllK/dxrMrhagZcNdZbIR2bLMo
LcjWrZik6pyLFeGWFHKBxeVDNlvyEBJgn8o2S+pGiWh86g99RbY5rUwAuSlArq3xk4HbncBg3M2x
UmkrKn/XF3ynyRKD6HYDOa7RNfMMBPNhez2/nv6bv0a5AlyOCsF9Chj6uxRmk9XW3H/YXQsx0RTK
IJObpMHzIN0DKx54JIYxAzi8pKMv2mz9eU7y03aBwXCe/+0QoESB6nGd4zNdggVOrgUuojNFFO7e
5mR6sXncNw+Wn1CmWjJ+KsBJsnoZer5WXDgVTR3EQm8X2aIJVMbEQk5uNB1HEzFTh8B+WBa5lLsW
2cOy5hoWBaqGEEo5jK5miutSb6MCvnLkHVa+KwfD5WOklyNfCBMSh7GL6x05q154/fdI7fnlhFAn
0nnGMDtAjtIzOyNHDXXSDNh/bCmcylHbNLSqQnO0LT1jMlgll97XhyZ7LXkuKFbPTHOqmm/bZ1JE
5EBA9PQd/7EgP/udAHxqpZMTg6vFSK1nelvivYshCyl+kQdOM7tLDqPDeXjCjTbYLCf7xdft+lYK
I7L3IDDoe60Xh/IrwscQWCLVfv86Z+hNX/2MVPP4McRdIcFmQjofw/HMzXsXpMJJKfRxtkt7z9Zr
pDL4X643Q8wcst5hmAtjmBI/TchWb/6mBFtWHVWVw2EVyiOpwRwKgFECqlG0of8mxJXJvPRzkito
PcLhwq/RVWIEH1GgVEWVio0ZeDfZ84JqLHEQVcRhsfX8o4D2vbY59aUpc4b51JztF4cNtAE2I0EK
jM9P4EW871ioWiX9vwfd3oNQEKYWAcCCyN+6/a/x1v5GXXjCik0IN8eott8PY4k5pJNfY90rtEIW
IPqHtXhV0U+70cY4ZAy9BxEG4bAhqDGAL3l7uW13wyos07VZ45hoqFRFFDayXrKUfSvMa0eHgGWX
Ucuc+83k5LdhZKrHptCdBRycUb1KQZoMAELdSizKzW6rSDktpuYQ2WOHrNeBDtd44g4rGPLuIG6j
NGy3LNWIEoMzejw/LoGECW+fLqQysFLjMlsoefgnZAiufvbowcredstr7rGYXPWBynw+wy/7MS08
sX189qkEfvAWZQZOpKkol07ksLvHb9OuVgJ8vUGMTOHP62+293WD6bFCbYTWdX3ulmhyaPfg1UvC
NOeF7npmT5bK1QVbucubLzDJ2IcWbh6gG0NOBezGAR2v9wcyk9xw+HeerG4k8pMtZTLlfl2rRVYh
EXmIJnXVBhqxMvz+v3sV5yEhtmIJwahrjxcM6TIh8ZKIYaZVvkk2yoAL7AuegRNQDjOsxX9fGcEy
ukBGLbh8XlvioA/FcYGQ3oY2gxAr75gpFfaCV2KZOOEDUUi83HjjZqKGJ8GIpa4hPgJrbc+AGVwy
SgG01RdIvlkrybglV/t/uASv6U+GormLYL9GEFRwbmtzszpPIMSRSMf/XN2+1dq0HdIbLAyk0EbE
BrvywEzpkwxLkDr35ghKVewkiQJVNFYjd1dMA1baH16q0V2OZcwrDdyyuL0fN/ZPrs/o5aKC4XgI
8Z6UrBlU75rQ2WhDyt/Q+ovSVn8cEouxbEJoCPYojee3U5CN6U5Ok4zBDkn1uQp8c/7dtRUt7KFO
QoYg91DBUXS2ObBLz1voqDpQ4fqglHIJhj/Q+Jrc4ilRN1S7Qg9imbl0uwWLnJ4wSu5FJ1ie8ggd
OjcX0T25S5NGvZLe8Z73Vy65k/GCFpFLsnv05JrZwP8+TFwmFdMJGUVKJrlLqWM5KM/HdrtboxUo
DcVCJH7n/9AlDExDcIO7rTcr7gOWRW4MKytGXevMiJD2Eh0cVqjca90ui8QAAa8u7ys7D3DpQ0zZ
UAiBNR73DaO9n2wLCSsVI/m5PSeQHO/BZ5+zda7p6gJndNShAk7FWcOUuqIMuI9kQmNBdVdGgiU5
DJRYab/mbXrYCu4RKtJnzPNtUYNORPXm/6duEXW5OsFZ0exB84C/BRmgP9guYYZE0KYgC1TllyEU
CAsl7uqctqPKfnCOj1jwdFscKxrij4IwVvPJnj4yK0RvvffKJISaH56qu+cxB0liFI/KX9h6qptL
omKFMTlLsvtdwu0HX8JkJnxUUYq19fO1raOIltg4SAc/mh7lAU8c5qMDZYp1aKbArrBnpbmsdLUI
0FcCcUYQb904hQk9IJn2WLYZkSAQo6ql3yeWXarkd6UsBu44f3skGwV23SBj8ZiC3ob4oMs3Fhft
5krU8cejgdu63iUUwzP4AMk5OXoLTHMbHwylj6jhR2nTEqh6Ky3X9r7iG+bzSRdjlxDUaBMkc3eU
veBizJ9PsFEXTzUvYalkVaSYCCoEsbcg8mIIKlwiBqSDehdkDEV0EBrMjfndo/mSMRK9CAHoPYyW
eVjyMLJScfTUCOvEDAWCUZ+GmlBkx5AcWn6lNqbN3HNDCsxXVe/tWa32AUOfWAmjgJTRY4LCmX/i
9ZvgacLM2VJn3gozSD/26Vql3i44hnL0YdBg8nUI7pQ9aPWjvXtlX2RsdVaWjB57DosYWRhaVhfC
0o32QqEziF+v/D+IEyK1hXQOWEP1HkmNNfQXrWxrlFkcpHzn017tDMdse5UJSAYu3/eJnlqGp2Ag
pLrOxQI2H24KHCHPvE6OmlVSh6AaWobJFda4zTKHdUlz/09jlSViPXEUrHQj27UfLR/0gf9Dq8C0
xMvgCkjxtQ0H0U1ae031FvVY4eFDOf2J+q803qa5DPtsbmlh75fXOL7QZceTUfLvrfD8G3RY0GIp
nyJVylx0KFyGZMCo91K8Psqi9QPRhyN648xOdSLgcJmdgygyeecRymR1pijIbyQzy0KdGHpCFU8r
6VbIuGEXBtciJZx23HtFZRh8dB+M+7lcHvqMeG+1jAs5edirdilT2Ct+MUNDpBP7+nM45a2C69ON
8daLOG6To3jEHydIOq2KVC466KOusdUtruxMfSrpawNcgEkGTQqsAD/Qn5q9wMfycxlw1Ikn7Pgc
YXCRJOUbO0RTCtwevoe8G0W8+8lTT0IGhwtHG0p8VYnM+CQbikgZFjL6fBH4bGHwVR92dak3ybZc
XVZHPvbp4OGcJxsdDOGQ2zru1ndD+F+M+7io9K9drRysj8Qo1WkRAKjDv9Mt6XM1oq+ynSqptP2q
Sk/iWeC7DYyQPs0aJOFtbc7wHFejgOnye7WTMzjsiEYhuBOSnW6JnoRp3nwQGXJKBGYo9bqzFXt6
GDJti8n57NY4AeccCvDB4JORx0ycVBcD9qtVzFLGhAsQymNayHoVrlFxtjQy1rb6rT5SLiklYcHg
0dQqKPhdk54Rh8a1Dp97cym3z6fCgSxfAtIkOV2TFpD4KHd6eUqB1PuHvHxdB2A9ANer4f9knjru
Il3OPoFZWMPFsWkZn6CHQOGv/vRJqcj7vo8g+1Twnl7sapC0Mq2sQEpz6x9NTatZljfs0kc7Nq1j
WjVt02K8aT2Rn/WZMz7resrQu3JMOWkMZ4aKschtU+xoIuWr1C/wTHR/VzFl+gLTnl7Y9TudDmjp
HP6uv1pVS/5xszuHMRDAS0gsBJcfI6cEOLZ7+Z3UPH6Pay8CVruFUbKCARVJHWmPxVbIBSezGvYP
6jKV9NIHEsbhjvO30HouXpvSacCWCisuDALe8whEt9i33DpubRd2nu6Qw+dylJ1KYjqotdHHzOJU
t0JPO/F4hL2cSoqVhXjGORbBcQFEX4AReFEXgrtNnMjcZrB/YEQHpsVhQATiLrc7yeDABK9qpsQD
6L/yC86Ng7aFJM7ZaQAIKhP19cLfavllzHngi6tTRmUKw2f7eAcLs+m20OcJZoEsOmnAGzzLp0p3
QeCLnNgJzh25nJh9LIa6Arvg551jjecvy877jkWLAbU0PrPvT36XXfXiYpTi4JaZE7Q9BJLfELzd
YNv/tmF82N8jRmat804bZFzcOxefqScauAfJDgAQrhViuKx6sjLFc2a5ditmxd1I4ee0kxFDdFdJ
nDXp2uWMtFiGkrwaeZ4jTcdyvdYWRoK5zqXqHKeyhMvkNsNlsEEjnwS/5oWZ5RjEigZLYqT8BdCM
thAwvZekA5H6t4Xw7Tilhpb4e1X9LceYa3RanAo4kWqSVEKfal6rJzCnTLcqUjSURlM/XZzQZ++V
jIrFX/kP87PO40eog4u2Ha+Fw582wZz7KtCFgfk/Lm+u2gAlZ/DytpG7nkt4oIngrs/WrUXlhEH4
PZ+lQjqeDQCX2tyIMxvJR9D3Wd2spKHmej94o35YCVNgLWr+ArH2vaK9HEWT8RcGNuB/SDoV2c2B
giQkL0Uv5bKko2I55ZftOEDOssST792nfHOpq0dWjvRwM1dqElRRfh44HIOfwPbXzPLFtoOp94hI
FN+SLtJQ44wGj8/Br2ZOgkLD246XYjIHUXHpSPKJIxLXO3fukTepDMDUETZ63G61dn1OYmnypwOj
ztBT4/kyoDJY65ciyt6HOR+x5DAR3cqca0xAn8BCudq7Is0aM3GkXtW077HVJ6tT7Z0Yq3dgVh1/
4pQ36gNczssPP1JW+a3c/qFJ08wKKz5xcq8EbEX8/3EeDYFgnPD4K2ol/SLcSEP3/Sa8+ZLYXQ5n
FivIrMRqwRNF1IyVPqqsRAc55bunCGSahRXwEAu7eTrhIdV3TfAuN/FI7WydAz7TJKKROwoWZyxT
Y2yNPE0iTbvMdT8mqDKyO4WGMf691a3C96yn/b7OiSFJmHYXa0jQXVe7JXkiZGDut7NvgU2pvSKl
zPKzdfFUV5dmZnC75fdHCkapCiAX1wsvRGwBY2/92nnggDxDEQAdPoLm71jbglZwxDVFco60uOxm
4dbFxfsqcQeERcCI0+vlDJU018kbfrWkr4vr33ucaNQ0Fe/JNEB0w14Wk6VZq69m57Gt2xppcnPc
nmnnf7kG/P8tUEVlOW5w5o8QzH9H4sIBv0XlYIX2xWQjYLk6Z6ymqHVZ8xQdJ0RhHQrJlEMlExCh
dECHFVq8TI0WIyS6q7ewG+nmbRzQ4Ij+MvKBAopQ7AhxqqmSxSNxgvA9XfnPCqPTHSwPVBWcyjkJ
U8TA1Py6AZXvcMQSFZ0e34g6gWsLFymJ6R8VmtzU9VagnW4YqxcugJbusnm6smL/xqUZmrKZz1b/
do3AGdpwGnelUfBw0uuWkDZVYZIRtQsRI218Lp+NKwbLgJEEOMLRw7vfWO09PlXBGVrRuACW9COZ
yZclqLae5tPyDe7fRRWSUeUl+VUQ/T9XDvrbv/hytZfcuiICrtIDJ3H8gWRUSeTs/mYoCFasb1t6
Ej0Dx8esVayOkO2TdNFBTQDuH9wan0Lmq7ZEK0SRd+jzSl1dmMj9W0TiRtg+gMf98pjg5wT9pkjJ
vxEdS43BI31bhoA3aEEBjlhghZj1PgDpAW2gtpwt+TewUSDv3Q/c6dK1+tCqgoWm0ihFD+f9P/sv
KJfU/0mxyeuh9ESzZjd9FHSI/k2/3F17lUw4DE7pDhQn3NfkUuAgyn89zzPj47XInCv/gHdnDkKL
tVFjD4MMI9HymvcSb5nCVw62bqNVC3ZvqIOCW5yfFinUjxik6Qgd1Yzh8GsegUJtR+ievB9owX7a
ZJH2JRlllcw+wguR+fL3K1X2BvUhBcNjCAIH34jGkfJHHCPvS8EU89RCmn324nY92CNXmFQwe6if
tNZVQcN9Blsa23LPQNJqXMS1y5O6hQ8QbOPqczFh3Wu9DdltgKjidaPJdEIhbySlitxA5lqaxpbx
ULyVWtSoDi79tYJPT5faIIrRl51QKaRyFOJtVn5+vmF4kN7FBWv17BqNfw+snbNhlSY7ze0tqi2r
5ST9rB/LkNxHQPORuPUG6pLsoE19HrV4lb5k0nLBAD+NpPtel41c+SpY6g3mMdgwmBd6dYXyypwJ
K/XCcukbMtVNlHedvwpcD5M5fnq/120F5SWAuze3a7RSZhlRigDWWubAigq6qt4jawFIEpi5Ld0H
I8ogrW4ORlNUUkRtzkJfF5cCW13ExJMmLdYax8Y7TVCNSJ4BcS3OkcZwZG2MudeHeRr4R85nxiEp
Xj79yf2gpTf/TGA7Fnba2QQNANRd9u0gOb9IxZukCPlQCwZfqT3tNtFxwPipxlXYjI4uJoc0eGTl
tmll4oL5mkJM1/yZt8b546QgkKHiIUxIAhHGMHaIkWh8oXLNYb3dqgQtxxNbFBf4+40/ilYQA81X
Pcbs3cCmu3vMa4IZ8Ua5kdn7MawXTyfXCUNi220cQFbXPA47UKWpBlH5ZRJig3WODOOYRpk3FF1X
sZepw5Kvigyn4FrOvpB0KreyKE8kfkVGv7tK3YiQehuuOzStsfM21JMsjKugrA35uVVr6CUtIRAf
l+3yybhoyp7UlVp4im2QxtoEnWZZ8JAjHc2QnaMNynnCbpMKkOGeO3KzvMWN+cO7EApubJuwu9KG
4KKtyd0VwwBS+bD6sJTACUlEpIAXbKBsci9Zm0G70sEBKvG2Jh9neC28ZWGP9KWEDM9cgYb9+ZvF
J9ScnfzAZMIOG8wAEYGAL7yy6SHNngbgdSt+1IdEgFEXzQTbHVfuIh4BKZLsoLc0qdEsiM6gyRoW
vn2P1PAZlK9qxx7eyXvFTeVyLDG1wGAxh14OmmmShdBAi2Vqj8yr58ThpaGkAcFE/vllMmV9jWU/
0W48ng2FD9jSdj7sfN0YmwDTz3wvCuDfYKWH9Cc3NaOzxyRd+1EOwbQ9Yd1eFA+uoMD4O1cDsR99
rlbrC+XaXUvnHu4phdqB4n7nUKr1QU4qXZByf44l8wpBZNRQtn4R6n0abaXCLL5KPhfy1yS7pg9j
0MZWgXg6OcR/eteW4+HNT5/9ZUGbSDRqTBRlpyU6p4XnqVT7bTIIWWYK8X9/j+kialKDL98jTQhu
5AbUBD9XMQzzkcAYCqsDwMgiXSx3VBC2fWIewJKxjRP0BjdEksjz0GP/jpFsWiVwYsesdwef3WkU
XgzYlLCIzM5aSN1mpv87WvBU9t1KJ6986pGEMTPkwJ88sfOD2Nd9V26/9IQI/jhT/AV/t1/Aa12U
6STWGld1oZ5zu0ebCnDyRCq6N3AiYVpw/l/sKBUJYtHLd7tGSv/Gk0NVc1goc1qYJEv7aZHlYCM6
XaI2F5BLAZWw3lI9idXu29oFc4iH03xpmptbfxj1s9Yfw+QBRpD7CcdRA1Rk7nO4wjXHrDqJSQO+
ZPextpxMP1NrnUPZC7129Ll3pcdMIIx1AZuverrH8zn7eQp6fPj+6Ht4aVDrd7MBYWtx0f5I37NB
HAmSkVAL+/JFX7BhxdVcwoRZlacP7i1NL943xhnddlp1OdCrLE7S6codL+hkgtHmLK10q1dbiyTS
nO8qT+rnB1JzhyO6BWN/5rmKJC/W3wamZEKZ0vd+0VSqGhlvsSuJaEO+brlVORLa9LFMEwPIsjmm
Sdu1Njs57AbpyZGPznPVLQv9xibEshqFN/beyEipikJkebkXyIIfywCFABapZ+uLw51JwtHcEvVm
+qobgUZCaOasXptVlGtujHega/0wUgPq5gkLxy3H6mv+R5+P/zRCq/eA7Adc6hmj7G0mRhPJxoHD
yCslV96EBX4Jf5hUaoEMliTWYzJe4d6+EZLL3DT5D8cTUBPKKVZeJajoJCpnnFk5/pGZyl8bfDu0
rluB2Hd4KgQSUzOd7ExuT7NZnGzecNAcWIc41T4+lyqCHo3PWXcRmd/8fNNLqS4dni6o/maA0Cg7
mKeGi8Qc7wzN7O6sbTFIsuC3V87jPsV6IFgNRTt7TyZ6ej7er0eJCidGHJYC52NcnwWCXX7nwu6/
jBZq7e7Viei+Ys/+hD6cDkGQYpXa4oe0/JhKZhqb33YUJX0O0vniS51ZV2VFUow1vn07UmmoGtqf
j/16J3lLLJtIXXr37EYn1NCLHPZRl1O5gSE4r2ctwvP1ErQkUCuE4KM4HnHicMvCWrmObT/mhdRq
S/O4Y+bESGAHymqP9iGSUeAoWE0eRl4CXC42YR2P8z04ePPoJCsiJztO1SJ2+ZaGdZxQNcBLcCxv
WCCu1Db4xttLTTx/Ul4LzgQ0nEp17QWj7gF42CtBhH8eocXDlgL2DDER9BFvMStdjPuWWi4TjjCp
fLqvlnTJ9FXC/D9QNjj1mXOsHQguuZMJSlqN52pPydQzUwOMJcrG+bnUAC8ykFF918/rHLru5HF1
HZ8MEz03Kqp/AXquO62rjb7H9mKIYVkpdeQFPmfJ8YME6wiMYqSkdoAYz1M2A4CZlj/xVzXBTUV9
wbZ/2Z5pdGaY2Lx1O1QowlFoDdRMB8Fk3E1fUF8Ki69QDt+WcHkJJIUmvXbkDb5srJ/hEgaXDcNK
bN+PItle5akGSHLoBuot+ocl+n4nWxykVzVKy68oELjYPUMl9U/2XRoow10NLjgtzP2FCKQE2ful
whMLhhsOMJx0Qmcz6ycJcFk6GUiGOVT0m1PrfGzKB1+Oz2gk0C3LD4XtP6sx2Xhg2D3nsDFlPfG1
ttJq/dCdZZvbZwKzsfdmzgmg9bXltzqab2qg8y5EFR4fCMWz3PIe/TL6Yhs9RRLQQ/kCCWBySLnz
0tiMwVxULpyvFNfw4MoqwylTlTInZJlCQ+rAJ0DX6TJT4rpsedhGjPYgfYYEuKd4lxwlQcmD/ky5
vtlQ94P6s0jleztBC+RdpI50PgwvkDl4BwMVaN3TV6+O2cwT2/x8rtrw3tx5sTHbPj3eJQIdK1T3
CPruDeC2EjviXjKVJQBYqq8YktQZf7VF001zalPl4OovB6g1OkZG1cAHjohGbKgLjTVmri2ekNtU
nSd6m3o8Q7WK5HAXwhNrlZAECNsKll/XRjPjw4oLwra1zjtshe4nxoKi2qv6FemWT+DoqPCNVTdI
LOK6ICaZtFlqy/+Sk1wqdtew4qQ9llEGKongvwJqMAIPV92k37BFrVzA6egHLALMXf30ix8f4Bpw
Qk+IpD4AZA0azwGD0R5O7Y801OrSLvubbK3nRfJmerQxqIxIcKx/fTsITrofTUy5SRXtUcbS4Tr2
0weVd5kpFIScCLBJVL2t8JNKFJ4ZK/nOKc/vmJNdh4lW1TQSdakMej57KpGlkEM79sOaIdUI4Ok2
BNBaGPkLiOY34zwqwsZnohUvn+XzT4hs6MUV5hVwE4+L2wSx2iy5XGZhjnKpVmrxs3L/kxoIYqU8
v2sA7G2l1t95Kxoz6Y9iuitbxMSM/YK5iRr6eQzERpNDX6o3a00Fn3ehR2CbMTZEt4nYLKxFBefZ
A5C+oqrc0sUYp/EMx1DwAR3TSumT2uH2Fu0lsFR4n+a6KoaVqvIQBm3l86LrF/jaGRwiSQlCZjR6
rtFLGfRDheGGrdT4KRF300cQw3a7I4TQKu7OGobP4WYgSe4bU+vYuk61AwbBw2rxw9A9cRflbDV2
F/HbfT8YuQ0CLm7vzKIFfVrahKqK4oaBNMVEbUsbkVBDn0uH5YpIQoMivzzl3jFqUl6JIK5XAESC
FaGq2uQRtLD1/JeibjYmB44IwvkKoEmytyZzq3f4XQQAcHmzEycIkqH1S6g8FGaA4YSaoHjwOOsR
Ld5TYlSPeYx0SF/Nt4JszIF3sZAZQhfMqOItVj31kwBE1JMG59fuL9ahYpbVGBOAdwnuYl+e6IM+
jVGeF517QKTK5S1wd4L3tSkhagSeRsCespGt0C7Ke9b1ND2vxZO9DgVzaMFtvCvNdfdSfdUJ/qQt
Bmu9Fi4QDv/y3DSV7bSsPoiUMZTGxX3t24/hPIMbRP/R41TnA9XoUKF1y8tpY7hxVZ7Y5BX05A9r
eqOz9jfAnsFpqnnU4/fGELa0iqIg8I21LbjsOOZY9kT3lNnn/KVMzH/0T62gcXS6EueOcIj9nlIl
2dxm6zGSUgvuyMc9rBkcDM0aI5KyTbSvBiJmR7ol3A6Rzta+tjqkkF5WQrOnHFoIvPFcG98n/dwM
hxrjDp+ECkPvS0EljX5UUTSn3og40kzmD7n/Rsjb0EkTQXjkb+KVuDzQZlpPHx2nUP69zwoBFk5r
zvcxeq5zmkrQ0pZqOtwajxCaOCFactuGl9YqzE1QBlgmmSWp77XEmPjqHPTlv7Ht8CKqp4752abT
SnrJnW2njhUpI2WCts9UVqqzy71ZIq3oW9nIk5ouXxbJfLjh0lU/QuOoNeL+VkAtJEzS+rqdgs/h
+R+3vtrNKR3UrC21BFxC34y1z29MsBS1vgIMCB0UW9CgZnL4Vfx08V1ajdkQJ7DFMED61QwXRNOC
cK3mBLY/9pM18HOM0IGMljB0dM3SoRfuR5T5mkzCFa0BnZJAAP27MrRzZry7ybJUvAD1QcxgO6XP
BPgsc4wi2/CYgDwzsxL47j7DqtXJfhxo32l+PDwremeLF4hspNXG2INNpEdHCGTk0Zq6ZuK04U/c
urbr3XEwUBfc+qpa0gJyq52hI+U+D3V9eSVQGW75dnIF/0ZWdAtQJdteSUEz7bc0mqsBNV0jZM79
AYCurJ2TMxmfCM2zN+vfZMxODYTT+dKPZNWj+STd1cneKABGpM+kFber9cYw0nxFpqWpQfAstKla
5AlCTpC9gKtACEzwQJG3kaigOev7Xh9TGl8Ytfun3csaUzhZnJ7Tkx0ITUTAaiAxc61KzgQpljLZ
BVxjybtVT9BYWrsIcGe68xutZNuzqQlcbTmLuVGPL2IeKWHgiyxevCxNfpl+VwkuwKk5Dz8iSqWa
s13pmHDIO3ZY1iLtwKXYrdIwInaTwFrP3D3VCdLj4zI5iMAcRNbylVqfiztpg7ST7BFRmPCyF3yz
M3fKPREvhXCJEaB28p1wLyJIMLSI1Sv2mS/cIdjqCAdXq+8RPsKGdecpQz3dCYqN+GBv3ytT8diY
iq0Cp1NKYkMMP8luC572cXO8vSLzSVrbsr8lmF0JJ6yB3KKfgwFl8AgreTZH9Gi2PXyEIxoDU3+D
IMRFqCRzpU9U4Q/CtL9s5aBDX6w/gwQfI74FxsYwWeTF0suVDukNLDbgdGttzZgIGhcxOooN97mR
+fjIpxcdLXJxTeF/MQAkGORiisngCH/6xOzxZoL4cyXAZguc5MLv0LlCGHdbI3NRBfs9Hg9jzXfI
h5mo3Yq5rkahKPEvcCcItWH47Q3xUOxmeUkJFDO1Vw7cK9IDd/WvOh035dcbJkTWI9vebAl4IuPs
b0dCJGxmLFqOAFBQ0eYQTkLfswMJmhcZF/bk59nh2iyAOA0btczQAPWqyEve0iKT1EFvhr6GMbxK
7Pd3I38/YleYICUy/QiNDS1u1eSTwBCVRFpXL7ENuF46QzaBbQkoK9U/s6ACnf4gF8Bp69YSwwYj
Bud9Dm5Y5oeED32CtHEIBljlYTY3OQU+HFUE3P1ckmCxq4D2YnRx2RrEDgYt2uRDbsCNQ4WLqQqF
kHc6Kg0JakuyLkweW4//cTP/BRcKyMNNoh8oNb6y4COhQaZlJ8faP8BOj36jfA7w/0qJAgZ5zHMW
yRDUhTMu97A8V2i+Obf9RnNirF+qmpGuSudtU6Dj+bT4AOTBL40FuB4ZFxfFToJrpGaM33CG6rvc
XYbA6my0bfMdBq5eXoQajv+GyaXx8rWp1CyG7aSpII2Er+X/1WtTn/vqTuy5UCYx3oA+YjZLzo1t
9qAY6GAc8NUB+MG7FhF8mujRJofXzOL9BLKn9WqRUC1daxdbWX/d3d7txHByQ/BLW1Et1dynno5O
4oA7Kd9hift6PkWDhwIL5ZAi6couBHe/Tfi9+4ZLJvNVDjzoMDos4FlMVvkJpUJl2qS/RQ9NqgVn
TPPBFBEludQTuYZz11/qE6L/3uUhwEKu4h9bLEjt21SecV9G2QyQO4ArP7+Eb2K93HLYU9rm5tAm
mxE9tpoL29lIUVsr0OTpmXaw5/5Q6P3PhJlg8M+6iwZ4XNogVzCwX7ujapeXfvTOMCyojaxY/CJY
jD4pkTqw7AS9E74U4XIzvOLGi/QN4pEZ9DTE+HIocwiQ5gjKR3HKF+fubWJcvMm9rVxDRlL7GA23
Bd8IXpN5zYnitMqHqwwFfq00AsRTW+xwS9gEPJ8cJNmQ2Ji2A8MGR9E3hFc14LFI2/P+mUF2+tEr
QQtJSgLW32l/9dynxu4QURyTxWeJqnYH9HAWl8YpikuuE/L1XwrxNpb1oeRXXPGQP5EE9clHEuGa
XebIxJPheMmjxM4S/M+e00xwegXyVvYebOg44c4qHNI4JRD2aEf4fhIMYrMmjQU6AJ4JXUCZ7C6Z
LBiQ2mPPYZqbou0Pw864axGIHVZgXOCV+eCtqWAN5nPBUAwBtT2hOdGIJsq7WZsedSnLaXwcGiAD
XwvcbKuwq6QxurbdedEZh3+T8La5dcIc2Y1vT06U2hs8V0a0g/rGV2xmBIXzD805Itx9rENcK9C+
nFfkpLHHc1EUJPeABbZ4iYXfArDFTdDH2yv0Es2ic1dhKN95ZKdC1iuf6pkBVbd0Esv+9/Np0HMB
vADdV5354CoD7kZNTR2zyhJ3B7BikyydAQWRv6Rfm/63BXmwCpfXfoPPToM7YWxbItyzPMAGXo/z
9Kw+pD/KNuuTyUPefCX0tXioHNKEHU/3N7z4WZU7ikJ2DezJAP86JnjRVJ2eUBNm0Wh0cjRhVMJu
874hLglkSs2+t5sTsGyGZnRqUNCj9eQ07LWvkFR9rTsJwr1kcreqkO2CglZtaK/OxhnR/iIkymA2
tbyPr0RftifCJZR7ZKBw45VpxMptEzMLT9Bd9Zfwvwd5OI5fUC8WvHkUXQMnz5uC1utPp7IUUWRB
fGjAAp6LEIr/fHMXzwLjwyvzGgo9pl5VIkSM75+3Xtmk/CJF2KvQxUmZpHfx8QxsXJAIYfujNCmT
ubD6FM7gALzxjA9c27lxZQr6XRDq1pGk3fJOvd6as0uhCR1wYQg6Wv511C+kZ+qRMcmlOI1G8Py+
Utd3P3P3JMqJO7s2fp0zExv/HDQioCSPjJrn3vazF/RwhGpJoxCsyrR8lyBwpQrViYpjljgIB/HS
tVu9EjdCDU8yitfsRO6t2U6rotNqHvghaOsDPdDeypai+QFwowcWaF23T6pV4MS4GeEhmk1Qhmqj
hPcFqjRR2dDhuwSD+Q0urkQi9pbpxyZZDSFAW3UYkYIgFduT87Id6rLPHZi4dlhAJw+991SVKt7b
akNAh4YTtcKlVqHuUkFV5k/CAReWJYQBatuJmuLu2w9MiO+7pGIVHnRjIZAaQZyurbDFG+f/1eBe
mnfqBuPm8+AfsqpDxW+f6EfvtosnJ6kA0WofUnWEI8HOGAeMs0Z6SQs4IwtLoduIYDvl/OAVSBbC
y4xScAVVsCFBEHa73rvHdYKVMJoyL66usrjNbkV8NTT5ZFDdtdwmZgQRhopn9Yl0qJlDouYH5vYh
GFIbVlhJClGz3vWqvSdPAuBfp0q705XoCdJEolDdy6Rj3JGuksg/QCInTSobgFlxGV0ZO0PxPEtr
NIHsWdTfQNvXRidTkpzrY6eke0b9kjAOjs4RnwPvSmzt095HpRnBWxpboWCSI1pnmKEycP3FWBNG
iyXLgGbbvi0twDi7rw3of4yA0UR2jV+CNKveBQ0czcKn2bYbvrn/y5f+f52dlxHTucLFS+gENPq/
eWUPxUil1BtXd0Ok3wSDMPwjHNYn4Q04XlCYQCWeqA0/CpPvxuZy2jUkNyHbiJAjDrbYo9EFdVci
NE6TbS3FPp77hChlLr3AJrrdSfWu++IWoEGzDButXf5nZPbNInt7WdHDqDsJsajZHwHfYZWLWBlP
YhuKpmz8QYh6vCpCsFHjSnfxdGOay1h0ISTyt1wRxDlstBCy0jKYeVeAw2rkUl+CdtmaN/67wjpY
BWQOG+Gy5QxvhWZEoO66qYwXl7oJB6YirlYibmExi2+wyr47SwBe9KihIsDGxqS+sdlMaqdujmex
O5PToVrVTs4Un+pyxIAdM8Nl0ABYw4krx6IYmvCyW2lxOIu29a1VS8qHbmM6kqy2p9L/n+FzfIq7
5inwYhZj12CKWWw0Gh3JrIb/26ioBnpwBDRYnIdI8yBGUHryB+2cNcJLuwYuPZ3dtov2VAJpfPuT
qZYem3p28zmgpmMmytGswsa2AnkH14J+D7MwS7I22PJmCWg16rgBfRoNViTn3196V/D87UG4btSD
dWXuO8ZohPE2/QN+J+JTOHq0JpEqDE+D6hu8pKlWAOsTdpAiGumJcITi1xEew8BCGKxYS6ae/P+b
UQCjCzQ7Zd9l43pwIM4WfRb/TTG46CwN30HHNxYAvmgiGsNpzcglAL6OE1tWsEoS1wb3ZBmli8Ig
3BY3tCdfk9maH2fQH71+94ndgdoe1J1/jFk9gEf45YTsQC4scnYeYkKeNLqvx6WHooiURVms8VyQ
QDn2ejuqKfgG7YU26neNBghyj8fZTAXIcWdRAiF4oeuuMHmOsMD8x6fAdK7vi8yX22zCCvbUXveB
KnbSSK0eTk05fodO7j+pfBQWlebSHQwu4OHh/qyRNpbtln6IRZnm019PZTi5vK7lcu3t4EL6UHml
w+yK2ol3CnfmbO77mZkyhKikbZqz94313ZIVcj/ewREkRxZTGRP39iFozKgBDWB/cB3uiictJHBv
8Td9roCQs3ngW4ZcTp/4myJtnuvGk28nZHQP/6rMq9SZSxulKeqqLJROpvtgB+N8FFar4J9SBD5x
GluT3oqHzii1wLxkPLpF9DvNCRT1MiFcU/cg9Jks1wgFfURsn9umrQ+KJxfiPgoFlasEX6/QX0FL
5ngEiC/MPB+SA6BK7vslIIBsKL8755s6OxVul9c7ZcjOy3aKWAjEhvK/4McJQEBMuCazuIbUG7pc
IcnsEP934FVmy1ciuIQMCF9u5SRh/Vw4gE0fzPA/oLr/Xf5eSvIDEx3lDp1V9O3SIond2ck4DxHi
c+s79UsH85bSdVwATfQCLTUe7iSQInwltSFlCvjLk/+Vr992/Xc8/EcCdshNot4/05A7uYe41+O0
/CbKVyEqGGqQd/QCfjUOYtArvZelUK7Qr2o7zA2vGJ9EBrdGElMYRwAQH/4lnOSYeMCWrmZbf3Oy
XFWJTgmI3OMhMzdBI890rC8qcaFxGarP122qmdZrsmBoJbOhYKnyAtKZIDDzWuwOAOeZ68Pkr5lP
EOZ1LeR+WHRueLyBBpWZvebWEWT0OPztQnti3MtofDUx1iVeN16PkQBfx0bVqkhn1lBMgzAcPccX
UGJ5+WSJmkFYgXNVXi4lKMDmVfyDbcWN0Tsl53zXMzer+8av1gaJs6m5ovTeBjmZNhFXlzdRMoOQ
LYNom46zogjapbZUiIcznMa6T1WLfTpSjc/zxpt7CoLMPwF6uQ5UR6DgM+fsZC3pdzEryXewSgQ5
MGm8plj1qiUcaf0VTyyinTOy/HjgL/SR0TZIkyHigEqft3OIcAekZCBuyJvwNz5RKsaw4zoLahT7
f6zsrqqgZ8d7zsZKsGE4kaVt3+AQRSjkZbTYU7RaGcgS2WAv5uYCog/MBetn7XXsiDcLmYSamTZn
WGe/y/24xu98oOdYLQAc8+5w6QlVqz4HgrHg71s8f5HnJg6BRoHBfyT6fZHOXAqJce+9oYy2vuyI
hsD6swWtXjRHQKuHV4Wrc8WZd2ACaG24BLnAeGCCsMDD5swfExJnQDYPWQLIVA39W4JnCW7FDw5U
/6SrQvXImc6W0KVAUla/L682EKUd2C+pQrOtVAT3QbEPDd7af+W1kyg/qpXD2Qr+1bsXvLBh5jbu
WOvbu1lMnbC1tSFkBwhQ0ukSl7QidYkG+iuRU5AyFxhgpjgN510HwHfqJBsmVy1qoE7pE2dt8CQc
/nnajwWqCZ+aou7ePyXn2tQsoy/eBWjqw/aHedAOI/Mw/Bbd2dnO8Wmkp6i3toN75YM/tQ0U8ev+
DVFmOl6iDHNgZ8stohGMnWEJc6vntA9YTRfUCyfbuRXVGHVbL9RRSQ09zA1oDs0MrxOIUHJeW5S/
WHTTJ8vm7kYQopSVQdQeFB8EdqmePLCBfuybGlggcDRy0DeEnZbwyZLezJoeYyF+pzm+SbSCr9Z8
O3c/5iGpytpeCOXlF1adADxXCS/+04TXpfbf3vM7G5pDcsD9G7uRCeaLo3zU4zqjmuWNO4sAMLAJ
sOz3HLlEeJXLxTCZjaK/tNdZ8lwVCb3GCRo1kzYFDkQRmnnoGP+yfZFapeViV+HX6S/PXAr5i1IS
A+FnCi71xPLPD/ZgkK9ZbIcbaKdhf75Qo/Cph9RE6TCEGp97s+dPkdPkanms6AqmZgNotB96UpYm
83+cO12yiJKm/li/RvkZRmvc1MCKTxmUUYbKFUbQKQ0i3COGIKrDLC7RObZ99hjeACWe0cC4CegH
oFE1NgBTNaThq4O2yHuKAgBlgBaxZTfNldBqZ/sr7EgDTK1A/E6yJIeEW+BuiMYG4Z+pckw/RVEG
8EzZUPzudiV8dC4dSqMMHPU2vhhyKdY0gLZx6Tzt/ZPrbFocX1YfYUB99Zgbb5tXW4kzSzffky8P
VqaHeLCf//f1EaRCKVBqqlcFoXq8zCHEelZz+ETtoB4Fbw0+WGidPYmxFZEa5Td5crodhKeWV4Jd
7pG2YB3Pa/roHACZE50b9HjvyHwtMOPXKSmH6l7aeMr+3xNI3ZaO4XIt6FlsHKLc4L02y5QAWswP
tovZgYDDR88w79Kfaqt3+qSHHM1vHW2h9wRKu1r7k/Mt5TE5AuWzX+U1g1fUvbQQu0yE+9b6IJUr
O9wu7Mb/XtFAu/eYCekgYx30esF+ajWvtHhRO5zck4os79gOEuQS1Fa891gI7T9A+Sw7BOxFxHpQ
W8XMS/c3RIgmZ2VKBUT7LYZq42Hli9C408UnRAGzHYVyZPuQv/J4i6YZi4ZChBBfNm/m9otzDqIJ
Sc5ODJNJPSanBhZUo+0EMb2kPOevhXIHwpIoneNz/OneBHlg50zUjF+Gr2R6NHJesTphVxQ38iFQ
z2O9D/l1xdGueUqFMco9oOL6SQYXbbOGLz6mcoUpFK5fAMFVW23eQ318VSn5/YclOt8cAuDzFMh/
mXQ00Or4j4xH0kE7D2s7DLT3r/bivoRpIflaz6+o/5C1xEEPbSWO9yv4YiBJB+KOYKEL6Nbcrvt8
5cgEsXQqr3GzIykoJ8QoWveAySgioLgTU8FnnIVLV+8O/m79H7YDE6I/rEITrTLdO/frasP7gkky
hOlC381m8gJjZbkhv5bLnnCMxk0rGXdlbgu0XSiTPOb5XpT+dXulY4hv00mIqpE55tmYVNS+sJ93
3+6F8i6HSLW4gWiPNlKn7IL+zrK+zC+fRQSxkgpNepMYatW5Obj9GWRqd93FEbTskVe4Gt1NsZ7E
VRsLiEjYP26iAvDKVEevbSozpIoVHDBUUTIA7LJEW3OEcVLscnQBOtEbneqPSetCMms6ki3Qh4Cz
5bBOTUWpz8fE+qVjCzxd6ga/sVKjY8sWYPv3YUja5EbAz00N2kz0e7kk68aF/Oe8l57nwBkJmYf5
UgAjDdvRRXBYCtEr5xLbCP3Lm6lE+CPLP3pQ0EPF2GOzDUiJFtNWG4GJETPT7VvYm/edNYWWn8m8
/nNRnauFwipHDVKD69vf1jFD9agiWdl30iTh+ln4OjxN3hHOsiAgi5ym4a75fMeXhz4elQQoF0D3
FpHIe1KWpr0zHr/7EOSvMo64dAMUxpxFJfjVUfrYF9+CHk3IbuWcx4pCeg3Nd6e30SuWMZVaFRxI
LF3DgMxWs4tEOHjVX+sU3ic3wN7wyb/ybL7MbRvHaLPzLUIk0zWywT6R+cZ3NOp9zG+P2m+PH4pw
uFRv2N+n1An29ouTS5MfnwkUc5e8/Q8jpBkkr1BxmcVDD0i9X00U3+PtvGjzOrNzAu6oBT1fmoAF
W8/vral8kHGVBxzZAJIaWqy0JpISW25LM7PAiZUdHfQmjanwd4zywZJznwAKaiSHPRMouFrlXFy1
BQ03OUkKDvM4IWJouD8cnllVxIyqgzXkJ5IDf5GrKRbqUW5RnNYWd3tg8PSPi/oNo5S4kUn5FRcD
olB65ydZgXod10Z3np2gnXB1RgRma6lHYAcw4BiphzOB5gMouMhYstqD0ViILM83aXrz4IOnaY4D
COUKj1erByMZj+DSjK7pH9/LSNkcHAJRcGfUw5CJnJld9m9Ufp0KjP9UtNrGUdAVVeICjE2ciUAw
Xw/7j0CVWraIZTEKOyoucVrRTK/Hge1/3ZMgLmQw4wrIDLVjb6LcbaACwPpBg0Iz6ZNA1hyCyvnG
h/YwgYMrHRk4aYxh87iTYpwW9kc0VZiNpK2g3pdetRhSmSLYeKYf/pcd6/zqFT0zht6KHELIO7PY
Rcqikop52XXRIDPr7FQIn0EJhqHhgvtD/GbQ1Oif36qFwsVuxzldLWmFWdwG/W0fH68ourE8ouNJ
PBvV0UfIuE/25kEKkG3754z5OoCarHgi9mfXUQ/G4Ei+qSABpUh1MDe1GcjTGgpCC17bejdwAu2f
CFf9Q1wsqJzTZmpnh1GjeM6Jy0FD1LLkbZa41etvYGkYU4qycwz/IWDrM+f/3yDeoTcKmAw6Jtys
zj+3DlXYxM8+DdlMyHEZfg20YDbnIaBibH1PRUN6V2x3IEjfURejZCbr2AWPoNP6orGI5yvo4Pdm
TW0VnuV+OhtiAjXU5oBMLZUF9VbY/1Tey9WYQvhbRWlkiEjCUX76mSKzC0hlYHLAOhZzSZAjN5FO
eCL8sTrqTC7wCPuVVF7fzFX3Oelczbpiz6//dTazebNIzu4it/inRs96o2SUIXpyyZ2Wv2bFvq2P
0TOkTKsQSU2d/vnFe4AAnpyBiHP75tNiHs7CeMfzC0uKD/2TXQYUX3w6nAmEqmVhCms/9E41Iw+e
fg1ho0+U9ulmILn6AtBI5ztYQHgUKsY2vY1W46g76oi/FGOFHDbDcwjUWWAcmfLt2bCGkrNwzdOs
PkpaOoRmL6mXxA30MQshQwF3OmTl81/7kzqva09rEZD23l8D20jcvxDhWQMKt15R8H7+F2ZK/0+q
QvXY7Tnt4hOCe7day9gOhCJANMfzvHI8wpFlbn2GRFCsmiezxHz6JIzlqZgbv7no24r4DGcrawJA
4nbymEYXk7EOvbI6wDSTUXtNoEh4RDHcBYhnuMCHkWN7RaVQxpU3uyI7sC6aqULBc0D9eFMgeraK
j4ia9oZ4bM/WBKcP+5Qpz3p8flOc4qLhkh5aphRn8J4kEoyV+RZ7iKERNZXr7JD3gT/4Zc6ADRz7
jE8U826SmE0/IPq8+3ERuRkYQzkY0Q4DGmj50d11yZBWg7vZUGCdrcV0ibO0wGax92WQLe+Z54et
3G4EYWORG+gz6NzPWI/biszESonKADP+wzP1jfAmXOTEfK3pKMuogjHFyvi/VBvF+rB2kXKJ58cw
dFLDa0o6grDuflut+JddxPvo1H4fJd8rtQ5Mjo6PTO7YRpdYe4oqYzunzf7VFcvRBESxzDZbYM+3
WCvcelhol8dfseu06vkq9TR9ON2+jMzGWUGAcXma+1NPwieb4msBqBgT0T5AUzh2v1SiiqJ48aAd
XLcwmVzb9D/7mjYtItpbDqPZB3JWLktM98KS/NReiO99G+vlW1M0AZ8wlFaUfcV0ZBQCbqvc+CJu
X5Vq3OQZV3eYyGOpcnQArwNa4QHoJpxULO0Fnl0d01LE4EMnfo4xMKduwwEO9a0GNbIWFB7peVbo
EjTsd++Md17AOPjMJ9coUP8BuC5e9lEzAeZfySmehDWGSHGQJmPz48eye9FwmfhvTUHIJkzDU9TT
34J6HUYhPmbrHkr04uzrf2r2iUNcOIPO4Xp0LbrNivyGzScpGyPIQddOCfjSd32V8vp+Zl4yWavb
b1veGZqwHVhOSw9oBTQQqDy48GZa1ogoxx4YmI3ZJJMdkH5jAdkwmsxDrWSlWM20CZLoTILQdEHc
43LAXw+IsWP18TPvAQ/Asr8x0EWfS6JS/vZNrKqRxBvMUOYTEy2va+jaoxBQ3mHvGer8dpxwAsM1
1XbKttv0ZtXc1xXfiaz76gSkSeaegRGkPCnnHB9A6bcMJ+u81CWP9u60WlbRXeZFAEno0FwdYI7a
vhmPwyjk+X2CY3/GzSbAhBLXWuYzYB0CF3bq1+cF8/nP2RUuZcSV0FOMPrGCPf9OHakok2BzUro8
cLfI23JgX/4/7bOgKAPJGxgVB9k+UwpByu8UmfqdPZxYnEmIOGjQrA0jHo/VNfohX08Qo9rGBCF4
+nXQq1fH4dq3a/RnY2VXb9Iepb8sEEBUAqzPPDFDr7QHDis3lLmO0eOrpqT7ol7pcv+92KVItJHw
XVRT8fR+i54Ek+qlILMd3q3q9kGXyh/+z/9jqbZLoedn/1oDHKfzD/O2ZU2OVJuPZ5qbdzrcyydl
+05cyM45LGxypvsUbWt+bMxp+9ZOuLl4c18IzqX9pOIk/k22er4CR7a6WhBeejzoDUZZ63zN2sOe
hgiQ09aK3+zAOQoIHhLDQTKx+1RlyLczHcUfqrsF7iWWu4pwu9JzA3lDlTVNElHY7o6f2HMCyMHR
zVNjrzscizbLUML6t3IdeMRp8C2CEgsneU2xw7ruMnvtZE3LTlPsJEDtYPQjhX47bMlmIfufL6oj
jABKZr6b6SYPAmIMnVdOIYsoXHRxq/M+SU4/T7wQ4bymoXt3DQUuwRp4tnOfhHwcUI7u9SLWjEka
iGU2LYdRzbS3F1G6w3NU2LV8g6bQTNOLdKwuSOKEHAh1JhwFGMljKFPlruX0V2u7LBUHn8RXGW+n
xMZjgk4oeEIuqMfIdd/bm+jYhRmaCmuBp9gufe1gl/dWf8F7gl1sV8+HW11oIH2bHoSQv6Jbm6pK
lbq36k0b+dcwFUr59W1C/4VG8iKGCjF7CixA6H2xbBQkVYeysdOoosajdk4uJ2BBxm2k6q/VFd6/
EeLE0qVPtdNR8SzVFHtGRdxfCDKU3Bnq9GROdTfyTN3Lrf5L1HczOglwjyk7dJOjhdtId5N0xJ9c
x1pLQubE035JN1zkCylHucAFpTKr+9O1NlScT8/pLAlKuO3sggbCcm2dZ44cEmSKmnlnDwO3sti4
pRQ2x11GpFTbKPOXWrnyErv6hSXEiRSZ8LNU11ZOBIVXU9JMhkp02IHnVott6bLEfgZMeUUO73eR
dAvHUEf72uK3uJ3JONXxI+9+3+dYh5pUqdYpicO0ZB27YLOAVFh9NZTnQYz0m7J84RBQTs6W2Ql4
nf1DQ4pCcTFd0I4uuiofW5CdWSYQIppIlfx+/OfAjQhCLJgZAY9HW2w0S/TXVVkfO38MHij9aeCF
2jo61YCFiVn8Lc6wsjaHOs8ZraAhaKIRutIIWxn53tfmylhdkL47NTbWkd0yeB3wT6O/9yoO3Vww
LEekLsTdrwE+YJQp9N+yiGiG09UIJ+y3CJuoNP/iIwIQXoy5Lj0pweVrFpyB2nQY2UOL3IwPFkhU
hW1KkPpgbYKOSLCrxxsS2jHVqRO7sXkfp/Aorp7n8p412tYB2XW7NsPav1DZGlWLqxUoHA6ePZ1Y
Rd8IvnMNkaRDOhHkNmuUVPBB75zO5HMcUr6yX+4VLuD+3w3oGClZE09NhQyTDixKJaQ4kCxjhRX3
IP6Yvlqr8+Y9T1qkPuXDh6fiA8+ASwj57apDhj4hiGPDP6+/HM0MvAJi+IPmpJyGrAeo+sbEC0+H
dLi9l604lR7OF2DbWW/cVg3jHkWwy9lJ9cAu+V/KLS1fgoD/0st6vTDAgt1snu5nHVUJxFIiNIfm
Gk/hV6NPpFA8ofPchxMDkfV5WanpEEsJCM7JAJqAL/ZTG/Wgs4nIAqtY3TNS7zvoYtrwRhMGIQHi
2CjZjr2KLL76lPaBduFjgt8rVjFlgPzRhYPfz7zbbW/VcMk1Omm8xlucwzSKDgZhfeKDIgGTHAXD
LVPk51ewWPtdqlNVydtM34H6CQBNCgJfwt8OcisSbAYJ6yEk6ccnqxEXFgiEI/Pny0FW2YizYLCU
gTGGVtjfuoy16exG05JK+LlVS/fGIIJlARgNwoe8Kl3tH5uQrFPbI4ZYBljnOY3Ad2DuCq3xdplQ
kOTUinjUz8ZRAH2oiUvuhcGCG5Y621F7VUPcuFM8Td7Mbj4lJRkUasdA8QU2dEb/rzFNHSIhKdVO
uhDShLVti6m784t0GAVmB79MUCqOePRI9DBT5mlMcJdZ2MZsvcYrmWcg8hhEZLbMfF/MDjNJ5ODP
dWre5Wk4eyvwMAHWWp+zMxd916S7FFgV/CgMjCxh46MJonUENiXQBkLP3dyxJJj6Gm/0Cgg7Ki4w
M75csacO/o2ChW6bHm1Jf1DH2FAmtJ5Uye37HbQXRlUd1znVXEdqIq+YLA3MTGX+7o5eVXLL81pV
BSva9qJP4tKmjducdp7YAb01y60F4yrfdOOQTYBAla64QELOOCYdQD6hGsIZ9fEAAlhk2OWe0Vtv
F25IfmXufpOUQ0VJlT9JBXoVDBknAIrNdJSg0VM9r72eIniz3XEsqod8dwCt0ToirgwLE8gG8lMo
6Z1IeL1zYuXCSNfcPLlHSO53wXoXyr6a+NFEOKY0b5xq09vxQqTNBP0jeiWNkJ/BBSPVlKGQEu6b
yjXFi3fyTyc1FHKpcrAPJDI2z1e2fS9NnZ2ed7W6h1T4eZk5fbCGO5bUnC30f+cbLkfegYFTqAMG
8uRIaJHMitnshHb88b5E/bJVhV/JSaRcE7x/6Ue7P63hyKsRhKClAmlGXHONLUyTqwHhMMggByp0
jyeNrx5Rc6ijQ5xwAPiMk138lQmkD3UcV2HZ7NtgKpnu8RjxCXRBm7v0KJwFBchJ9Rtq7o14e+7g
7gCIzrE3mKqV/Swnkc/k4aBBX+VP+7ew6+czIM4mKfPS9AUdL1SSN5jzCgZGA3FJmOZV3ZQ7vR9a
o11NFNkB429m4dHrL/yZwmzRag0Z2fM5aX4tYKNGOO/E6Tr7Y3X+N6KHDcalMy6DyiBCtbbIGSq9
5RufktRnmHiGdBCmNks61oYOOoTmnH/nA+AgawNudfxi53TcPVoGla6SHBVpTKK0jm9hgQCuN5FW
Y6vka9dJZFh2503zqF775iKlQ+Gd8t161FCMEfJomqHYrW3HZfqaB3UvioYjoMh7o3klj4w2D0Rf
xwBS+ERhytvfuKwcWfjHSnBHnfwu7dBjtUjoHyDivHW6yV9zq1MxhNGYRvpYFfb21MObOX9lA46r
X/3vni2LirDBDzXYilLVrRZz6YUK/QENJJouxqDfbUbZjAfTxXlw7hpc74yMCfxmbG5b+JfB9wi5
XHFvh+rCFzwpVChGDC/4wgdhz8WxQAYdRnAbfUgQMFspNjfJDjDJIC904Pyb9TkcFcf2aRmmQYqV
drkytTds5cxs9Pb6bZD020UmRFVD5WyuBj//UlJ1pk7K9KZPm8Q2MdKqgoPCS0BQWxCM+f9kNTOT
eimNnEoZ376LVh3MqyIvJ63foGtFKNcUrA8c241BTF8q6BIuIW1zi1LjYW7GoTg9BK4HWkRDg+W+
hwMO0bZXYAw8M3SWr6/t+zrDxuyGZmezGPlyyPBNCEQ335JNuDA8X4mBTDC6T7vTXi1KzRleVN+u
nVwYZ6FSCDcklBPpdhggLadFBgY2M/OdwjNy1T603+kXoTO3B+MSWpkysP0CF02A3qWUfdvAiX9a
aQzKc+22mc4u3TCNw4GDAbjbj+2bQ9kEk1PdRi/hvs95wN+YMeICzMx33OMm2+WKjvQk9g17CLQh
vWtgEUZewfcpjrHHNaN4uMFHiCjUbWfuDiCRq+MCxxpTrJ4oPot+vVHtIgtVJ0/sObf3CSQjgSFL
Qv6NwjBAGPJNHu9R4br+j8l9ej3+tTAWS4+I/985hUJhBhF82+hTFSIlHCQDjwzEPGNQCcIqVszJ
vxlZnJIkIJkC7KA0tqIpzcuLLZwhRE3P39uzEG/B1du+u532eZ2423FgqAF98V9zWETXOwx4syJR
A6fSFLOYLAZlzcF8VKoNw3n//uBMo6G69keh80ViwMKwj7zJGPRRIonmXNQr4uJBPiS+Y8Lansio
ng1KGiNu096Do4D0cFo4kXci0LKnEKlf3/jgv7Q9ILVFh8K+BndP27w59UAdPltJakBbqRFc0fnp
G5g189Ys7nNITcD+1fk1h4KxrBwlya7AGwyKPeK00FAxX3HPi6pDrqE9QFi9aL9a+kDxM7qP9kCg
2hcYATi4cV7+zgPpcXTUvotWYbQgHlhs5TSZqyin1ZW+Vx/dmlxufIZW2W8IKOALoJJTEE6EWEnS
u1c0yr0KiVZTYVWWPaLz1U1ZHb3Ddo6GoZ9f8k9yzyVCSsG8HXCoKB05Ywn3WmoiUzRmporoSrZs
f8mUf8vzP52vbqdviIuscEVuAkjnGOySk0JYRXlp9u+yVLG5ec9WW3gAiHRU7lYyXT7SpOk46zPu
mNUHo+muOfRqZPYsDX0VIe1JZ96A1iDj7udQHe9bJU43zQOCxz6nzDoc0g9YhLNINQaJMksjFSVQ
EpmqkXbIHsK3mmNGGmP8/OgY6wFzIoNuEGX077UAFId6uqGvM+lDeTXKxztWp/veFqXTBG2XelJJ
8FHuM0bdq4wkpVcfdj471OBymhZrcT9CyKMl9CdxJ3fjeV3Q4OUR+9oJSkFEFyZuzN7SX+nAeRo/
arEQAVsXJJAbqxKfUy6J5CNcpHVJmFZfX5EgrZH+6gUOSU+bOarrdEFzgEaGh7fSkH/YVArFEYvO
QvHw20UEtttP/jUCUSxxnveCYhu0HFvwQ8XfSGW0O2v/cjJ1IGdgyMmhZ23sNsiYSSZT3eG8akTS
uA3N+R7FghAK3F7SkRqXU3Bhbc1/7i/EWO5tlIH8rScj/VYt/O79C5OtqE20u3xiKRDgv563EI+u
4hQHEuhHGiBfvuAtKNdXhOszHfeetH2N6IzenOIkfRZ7j4dlyFO/aKbH/V5eB8TESFRVRkrOOsLn
ICM3JGDnnVG2brQUu22LAJp0hQe2pJr8RhUhREkf2VK+vZBq8oZbG6NsqIjJTVTp1KIa0f14tILA
EYP810bP7QG28ACr9CEW4Fis/CC5NrJDzIqHmp+TT00sM3rF48IsjpKt6DU7XxnviinLcnwBpQeX
KrfUpklQWfII3DPTxU5T5CpBCvrfQYBqHdIelzBOWafb7FRsAtF/W1e2rASPXluXWDLM/Ih3a0hV
59fplahNWiaBwaa1RJqtaE/qaBt8V2/njs8/qgiA9HsNuWukq9CXEPX2mUWCNSEkSE++IbLVF+6t
YWR5QPnHnU5rUJAWU2nwycubnZi2jskpYytxeVA/ncCb819rALY2icpJy+ZoqEzeAgvSlye3BdEZ
DbmQ3ma2ysoBHrB8VHOXjm4zpHkjdotDcHM5fAFfr2d+qTXpJanCMVyzBhVtkZry2cJ9LFucb7eU
DBdds9xyPgtOu9plOB+ymhgQA63kRoLPjR21QIq+sug58f7cz0xyQ96CDhd3i1JmAPrujhLyOMqz
u7/2TI15r9HWC9d/nnsymJfrXSDchIHvNdGbBMBrcJbhooeEiAzMR6x/1d3ShEwpC1efc9+qBPQb
lZZoEwPjcSFMkNa4GUAvGgKWBd/OgkE+T1aolR9+hPyHRhUlHNLT2xLmmNFd+hqyIQ60i9adOf8R
hbj8uiY0oCgIMEejNyglGNG7bSDB5ujnWDNHAgzB0xcqcQk19bAWsHXHLpu5jFBHtj8MdeSMdWxs
y1rAgWTExQu5ZwLOHA3gt2hiM7avKoNiDqUqX51qHBvfGqaCxK+AO25cxgW1bdmDab7Ck943tyyA
hu5NsNpXRzNfrBsF+hxR0IFhDx5/oei/9c3KIyGOyp1Es+GwCVsMxVW5W26lfqYeI/V99R6asKOn
6wceY3K4UkR1U5WHTLwRDMW3UYbsfJwhm6tVldw1Lvl1JFc0S3pJ3GhOV/1hhecI37rLnYNC/PIc
8cE4Uz/icTpEtdUmT57dWhv/32zT4DbKzSCykW5tTVltNIOhEeGzFXzxo1qOluYoj3jgAank1ntF
3xH7Kok7+LgkTxePvnDMMHPBUyywHp2CVEqCiL1jsX/WZf62Uxhef3SM+5etHHPG3Xrgh+QIvDsZ
Cd/bq07jd2VMpj+FrVHHpdYK4c58Md5TvkLCBjtqkr0sq6PxY9b8Z1rB1ZroLJCCtg0mUhQ9uoDu
9vIbv4so7L7vFxAH8Vx9Sku+IfjJ09lxto8BpNUZNYuoh0hEu/tL0JycsOBfzZduU5DvFb489+W6
pl0tasJNxhsLbJB/TI6bUKJcEXk4Fbkr7yJDsGTWbIflhgpIpGJEj5M9HiBL7ELCv4/O9irmAMNx
0PTBsUwK+9W8fKwFBOH3bdgm0tp5BHKs8TfmoKdDaTjZN3A7/Z/phBvmFJc8leY8rke8LCWQoTVL
M3alQtWgqoG+Jp+9XplcH+mBNTTCJmE8035pxkpWGOBKlQN8BWwd+wA4d/NiH/mMvHFDn5URPfIw
TfwexHcmu4OiKmYsETqIUflAuYisx+DX42eStnepQpqva2gHKbBhK+QU/p2XPi66VYBmi4v6blJ0
h5vZwpTkdeH9+GWwU0X7K4mAnDWARpoYIs/jtFofwS+spNyp0MYJbGbtpgVKBBQu970Mi6xQwv+m
1WSFx/pF5iiBm6YLWB0mI7W9h9FeQJV1T6HdJ3+eQNN7V+WFB2BIqiVTIYs3J/+es7hjkSeF1gks
XRKQu2bPOTf24/CZ47aGHgtzUy8EDx7kazmfvLy24n2YPFg8ZkLVXowyDs33cmep3hd1ecS4QhAs
a1fl4PvwDCG7735Mqe9rmSwwZO3dRSF+bSOfPE8bi61gL42TAhSSPNQV+biwe2hMLY3IHEvPmaqa
Bag6GXuu4FFXh26tT64x6ZtT6Z6EiT60xpXQtGWjGvV9i6yH0c/Q69GgcFVQqEcJgAzYAJa9D9Am
XN8F+dugTLNZWr6WHLILXFoklN2HygpKRg2Ge5GlJnoRnsxYhHclZbriD5fhvebXygc2YtsKChlx
yI6LrVs9YgIg50m4tqSuTP7SCDrHtAzwPXaWJVH1kvpCL8uVeqIWIWsG2POFmaFzDlDIodBkDd3P
qxMI9UGKRl5DD0rh2LujIWwjvZEeqgM4KrCgNlgUYjku+hqONbfP1utVVyZDcyeY56Q9Ab9rXWmC
XepZsvLbWfXL4X5W+AM0Sli3Yu5I2kbIGiQT7u9mTE/cGQJocJB4MYYW7J7e5zPsFAOygg5va7vn
+jSvQ5WR/GJJWL+AX3Y97OR8aZFJFAVw/BSHKgejZBVtJRp+oBOk4hX+edNnaax8dHjmmXN7XSkl
AgFUk6JY1Nu7aDupfdZNsMTYSZa552cLPcywKd5tTzL3L0X/+Lrb87279w+MVVJaDwgP0cabYAAe
8pGj7Lv5uWhKEdOz537TjcS34EksO/jCRkWntLJSLfNpIAsP1wIDauWCo8TFuJtK4wRdfK9tQ1f/
LaqyQR1oQ/0MpuWrtuA+vmch7CUPgK2pFC0F2AsR61zvWhz0etmxG/mp3GYph5BUqS1oiAoqKOZE
V4ebhDSmBAQh+rG/nq1fTJ0BcrdNrJCsV7yyUO7VzkLsjOYw9ab+sdptym4U8W5tjWnpvx9gD/Z1
J2YC5N4E49pkrTvHGx4GdHRiguh93gjQq2J5eponWUjQjiewRGvbdFvl5mMcT5W0amU1DaU0AEY1
PCJANVvr0LWHQ9kCzVqJkDl8xGny0u7Vru0P03MP0luxxzs54DxM2fww/Xjq4BKgmKmXXyWSHer0
jgdMD4VqdKeWCn1IYzdUzBowH5GLKgv/PvyU+QX6QL8nQ9NOZnsGTwu0hPJSYK0FtXQJWdPHITHx
Plos3dBOQyT1yGDwumDelremQ4hIabHwm3ekpREbkyC+fMb5f3TrwHok1iA8Uxk4VVzQt697Bz8O
F6XnGKN862b/UFb+Tkh0XCKWctAEniA/WA1oVq1TPAjGC8hZWsa4cdYaogUzhCwt4yG+QUn5wvWt
nl0s0BYck5GLLrUWZkoJHlV+beCkBUwCQoNwTzjjrMMbaxJHhfvzUHD7iv7jJuftTOVKKZWyT+tI
vf9Q1GYLTz+Gn8gvG/1Avt08CkkUII9AbUk7cM7/JoAAG30sO4ODPXd5vjiSHbVZ1lkKdpDK6rPt
+fN0OIOZJo4A5O5/5b23vxvBsVUoeNOLdiZ/W9fTa23mFaJ6OvprlyBNREU45JUXxeNq13EzpCuO
ZdQjbu/YcgU9SqM2C5K7yk1Hc81XuDE82syBFX88YyQhdM+FufEPuZ37AmrCOz9Y9ybAg1tlLw6R
8Y3Pvk5pmiQmTgG5NmJZfxGw2a970YYRW1GeMB4qwmWdSWbQPZuaxg94LMWMyadlIX0woGNuk659
mTAH2vptJonzBak7luPRTZY2Yjg3wwZyf12TbHeVLXgJzdh2oliUlUfwwCOgs29vyt5jTJvYkgPR
lwlrrzf7emITL4eGQ6EedoIPOTB6SC2EFkC29WMV5Qc4s7Y0xeRh5xjHam+UAm0+bkE3Umqrw0KB
9wTzoD0dtV2il8GQNzRn93UCDRRyTsmFI0Ic4u1Fh7Qd+oi0wZ6JIIQCOWOyp3XwwaCkxJHu6rT1
fjwdrtNrET/OP1g6KYjhMwCIJwN9GPIssAt8waefmvU9Wg9IBnTiN//j1IpY/zfg8w3QLIyFJmVX
uJOLVrV9ZpAFPnuUWTnN5NRBv1sjVd2bahdwdLF5uHscBHAYEQq/RKT71tT0nEJ5kHrlL385AgDN
9Z4mtAJVSBtiMLgf0OpuAhPVM/OHO0al57e/xgirHCGwYbLSy7KWX1ivu236ugGnfuNYBrTwKKkC
592EqjvMjDM4/xus0gvBquns3EY4yjVKxLK5iF7IYQpas1H07URWLbMmfjeKPzH0cMlKDhDdDv2w
hLINOQV7HoASsE34uWN5jugJ0KUVwoK6Z740Gg+ZDQBUBWzW/fCbW3lLOrhsJPgg/Zro9slsox5m
RoUqlUYwoPYA7t1i71SogaWcmfwB3QJcUkGABIW/SwaLdpb8HpGboIrGlgqW+oLjL2w5NqTcSTF8
XrqhhD+yVAF9zNeAfkXcbUICHjXm3DTo2vhog7n607Y/vvcG+RPKZYc6SiE0Ytv44LjVoIUrLxHU
hehW6PZtVGiB8q3A62G4JZCdY1YZpGpUjGoGgmi6cQAARxbd+h0tf8Kus4YPcdU9P0rPYiNHxSx9
N2MgHZFkeoW1CF+NdtDvICSYRnsEm+42RtBJJqOVgRtSu/aiFzmT6szxfj5Fut5ZEFVSOTwHScTC
a/VPz1tAWHDh8hDsd8+Fier/W8vgfP4CuEGnz0Jd9HOpOBsZVJ+fOgDLuGxv5WaxqOzFLU5c/Idx
jHwbbb4IDr4727J2U70IY8CE1PTFPon55PFgTagFtNut5amzY7OI7NO1sz45Hd6UyDem4lMiDOyn
chMy/KOuCRZvoyOiOgqUrNj3R492SP5pZmFO7I7zeZDCZwgUtYa18Eu3CLysZ1VE6H4XjlQ1SnRS
FbuO3Lw2ef0ZGojBYL9Zt9K5Vmjr80cBXB69lj9bwFtOPP6q84SeUnFWr/sTXjGXDkF8JOZw6lqN
KtaUwOI7nEUJMXbChfaXh2RXGnbMRwtA6K7IXFc/xJppaGHtprdDoFtFcewhMwpVJAbxuTTY44RH
RTbHukxYfUj/hLnAOwQRPvxC4myywkqMGC9xlOQVXeoM4py4+oXNJgoVXOV1DTksFK2WpepdY367
7seaYX6KYK4GTAQidTHiEmfWTps4gfe3CddKX/DDICI1hqZOtW/m72CKVsmbC5+wmH0zz2E7cuVV
qZ/8OIBmPaTFBqDicANxS+7JaUAed89DauvswXoyRVYq+icg0r/Gte2MIf37eSbE3IKUUmHPg1dy
IjDuV86/Lq+k+3/PIVXXvKnVLLiZSC+higkrYR4rKSGe3PuuzvNRrsx0qbzl/evoZxmV5xyhuNJK
R7J3rycJFOQuQwv8lccuWBmJplrGPddptFhJkG+urjYsqdVExTFOtKVac8tiZZ0f1AIeiBEXRh0a
aIfddq+hbLFmkErTqzN6pGhd+Ko6lRYYLVqZYsaFel0OCmBSY20hoM7eG3fqP3kslafY+2GHqQcR
d/Kr94vN+8VTmg4e2KkmmvUVvT7z2xuZHE+bmzCZjiezQaTCq5t6VvvmHtx+Pt00Q/7l2X4dVel6
1GKUzq9ARUgA6vYFqxBSttCRpbBhPd9UItjtnmAWwHGWOPL++/d2p8oivaZ72YUmbx6Uol15WlkG
bmmAhrsuOM51Qfn1u3AFbSzMexFH2VdkdHpRZFMY9s2C7AGWKhSJoZW7zyyAdLJo2NHvjDVygA7l
pEO1MYS2j8d24Kj4rMSjFMUXH4Ed3SwhkNa0Jf9Biw4yL9zJNBEL10EQMwLZDOszNYUAwN3FIfh3
RyCV7rqzol0xjXNvQlAL0il3N2Bn1IjQIkCbZq5MTTfzfCELX3ga86LoYLzlEkDvgwhsLptu5Z94
9kxw42YhOfhH+8hX8PAsKuAk/z1VvJJD4g3yOePghENyOSzONjU/egYANzFkSXDO3OvvPRaC8Vr6
R8Xndej98dSrIFt6FI0j2zdcO6Gmy9Cyja/pH28IkMbPitZ/xGeGYIDOIQVFd0qYErSUW2Bv0i1F
OCOeIMuKjaV3oLsKB4drqviUTzRpIXQZxBg9W9H8i8jraBvYM5iY4CtWTd3IOdr2rAOUtuSZ/ElA
rPF7g9wdlNOfouVvsx76+kMqWME+oRyqmsD+eEL0kb2DSM02oEmdJkF1YNW2JYnMsOVudG4wzfBT
+fHedIHu9uxbAWHOoaJOeFkpWaTfLp8pr2vqPjUJNxXnoU/ZtNlPsELY811hXNVJjgIPrX2OzRY4
/GbWFWfvYlVpgKfFgfYsi0lIYsLzQsplFkjK3w0MYRwKiPODwna/uy5pycMX43nXJLFLR2w69osV
RdQGcyQJa916NKafu1OozvvtGs3b13ZLTTQ1o6ZcIQFlQ5UREX0K+St7JCPYk/S3hSFwTOuxqTRd
0NpwuY/PAdNsG+VEcBJm7czmgsdvrOl8Kqnapw6VJrrbRJaEqdlH/lP09kvZ9ITagW41uj8YrFjs
/zfN0Ec8bDNZQukk/2MunMTjfWUITs/DVJXda2lAJsuoawazEaDBjjsXgFX8OygYd4Vcwz+bFWwp
E+Kgw+83ztmXn+D5qt1JFuMZ96ELpWkJFI6vzEyBhP9Csfx198sixRbaVOIyMJqRGnT+4KPNyUS1
OMnteXe1+V9M7h3xD/NcALLCIG1+4+bzIHUWD++MNrOCbxL6RnjPjuMw6sDnF+jnRAUgu6ZsJv3K
J9SzR7WLg81i6OHIRwCkaJbePeFIItWbe+n+Ym8M1ya59XQyr7Ok+QG0n9swaEue3lsBRPkH4Q8Z
7t/pIiiOCaYUmW4MOIAJaMtWK/1gP1V9933v1JNbW6VAPKsYwCuHMv4CyrWj7eszir/xmwy4Gc+G
XjtFGPgyae9ME4TZmlVtJuBJvfvvbkWWJtXnKoIPtRuYTkkXW7o8yzoR1BW6ZuxliCWREaVzWzYk
MfZpHjIW+O+HLfmvNuixxMoZnVuX+x45vYlcmteRzlPw3UItzfBuLHOezJ7V4GUeBAogHInl1HPA
7U330no+wid1wASUyWl+4izhc/H7MgvXx+ZIp6tLx6jEglYEp70I/ducXZh6Iek8MU3FDdCC7ZAv
wVz4pqVpfDwGOa/oOfB6bwWbetuOVc3WYhRjXU0EKBS1Rm0RERTAEmwVcW41auK5ht7eLLUnfMv3
yBJQfmNGtX+B+Idy05zQfx5pq3AxkXgLIhihAdalX6unDVmdeKh8/g7yITRwu60kyJKFijPjQe/E
D6Yo2blLFbdaqVbKWm5vTTTfETAIKPH3zaIEzr5bwiMXaNBjdnaDPnjAWKYvhN4Hu7c9lWSOCZgU
BnkQ/mQtNg1lzsJWN+w91e1e6qy34k4bd5T6MDsbyqsIpSw+/GyftROuibCnv1wjPv05XioG4zCn
6teFkHJ73m9jzWAyEX4zNBFifu1zJk4m7xR917k7ghye2520ifDnT4BRreiND3bVVegGxCglQUjf
av3nphebEbKHGm5hMF81B3kRbN34LXlNpKIQbx6R56PGYHrn8GBZ+gx7QnSII4O3aXlVjjnRhIRh
8zvSM9ehMkk4nKEgWgmsK3Ng5OR/H6Av94q07JBTrmDHvX/iLhOZZ2i9ivpHbTtWp1WzxZ++8Av0
9+r+GqtRnXBnw5tOqh3GqOihDU7QbblJTFwge3lARn3rudaek/ulg7Fp3uyLniv4y89OdMG+WmuT
O/TdagA54mg9ecDUfNqlxryMEwFVt/+9+0prdRFOlwTLIUrcLRpyFJGborvEnuGfkt4hW4ljKbtZ
JQo7KlNQDgpUkbZS3xT05o7hhWEGVB+VbB5XjDJ+CX2r8iqPheOXR8ExAp0mOUtY4feb3PpE677X
/0m2VD43vH6/G1Y/P6ofbCZn/Rd7Ie8E7UdfpCPAisnNqD5Tgni2xRv3BfVTDz8DvmY+sUhJklTj
cPWSijbbqbyv0LzdCyCQmHgrG32u+DrqIsBQpTutnLcBMdU8RbhInKTYr75e0XwrR+kdWTXqRACA
bdHx5dUN28e8AZphuFK6TkXIYBO/RiPrR8DborNc39UxI708TT1VrdQMkA8Pbaqd2RL8LUQKYRIB
mcfkRId5NRks57QjF+jJ7z76qXBRcq//ceLiJT1ANNvk1NQHpriZeAKYTrs77msN22bCSMNGSvhv
eK0jT9soJvr4cQSOIw3qQN55rKuuFE37ISf7xGoi7qWSlVhOqSdstrtZSD7d/on9vC8VO0RT2I1L
tEiksYZyjtqIU/kZPLOulPzz3vyOtz6baw2ZuHFy779+pJ03LUaZWMjMjMoucw1K3JYvuMHF4C/d
IiKVGZYusLfVxEmPb1rB7YwnH3PL83It/8ULzWeDolU3SuGP2PiE9n4fl+if1UwhHcNmfOF7UhH0
sOA6BD7A3UF9IEamd7pC/zrghN4DQiCIgSfqW8SIXNlnZ1tDx+kQWFlk+DOhfvnH0rWeVDPLI968
EWR6r9Q2AlaOqVbUHQ8HEnJxa4NK8jVMa3mMrag2n7NA8SfByKXDhtTZbwzlZh9vRbxpFOsU8hUM
eycB7TwnH5b2QuBO76SGcWC8DNnpoamrcovy+LahRaB+qK6ZkkCQUynOrhdPHMPHCRwoppUkLuVI
galXN1hn3VUyiH07F34RnymofVxFQMIlkuo0bmLWpCzQUQkC6mtuGvlaWKKTSf/S/bkFU3mPnEv/
S4ElXtzey0i1k8ooUb9XPUW1lzoreH0a9cdB03yPvf6OZneEWRVA6Em9fV/7YIx2Elwfs1GIR55/
dGWuJVgo42wwObEACcDoTXeZLwzE5tiXh7HLxJPX8uWGrwlJm5iyXyvqJRlJpGO+SG4iL12sO82Z
/wzmX8nX9EsOJHEJ9CbY6tpW3JSaZdE/V1iBoJVhm+A5DL9BKQfXh2ll9XdViXhu2rm4+h0+j7Df
E5EiTMaCDyPk5nKEZpH7xYerPFPRRIm8tQfxT85agtomBwJQ/nf31XaIGCPPNswjQUIT6e/Uf/GG
PBylbtk0U92Txo4p2vPY58UMuadVxRZ9qQhAigvd0kiuZqyCW4UIznKPK6T502eZMEV6+OEiGyj6
2RXBnHHoTU70P1Z73T6u9Y37HnTj3EzYbjP+CAe6ZEVZqVpb+dY8SX6BNjuMNBYuHeQHHJr6oDx8
ZTDYB24Wom3tx2CkCc/3fU7Diti4C2H1HFd8MoeVHsxchISOhbj07HFVsAYML/c07Zw+1yC3IpnY
ZWwKeWDkA5QryVpo/EWuF80Fxx1ZXKMrQJRYHN2Adjz1wNmvVBGIzVxSgsp0mkyUgqgx5lOVR89N
TDtG31iaKJxQN2TM69msqFZx7PjnuGWM/YTlj6poUHV259yaL1mS9P4jK844z5sQPQ7XsOk0/VEv
IMBzlx8VWUJuhjJzpo/sUYSEr8kSgHegNlhdIDYsIcIggjyYjyRY4drmPMy3WASSDVAbrSnLZmWH
lc0tLXYwms1v+u6YUMNZFr005mSyTEoR77okRqyXYXIHs+tXq3Vvt0QWSzvNGhNSQJ088V9bs7sf
Idxb/gdOgGJA6FymRItpf2In5kMOQgbScbktDgjm83ZsRuN1lFS9+gg9fYdaV2Gs0i5hsKZGq0gT
RNAqJrMLIxZXzjsy3BTtJuUK0/astvFede+qZ1CGT4vP5lJ4OtBhKnO1vc8WaU6hXWViyyDTC8Ax
w8d+t2ciQ8H3WfVHDxkm7vm3ITbcSwdzJCKczLzGL4iu1JPkyReQKhvG0A98SZrXNZziJ0G3mU89
1pDc9UyDYGPawE/+i16z/R+OjwgC1sg7zCkPhyd0+TCSCr1b1SrMbDrXvcS1lwH7YYDkpQpnQWxd
Nqc0DcInHr9Kbl2KJ+/DU/DiN9erpGIa1iXybWu/DNukrxdrSBJnft7+3wI1vf5RyMHCtwlJZCDB
d6z5OQ4uPXNtUsqnHqhNt/EHQCtWyj73zWAb9f3lcxT4/7M/nx/p15g31clox4emIS8XebfDoIz3
lSnAjpKDHMU6Gvvk5lDouXVqNjsTzvY1O2QOulUsDRkhBaooywB2hZmB9m6+x93lzbGIoZ+YZGHX
6DCUEi9TjK5xyRfi20ro0xY637+QviKxrnzLUewX+T4RZBZRpezT1RuVR9TkAT3SDnh+Ubv8U6Kk
ulfDrnSH2QSydhb2M9hkz4cKGZyE77dpouwxucpcWTQqsGFbLXtPXji0JvQ3NGH3oX7PNC5aNrM+
qCQYmS7BZmKUi5pvm5qvW1ohl6ALFz+oH9i7gfIANJL9cSFBDfgG5CSNqNsZ7u1Rj6N6H0iQgwZu
PJTRtUEImx4YemjzGRf+m++SdS1RvfM88dHQaApb2w4eXPhia34t9DYogJS1/l1nRzreVtrCSA6K
PHFEd7wxYlQRo4whujtgX/BPbmXUZ0zWtRmm3fbmljUp0lur26ZbERcTCvhI/1Jw9QjHPj5hKCS1
qO4fBt8pYHwZgTknyBdeivgPWn4I4ujmtN1Y50V9gWfNAtDTQMR/sNC+NOgaK6SiAF3aD1I04byU
eXBli6Yjrl/eJIo1ipDZrVp0IvjevIo7Ep7nbGiVXkCzAgb3lunj9vKyugfnTywr/zZnIrJCJ58u
6+kcuW/j3kZ2EPWpCdlnso0V88Ac8R1q56+VLDTsNM3nkeH9imvKxfg/3rwls0MallZGRE8VIfZ6
jAjnD5fsJZ1ZERfoHYWg2PgQsL+7Ou2RrGYBJohczyyPbSbKca+I8JjwmhP4FtCwBEKVcsD4UmnW
cRTRYyD/Cvy8mj5vdvK8xrsQrG1cMViR8ZYbWiqPkgJceijbTXBi7csYP6PY1qwaH3IolCalinT5
Id2LP6CRX7jCHirbt3rET/y8Ap2q35P/wm1a1r3Vpwftf01JMQH2k8X/Kk3MVf+fbrK54z0wT+Wv
m7lFbAeBAtkCD3wVSX1widZ4zZF23cyZDI9cXIHt8zLCZz/4J8alvo33+QGKENXqcBMF/U75DMVa
6IdfZpsW+iaCp3svct9+BpGZlkjS8aOZxmZtZp0psBBf1lWY34BfxN62dbjjTD2sQ9IqJnmpYGll
v9qS2FzZn4CMaxHREGlBZHw1Rkdi2z7uP23KlCLWR/l97sJZaJlHFEGB1kCduXqOG0fiYR9bbvuD
WssXIIaSDdz6up33W51jmhrOugE4tlcKGFovgXg6VOOOZaduikCq3huBxF+nqLH8+sg9SO9sVMmw
54+9eaLo7SKRSFkQbKHS+1zJn5LpEK2GjF+lgE+LnaALGVPRaDF3wrKG3UZuEx55ltYknbFgUQvq
ybEilVqshTUTabzWOrEGj9Mf2qDwoy/Ve3RujX/FsQsnsTv9wbccHXkMKug8meKDWBp3xzrj0D3c
Revouz/b3glxykbQmAY79im9B1VfnhPAHWBZ/6+XPkz8pvzKawSVD0m8W9FhVV8Xyjmi78SmfTjg
nZ87o5XcHt5CclMfts92mZeszv8rHa2FWwYsiDOjTnagm389TnKOysWABeKRbhlAhjB+3Y9+TtYW
UAt7fkOPFflilb4KfUSE9UgAyJUDWBrTSjpP1Hse7vs/DBB4aQB8FcQaLH3dcqJEApFCqpcIh2PN
KYu4YTYu8wTUZT8YwtWWNItfpNPyScepZNOqu3seFK0B0TELia5CQ9oVfLDd+ItbXXDqQs5NwAUB
EvppcC1a2xN00Td8uF/LwJFPf4zewApAwUbJmHxGSaoaGFqy+JGmvWgmNK7QIM69JXuzYFAFmSf8
As4r3dIowKGCW4o6Zk8gK7VJadwA85abh4qayvaX5k5aLDXwmO4dZh49Es+xV0LEiRmTDKvnA8kd
2n5wjXkH6fDUD7Y29q+mPo8ENtgJ5EQeqfP77O745rzhuLcek3NkAv7Bxl/jxexnvGpXqMHQzxZc
qQ+jCLS87K9NUp7EjgyXUMcQGWOFMyVUEfBZ2xBImmUnxef/gG4Gq7KTWnn2K7KNLr4/qTtIoPgI
RjhFvuhZdKk2VNqYyqjEvsfB/dVeNVumIN1sP8BWnrXMK7xMwLR5avTKGgqmHsG1O4/sKM6BQNas
d8b+iVlg5yYHFsGRJDiiFO8GzWlV3GRa6uHmSA52biAW8eSrAQMRWoBzBWBH2eUZYeHzBlK5LprB
ecwoeMQDBX+feZNK0cmRgPZ/f8DAckAI+1st81gJTtGZ2Tdy0te/56ULK7VmUri6Kf/3+wF5DZ8L
Vzw2Kr1Lg/b24yK/R8WpcPs3rj3gPS1O8Lm7L97wftF1lQrqXICAvvqnwaqrNiir8nicAQ4ysKYL
sagVd9a9hpoDRWFiKTagpHkTRwZqi6U6N8v/uv+pf1XbWdOUCgCog96cWfTQ1p58BuT3dO3wGsr7
xAkoMpunJFEWuYRowbzlo/Zpd0ZsG+mumzFYw8jqt8/93iiWDnuuaY+q90Rc9Ow4dXNQuGIokRup
SJ2XOqo07sf02kribaGBuRJtq+ogi0dBD5CIGyy40jP0NU+89ZmeoAjUak/VjB8kQqjOZviW1V8p
OIlwHJRUqTdvN3JAoAzQzUZ9jyTXzCaWjv53+eENb+yils5E61diZnnOUts9DL31dBy4DBjCpG+1
oin3jx+zx1xkhwR+3U8CCS5mWy2CHQE9TC6FTM2qup1bebbPbrb1Hh+DN8KQ0aLanu0Z3i16O3zp
srnyI/0q4ByxUATaYbG1yw3XnCdvOBL/vLpYFO/CvfcsTH0Luooc0C5Sv36yHDYEhKRKrvj72oYp
PzRAaTBwgF80vvQeaLSSrJeRmNXmJXwx+PXTVWmRTCsfRJi8Gx517aywtFlfuD9Jv7xp+U802bpR
Xsv/yHjla4n+ose9FpkN1SpGrvZMqNkq2Txerp2Wgtv0KwbF2PkofyB0sDc1RizvfQBTqqLbGskQ
TvBGYSAn7buRkhjR2frvjPKifA+pEbyxNeJPvLVpW1Xm/Fnv9ccTKHta6kBppWrBEZtYelsr7hch
frCr1Rn9edRshb0/ntYe8sf1A8QQvORitwIi0/1hpFnC0pVUwRRbm3hgb2zwMYWVV1A5OgHzNYkW
F3RDLy5Tm/P6nKZsr+dpHeldgi7Bc+WR46Gjp+TT5YO9dco/ybgmIrJQ+HbOzj6HxVz+MYC8a0Bn
TQHwrnRhXDZ+f3jz45gyIHpF7LLmsKcvlxUP/W50rzXmyBZ417n0UJSDah2UMnIk4z46EI2u9YMw
EIWYDFsmLiBUD/EqceINodDKBORWidvBkxtAkF6FnMdg2/vdSDYGz1acLjTJlhIXj4UX22ZOflB2
wzgH2/rqFTdCcn4xAvmHfjdbhehzxl0VkHP2RnW8qM1khJIZ7FRPdM54NOe63UIunqlmV7hDYZkL
CPHXp6ykzoaqmgQ3vq2RBAp6jKJEdDFETsh+gwlg6p4W+zMX/BFJ8INs/If3j9lGIp9pxlamWCJP
zo8tqAjg0QKPtZbdcy9A0FT5j1PIcVfnLd6y54JRSDQtNIrgOWKgb79CKK6Oo8IsEGhBrkR/h6bN
uC6mcIMfKfVXQEoO6bGsp0FwHgAq5MaJpVE1gypQGF885kDBC0RjJq3rDvpIYwXBlhE0CgJSayO6
KEfD9b9AmbKDIL9Vcryii/jQYz40mNaFxqSM3lv2hiodVSPCCxHsQa3peAfWPd1rKjPate0KaqH8
m+b64IPnZEy6B/CXbYCy/1Qnzkz0HYOiNFwiiDshI2FNMvW2kyu8V9uBgFc+D8y2E+d+rOP/vavp
FjcLh71XLnX+Zlrt5V5jNDaN/LKMl0rnpsXDL6PzLdUKTG773ACIdXVkg4cKWe5f8YxBPHnwseZE
4glY1fQ0RtVM7UyIzrVbRlcGJ0UD9UN2c4QPn7A59qxBiKipf18nG4OMq3hD6JgBIm+7Q9wmnnzD
+CBzocfe9SDT5EMrLydinjJyfjz/hlfmKHnXmxhdX9YMNIMlnVCtd5YKJjmlYDSLNfAlRknXfH33
D5Ee7QtSYll82bKpBIcdXl37KBWNwDItu6E2qVkks7SEKg6J6cZfKs2UTl2aMxpe/GsFAUwiX6mZ
Sn2JhakHbYIuZcH+N1u8JWoNHRIAwAe7m4YNq4eTzkhw0/h33uQ2iWQNbtitMmiBJN/Roa69lA6I
PvXVKwZ9he7edDkcYwZbF2KY9znq4/rdzpfyq8YUiGQ/f/pgQsY0drliopqL+ifeFO4YZ9GocY9k
B16XjE5E793TZysJOk6gxsZJ1rDxO3XG3Lx4WGrLbta5peLwRfq6vjeZ7zh3mo1QBL5FLVTJXC6x
flrFweac6tXNB4OQUSqPZgr7J/F8a11LZml486Oa4rZ0xifH5PkKu4R9NOu0f9IoexQ9XIUHoDpG
8vA+JsBYgL/lNr6jWqkNIPB3NRrXAmZUHxp947VVBYcdwGxpiuTv/MZeMp7Ivtc8R6etyqV4D+R+
QR5kBG6U+wX/r7dpn9yKfLl99wjAUarqQC9NzqDjzAN94CmBFByRy/6oeKVBmPGryFh0WadFcJB/
78I+d4R8XMI6f3KabgX/NoJxQKXxfCPshsv0BgQrn4yCuaVa4/fTIx1GRzsQEDyohhMdQHixflWQ
4B/dK0cZzeV1kllveoRfWZTHI/XWz2MWMVPnFPOK3W4cORVFRYqRG39ze7OvTJc11KQZA9Je1Hr9
/joKtrEv4yuBW13EcpPQsHA0VLsNw01VNFP6BXRV8ywTbfx+Q6ybOcdvl/PTDh3IaakNNM4Fowp3
7Ac8Ns4iPa0NgRj/PjpqiH7GJDu+A3xl+hwPmq/EMJb7WNUVJlXWzp8IoBVDzrJcu59zfaIDhJjM
PLt/Nvy8GqdcJTpqEX2q55KE7UG+Cm2nnSEGanPHgVRFMJbYHZ6Ur4LIUlBHSqOal5XE6s/qkSpS
uN4neTepqbmvY/950d11BBxaINwMNOeg1s3AYkhoErb/CyzkQy2KbTg8nWpejVio+3kJ2UnlN8xb
48hIK+QKXvBHSebxwyQQIMofUnRLZyXD0MHgczBb0C4fBnCqiTSuyvfhFw7rXc1K6OeGxMCqX9+S
x1pDrAPtIuLy9Qdq6pliz7/C70K4I4O0RE8pIIPsH/M12/6UcS7BFSl4ZWpEjkw6OQSTf+VRacTi
z9h2PvLtZuC2R8ogxJ6ZmGBMTku/cp3BEv+V32Tz5+egdJH8V333mzqm63rZXNElWKSr4BN27WGM
ypw1+V8g9pxL13fiy5NK7sCLI25pYKH3FOyrbeQRMy9TCjUId4jkHQA/DymNYXpHC7AinohC11IW
pHj6WBjYssih3DYTCW/c1QB1mRSA7dYzfRPfN6h4jF86rvUFNOdy2WwIe3eDebW+7j31aqEkmHjz
YLZSrDar34hNOL0IDQ8OV4fTT75clDVzpiMd4kxUUyy25RsHK0xvhRBalNAYf+GLNZbykNkxD55O
CE+6fMTTqFEGynZyFagTmeYfuLCqW8DuaErMiCOIDcF/pstKX/nKLyGc8YZUiVIw2MnrIcX4FvdP
4Pcl1T5+MzXpIuZD63Lt3eTvERa4BL/baPNfrdK2xMWA95gO7xLKY0SK7Vp57C7NAX/6tFzn0v+v
rBCWH9eCDIbvymqxY7/cKj2GvFOYw+vEpF/pmdQfMxDV44osYJG8wgeI8XcIatpOpv1LCejE9sq9
PfJ/XGal+5EsHLC32yH8BVSrHzPrByyyQCWOgCoEOsqPjYMnWUDzFio0ysJg2sm2QqyCjgFyqk7f
eZ8ZMI9V0c/F3cpHP1cC2C7cQN13seakK7vBJbAFx2KQUv1D1g+6O3X4HKuLMkRIInOZUUhyZQzC
v/ivmyZ/nlp3sfQ5GNDXdwSGWbUscA3XYalJON5KOMlnKqxRCxXC8PXSFG9trUgEpuEoXZ4zOy8X
WQwKtYDUu2GivbaNN9ATw78MZskaWy3FFQyTj8H7SvqWDx7FxatNN+0IsyF2tKDnoOjxiOZfo4JR
40gdQX+u1SXCOHYNqJRDoHUe592TBS4e/iBxdCVw8JEzioFkEzncI10jUrnKMX8KdWdU9IqLmnDR
wgnS1aSwbarLizd8jpt6J0qndDOvuz+m6lI6S7bg07tskAjdrwHYJrmOW5yxowTvL1lMkHbNJjL6
QZutzipE0l8D9vqEIQ6KY6ni2oKgUEvzoxJQu2Iw7XR1pz3Zacn2OjZoNSJDq/InzxolKFC8nuuz
QiOZMtYaLs7R7YgZ6YB/e6uqkBxAyuRN95au7rLpYz9O97WJGa88F6N+FkXqH5QwjfpUsCbunUoN
GzW0SMSVkLOT4Gl4ld8PyVpRTrIw6wrxD+PKGLMA6g7KKRwRaUBaZJ+qTmkHPFZvveRzEo8Ysdqk
O6zuR84q753QnKws2t/yMb0PmyAY0TobW9iguY1hdJdFUtgk5SB0bKw558Lh12kI/l6vFaJZj4Jc
LEyYBvU20KeAQodv7/dTjQRc8b7Q/xi5trMb47BCeyx/vF+zo+PW4F9MkQYLUinu60t3fFEF5fyt
z5VX2XSXOfqAWe7eVoJXSnf/WbOOr58VemNOfUH1lcz3KVwgSEGgW10ZhSit3RvxAXuT1ORE0x/C
/s8vyBwdByntlhcPMxsj6XgR+eiXE4CMciBtqTGxBVt8fJDWCbimR20TqMouwDwjlUmLtvyBjR8s
qKNaWdXdUS/MSNEjpg1k2XViyqAaz4VBSmVlkj50gey8MPJLHhTmskW4MD2s7s19xae31+SaQF8D
Ri4niLqRswX4qRsetPgA4PL1+dl8f2NQZ/N2j0Xd+YVmzwgyUeG1lElqf2bZ07Lk0AMHTvXM/zoA
SRIE8XoCW6cPYc/1PvbhEZPamTJUbkygH2X0WxVncLIhMHzzWV4jndb7wOkWh7CMhAw2HRyAb/Dh
XT3tUyj22MwSliH7Cx29OETbo7hZ1/H3hRSgsmF1DqIafkN+pPuC+UrtTURLQg6H4kLorZhxDIku
VSmWkwooL1720R/1EJAOiw7bZtv8AkJ0YKB0VZ1IzmTXOWg/x9RspHDVWc0uEJPrLOVrFHd6y3wj
L+WzWi35SOVu8KZ75PeZ7UG/d+PDxVgqy6aOkOtckR9HLCYvKAWvJq+E1F8RxgQ0LN7v6xRu1V/f
jpzYxxEWNQHKBv6b18pazWaKMeRIvO5O0lkYYtSkkbY/XBCfhedDGJkOUVu6mhQzVbME6sN9uhmk
3hStvdNXsbVWrPEYuAVN8j7QjK0IGr3TNFRcn0TbAFoDQ9/3sVtDoysgs8cc0h1BNDjToU60W/Xa
aTvqGtbQvQKnPahUUylQEl4WyXiUyw15Kobiq0iUXAVsg12KiccIBuLjzp45PKnYNKzqXs0z4D1L
OFi1qrqAIJaev9D+BBdR7kAoz/BVSQV6zQFUMsWaA4zloOXIGAqBt1l/azijY3k3k+m8yX9wlz/T
a6pKEvcei8Av6FaR/RF0WCBfY32l2F0iRh397OA18gTvq9KngKuUtOAoOzcTsG8ElKUh6zjN2Fuj
zJYvO0V4VzIZUYK9S5AxohSxNosKmxdeqcO7eR8RjB113VjqLQxU0Bu3c6WwmGCvEpsktDuoPzod
v4AdijZcfQdlHvzgOl/ZstsChNXnLh5dlejaIxgBj6X6Y4vsEXZFfBiknAOplN4OxP3TI7K9XNz8
bhXYpnSQmvq1t24rdm4WbArmWPdmg1G8jQC+HC8tbsD/gpfS9XCTYFn9yslaXFSouGKAqLeT8h7n
i1j63Rh8X/hj8+lgACs5G+nOUSD89FtpMXO9DsEbtYtffjz+psCCT30v1+puCaZ+O1rG1nvtrkkn
knnU8eSpu9bQl5E49nFQDIicsGE+vwPU/PdTerD5bpVREn8aLAhbGHK09e4MvCElPUf0v8UwXNrQ
jHB7YMpmZL3pYNLPxVzIHDC1z0EQ4OkkLDVgyUwiezJ6nYhpC0UqLOWOx+8yGMqsTi/LZlX3maV9
RM8Hl7AmfGedSY6J5azBtfEJQ0acENzVA3A28Ngyb8zOoF3kesbpWFnTep8L0nBv5KMMNdRH2JFn
7wYFAk1pXSr7OxEkWNlWKOnuyFMWDaba/DNlpWOZ2bNBkggaBpFZy2FMs7QqmGkU5WWqHUDSb3z2
LPPc6XtOrmx5am0h1f+LLgbqx9jnM+/dEbQ9LYEixv/PnDdzRs3KfKAkH/KK+ZWuQxbk9GXFAcQh
AoCQsprWSoVsX1Il8ZThRWlnEbN/pKVvIsI/YvFXS7f/Q0F59A4W0E9MlnvzSM1NJD31G4i2LlwS
Wnq3sIyloCR99ojyV/gQ7aDmbHXLN/mgvGznymz+X1JHq5K/3MqVNvY47MVS6Q5ONyvVRQHF6thT
8/nvtwUfHeT92AqbLJzHQUK2DgNwcQYa0z6aMFJkapOlUS1bKN2Qxw1rPBlFwiz3cjbaEVAEgxiQ
koBwLZDh02PqUUzY0kj5V0i59PKNBjVzffyDNJfZ99L/qV2CHDgobjp2hfgrmuVnyMpDdwvG+0LG
uPRHaTMCic+YOsTyB9v23TjAiuyqz0krHeKqRvXPi68o6G4kb3KXs07NFMgBGpuy2GZ0I4NXTO2X
7nJ3KrDxYiYe5sgrnlNqRdsY2JPus0v5owzDokUSlLyO7GgvS1fU/jSv5UIaBlj1e815fTgCi/VW
dBn2cih7UkSARtZG7f0DezEw8RKstt233OMQ/paUgez1n+ieNu9lOQdlYzjYWdFvkpvBlyxzBgys
xYc0HcQHge+m7LE8MAtRb9OTGODwl1L+njnNCbv1/mHtqdVKUfUkK9vuZtC+PijOZV+mx9aNwZGY
g3CVKXa71/SOrEamLdu3BCAvwOyYrW7rND9eK7gTc/chG6fl7h6pCkNvMaV07+RyfMy+6boGMsTz
YD2lopZUlXfGECK+Pkj/JoRLTOBcNHuBh/3yPeFXCKQr3LJUb/WQCz+4HFskLRfHWjsDA7VdlW4t
d/gtL3dV+HAsLakHML2ezTSI0Clemm1O/hkanw6cKrILnZP8spnf3iOTMWrA2VH/Zc7gkWty1Fkm
XQwKvVea5SddN+5mkPdMj4wTvx90HPrgPH614xNwXkGlpLQ+dkLYrk+mXkgyizO0N/2MxznBECiW
6CqflcJU1nTyf70fAdnxxlkw2juSa62yr2c10gmIph2hj7hGlP2SM3p/tIjjFeGeGt56TV+mNW5c
BVXWzqPKdu0kFkZG+WuchmDdqkld+O97SFTj6uui70/bzFVQQWjUsl3XoFWFMr4ix8HkMfHCtXRV
CcAabUMroDwLw+WaGVkxIRFdmeD7+TjOGUB8JKTu/HP1KQDCGnMslEqKy2EsyRCkYyQzcd5lUOX3
TpCvtw/Pkzz7iZUY7LXr3LD+qf70S40gNSVB/sE1iiFVr1YddstWefSEd2dXHd4QbIv+dvAaIEGn
biD0LrS63DFYI5IJIkObquejBmD+EstCFZAHj1KhYr62+iMtUn1ozvqz9Po/GA+s2yqq2dDc7Q9k
TxME56t4s/Fe9FH4slkTTQRBjCVu8jywJSBh5kNluZQihP4NSq7D4j3DCDtmBHOKdSH/SmWwzjTB
lFU80bqlW5PewiLeYAJsbxVf/VBNZk82ogoelfRgXbtWVSTQu6H1S/3RuLdFBLdZ0kNUOIluopgc
3W9wTMJWE68gU09x7YzNIxMEJGDUlTbBJ7Ip9P9CXMYHlnRPCuuRRb2G1WwRpL4IJDhtg0Q3hgGg
pa1KWBdhDQ22LSAceW/onuwT6sTJiP7yzsCoFSG5fTKvteyNEqaz6bKepluzEvQfMLe95+1+BUpL
iwNRbj/JZDXvjG5ZhohTyZ4M8ph+uR15dLug3hZJxAbHbLH1PLeaaBcnPY6vlAmHhSpsXn+q/KJs
sxwb+gtMaVTWINpau23Z9F8Mp4iYUuvEUNmuG+5/hHgUHleUgjfIULqXn/TjIg2POHri0hV/3D+Q
Uqf3G7MdfUYnVla2JYful9449dAcE7U0QUHpEiKjCKfl5c62yhlAERURCHCaQdE8arxNwFPsETaE
oqolKInm6P15bXAge7HGUgPKvM10Zosl6Qs0hyBvfgGzXmR3TqdX8QMDUfZEyH2gAGsTWxcmhovl
pOa2pCTUTfmMdx0N7cDLYkX9D3JjcOl+Ye7m1/1Ss3uu5vMxopSaG2+igCley0dr/MGifppdH3kG
KYPWfDDvfKI10Wfp7rfJy2+ZYbwIZTKPkap0PbKi7ht7zfBaX1l+aN13O3DrcW1J8LouM8Z6VILP
9BLM2Pf1eL7i27IBIC7MylxmoG/3SOLLOy8l9buM3B/oTBkl81aVTHcXLxCHfKZskIDj7Ge3iiCh
joELMLRQZW6JH7KfnbiyuAfGZKa0Gteag0vVGx12+EEyUBJ+q2CLjKuMfwnxNCocZRDWE5RyLhq3
IQrZTdguFGdXHCNXjB5gJcXtoIWEtn4p/Q9LZgUwQR3Iay6MwIbt283UoamiG60E9MpL2lVkvtDf
a0gopZbMyEB5hYXvIvJnDMIVekcA+cIpea2xz6DSK/V+zq+awimw/7elDT4TODFllaywEqMYvA5X
8DDQfqrpiZqn6LyaXJBVnmn8ykEVCrfjvWrClLgHuUe7pcgmRk+n05+LF4wk0xD9MjysOqcCHwDB
+R8vA4rcBBc0EAg9iaSSqanG2oSzJKTRmITS4bM067BkL8GD9PWOutpjY3+hoscCKYnbHcJ9JO7M
pyOdMaSiwikk/Dvtc5oXyoOQ3R8XFhvqqNpHbzyuzknNcuDKFD3ZC3lKJqsEmSrdduPSIL5J0sIY
0xNmYjSvndymLa6l5DzQgPVByljWtpqyA5oiSK8TI9git1yHtmTyeaWAJH4ahZ5/jD2M3LqyzXf1
WBge8agfN8ek43vzOcLajEmugv/dNvEFU3KdOdbFRitw0O0DwkhnGM73Ly/U5BtTM48k9MfMw372
STGRWIwo3OjHcWCSIKHwjh1+UNejldgJswscKTeamvdgR12ajdtbjbKfve7PU96I2a/iqsXJFihX
TtG3UJUb9bPts4VN11QixxunSLQrVsDX/v82hkwLpb1sVLm9sPBM7KnPhuExcr2Vxn9EUw6lECMy
c3oWlajvAjUL8zKXDRwolON31ztr0tZrjOIb/UJk7Oo3VE1EZZw61pBn72agknkJDZqddDz0M+aT
ZdT/Ls8BxJYDJwPq3od+qICK4BjZnLe5VcwI4jTqpJwGpi1GjkXqf0+4880L7c0fq7e1vUYzPMTR
T2uQaM8cJP0c1UTVSCMr7xnp6nj/nedYF+c86zOWXQoMdlsAmeHHJsKpJRiTwWyYMu198ihSAyXK
0N2Km5c0/zyW+uYbvEmZNX+s4ZEYASCeCTkyM+qsENs8pn6MAaBZoOz59ORqq+0NTIbn2BV80lND
sVSiSU8A7RZ/sHd/i4Tlw2ZWqxWChOfaTm/xStapKrTpTbR9zUC83b6SbLkpsSJaU6ppgrOjnvAB
QeyhKEuOG7aBrqKOvq0LnMwD12yz3epUpv8VSmQku6ExZAW6daWcnQkHoi1HIuEffJ6ZTogGdVGz
gT0HNsIvEbGb42woJbnf0BQWb1nwEdQxeM/pJ/7f7f9emMS0vXBCLnGdvkxQoiUpzyV7+HVF2vGf
n3K4yRBpH52bFbbJcJ4z6GE0PNYIShl2MmdafDLbp0bOPCMYXO27pttLEt+gPl/14aOGlo27rr88
dCJ12Tt+a28IjbpT/YPeVn5dGAlTObvxrIx4cpLIKPCCyOgwomQ2qfecU8tcDAzQbihufnP+w63J
T/Vo3xjmEf7qQpHWLZSC3K/Q7hNLcDxLflSMMKC9l818z3GVlNR/Nu4Za1zuZp8be1TUSl02Pqt7
5YHEy4GyitBxukyiZ4dc26bH8J+0derLZ05hqTrkXtRt7W/Q16ta7Uq0Llz+tWRKdJvJPsNJ1l1f
ulUcpG/Bfpo2wpVKJbQzqur7SJZP0EAX2VKLkkBG1RDud7o1goB3OAnRLhcu9+Uctsev9MZdvUxc
E35R81qUNtZ/Wrv6B2EWHLTytlP04jXd88SB23Y8KCQS5CF+PbtxpbPfv7YMAx6BSWiQfg6rgJyQ
RXAdkYNlrfmUSI4VjnDOd8Pd2fTMReALH1Vo7EAKAZdVU5/+Jn3FYI+kZbf2zEmnMZuwjwWOpGL8
QMk8gfIbEiRFvaBQ2g+9/C66aFn5/64MnXjqtChTUYzGJV+fAkrvqCrla7dm6UGnC30vNi4L1zlo
dC+EcZPQP0TY/9s8MScgJGnqCEeytiGy56H6s2xXSc5ZJhfgl4AVCaYejgbsYMSBjwh4f/ZqgnPu
NEX1pikFJoM65yrZ+UiIVoX3sPQgRP8i+yDF2ZE2xOu9u0s4UsBNUqu9T5qk1wWBbjB+5tZWyJ4T
x/OuyrfjZ2VgW+RILAX9LwwqVF5/B8rXx0sfaQZT6Pgz2JdQMMK9J2pR2JTf3cvvkEUwqTQbnygY
i8mNhplREffyl2y8cAxAks8OLVZ+4//9rB9tFJX3+s8NPnHNLPPs0JidLq7qwTdheT5A4oG7BtAj
btbL3ZFiCpHtbrApvltVnTxprxOZyWnyUC3e4HfdwPueMm70COdLzfMVI+rPIQcIpCrTkQXQa/pc
OkTX1LfJvF3B39AkEaVQ+IEBNOJnl/sDhw9ETYNACC2qh+J/uk3+YMr/6bk4klDALEuSrl8nsmXk
jiBLlYq64NEf7g3zAZinQY48zxkarae7Tl535aG5EKJsn4C5i3j/F8h+gizT1UTZgu0qbnzwDB0p
A6M20xrf/FcVOowCo3iWCEL8uxLQumHLT0/w58vuVWBiOtsvbhstTzlmg99lx3Ylrd0DA6FofigR
4hoZ5/82fgwNTHAp3XgKou0PkC6LB4UDyu3RWdPqT8CDmRw13bh2mLfe7nu3PEFUu8gMLNlvcEnK
pDgdHQEakUMs2JP5QZtVrJ7coAfS/Pzu0nlBrfXlT/3Vw3wiA1R4rHTqjoIK+BiCjAiy/HJzkWCZ
ftoiMkMUQLdGQqI1wwiA7QYE4N75h4AnZ9aO6NsGtvhnNzKgKEmyMUzsb6nf4EGVY8HIg9lYuAe4
BIx4VkE4VItoavvZghMMhsQh4im1jso5gkCaP/Rz9BZUdCL7S9TiLmf4f+e2g/oMFLQcQLaK2X9K
CkNoCxEQPpPGtOENi/ifP0onlRlej4Cc5gHD4Gq5GG6g7cjfXXbo10b/2DonkRDks2qtQWMRXFcQ
6D4Lbh1Y56p+buJXdnE35dYgmyGFVmv4y9qPQ95C53t0oJd42uEXFzHbAikXFW8VV2wN6RlXDzNz
Uzg7diXYjy1c/ZIyp6S0ZVA7wq4MEEsVt63pKBYEzXEBpZTBbGYL+WCRoqehv7XJvfyI8pVI1Ojc
UTP6kUNu1YSo8LFIvMSuU3G+dCaLkOy+51sg7eJia5jwSs8UZwF9fjUcq+OrNWcVhkNzYFAInSuM
sBoFlGmQC5zkwwidC9fZj7nVXe7VNB6eyOxIObaj7V72AoxBlXmQvGnjbWXk6sw59Dst1ITlvGI/
SL0Uo1aV6y0mdG+XJQ/Nbct4SrTfn4rQ4JDkkx9e9uty3bfxx7lEHxNJyztKBD+IWhGKoLO1vY/Z
KgTVgE3VPU7yM06AnscfJPwMtoVhp7Jv/ZkXgfid2pdhBuec0fzLmCWuxmkD3nGG0Z8PE6dY8Fdt
XNPrEYhUePbdlZO3KkKcKThPHn4snISO83Ambgmf02FTbyfgBkaohmdFS6OqaQWccYQF+1MjBjoL
w7yDZFC3+2G4yZoHF9+Je3HtH3qpjJBLO3bbum1LXq41RxLIRmWq4i7rx2e73Q+2ccBxuuFUYqH9
3OwOTs2l7zcI9+OQrnzxFkCZkuzH+DvLwgpq0335PAcF2ctILjIh/jmRezIrodGxymOONS4w1neA
ib6nWFBZFfJVUP1wLH3CwJk7RrW/6Hy96thHW5+rTyZFNtZ+1TvHpB2+300o8c9NJHAdjkYP2gQW
0/n7Za9OzZQS4cZg2zh1fvfHVozoQy609NT/wOFRlhFxgPKrBGmkcVbtE30bjtVzudOzp94zGuMx
61mNB0GeE5VGA79FRFsnE4Iv/QggCDAbv9agGP8rAYFS83hRo0N///ScAYLnNZGshgucMFNvdMPS
iXHkioHDSt5lw15yEq1TO3uz5Rax9byZ3N8btIvvqH5/qyPC0aJKmye0U3ps/+EtxxyiD/bc0CKN
gWKfvg7IuKBSZ96gQ7tcIGn30JRJPNXraHN8F3ktokRkkWEaH1dkpV93QLW6frhqkjtmyQ/lojXP
0fanKdOVhtuU3cVMRaHMg3NAv5yEzjVbW6F1TN/rYYBfXwiavzuD4716g55zIR0P5NxipQ66g28g
BaAhj96eFqBDN5VknyGnVJMM/CcaZcRd45mvuPyj/DM8vvBowIvRbEoUY5s+A6PcESOrS0F5Sbv9
rt7S9vvlQyl+0/GMmk3+wnmtM+Qs9a/UzIN8z6MZXktPboajqAnXYxdaBfJw3GxeplVW7Ia6TqML
47P+g2F8lEQeQUJHvGSG/Dpgz4jHyfZjJikXPbGfT0rNcsWMI1f4YUpWZ2DPRGL+4ReuppgXHxgY
jFqXO8nHn2iPbhlqxmbCO4aAqnlF6KaCyiZ6Kta0NYP3hCgn6Fl4FjZySObyF1s9W5NA7UktBNqf
sY3aw6W1PMnPwKjPYZkokjUBSH3gzbZllUnZaWeH8WlRayMGq7/41LOnS9pR8qIUZQZy425Epol9
BAOJ5TRMBro10HaQXPS3hrEmaB9VY65PNQL0+bjisG0XnmLlCv6utTi8efdPfguOGO1Ictu4qi+o
RF4aLaifCFJokjglkxKy0qXEqQinw3hkg6igoJWvxO6tZ+yZHkmsrGOlXqOhq8fF0RGwUVHj7JwK
jqhY9roMgcxn7tNrRlNr0AWmU/XSbgRy/PCdHOKpNkPa9UQYpGWiAWPJyyMXAtwHKMzGS0Q9MUfo
TBWwzIHFHtWFf0Gni2XgLkKMEY2d+IBxflxljAZqAERdj+xNjTztabP01iYUCLVUz4XLhv9Etge0
E95o5hk89XqH9BjqduejOrFPwnLOr+81yR906tRq/NURvikE88eGvC3H0c45CST7sHmLB4iBL7dK
4pMg367/K5Zzkkaf53r9AKsDNiMAwOZwvpiNXhgB48iuU0PuG9+h5mP9bKpIFPmznb5zv4knV6Sj
BpIXTOD+UH0MixYK9xUlzbgKTdWRXMENYWRBsYYGBJxBIFKIn+rLVsYYoidTiA2LEu/sGBJhpEtW
/UxkGaBIFPn76otzcbwH/3hGMUBl2ElrXHR3fp5gZXb3hfmmMRc8zPGE0v0uNvPfY5H/L14Csd/s
xuX9MPiIfysQhEUaTaJIlQhNHULPH6bX98Lpyh73Z9hRRUjSZm+miyIQfFnHtGqb4L4NRLfzs9vf
Gt/9OEfoJQRBzeJPN7xNMwA/fSBIbH749C2gTrFM8Xko+zsYxREvM+cczsbg8F+mr+z8AeHVkES1
I6cEco1c2qNuFs73t0bQFSoD/JKBa7OfWR1p6dkCFVUgLcnJTZLX5FA6P7dbo8Nqm6LXY3MhVVhD
x6j7v6FVwSUUHAKUo2+fwcsO0smlBDTg6/F0VfY+ClPMVDicNpjmFJYdNRCUonkgXWAUxl14f8Y5
ozk5v40Dkgd0UuQDR8DW2qyNKkq4rwR3tG7ABjiOOBQJ8wD8Np4Ggf+RtXY5LbvkhyIDCJW+I4yF
2thdU0yAqrH9VaJP3nVz3jv6JM0nm8X1rg/ioFz1KOnPfgLQ3y3kJ2BGIa0NScBaCq845owOHREe
q8BVg0YovSaaFXn5OWFMyYtN6caFn0G9BWtKnhxnS8ehKstpN2mjUof0WAO7jWzMZVsjN+YK+rFq
ZBPh4fmRbNPit4dUe49Ce7OV/YUD5+FOiJFYUbnAPa68U5t+3cqnYzPDaVEwinQVk8QEfl+HdaZW
0RUUAJvi0FtpFIQqdtQM8WFjuGTGtDToWPOmr7pb0ZoDGxUxw+x4pY1mRVc1JDr+GK3Neq2eP8CL
n6w1m57JVIN3hI7rWsrpftHUptACGahm9sudcCqgxXvi+3ltQFAc5lBFZLZGuB0nPXNRduhvvmRf
8JU+z8SV8M4jWTpL7OCmxjdUF7uYEROwIKKcWf4f6sCuHE/hor+DWeWvzXHlXBO/qFnX1yhj+cpy
D6Fa8hAjIaxlvQfMkmAi7BQlV21febfpSQx5L7YF4UsnD51LjtcsgOOy0O5emkdZOuLFA21KYtLK
8lbzZXIdqOldfzjNBmAV1l8nlWV5K6yShp9JP7WSHjnBN1/k869ZSl4clHJdYQvbfQqYhaOqmQmu
NGX/dtR4QFY3tJyvm0fAdVieZvY/gxVAQ/Y630u4Cgvgmj+ptG42dvYg2wFAm+NAdMkW30OyyLLx
E2NgCLATaXFUw7gjrjB9k+a1hk4fyaHr2WsbrYt6q7uW1h/0/h0BtQlmaasxViP3PFTrUxu2jzzm
66K3wyAYASKamUs/NuV6cz5+MXfW+VF0/nYQtW4IGglt8hUA/RqSdragH1nldpy9/n8YbXdlnDTP
8quXlTYVNAFWcYJHTiG7Ls8hc5wQMxOs9DM28X4i+PT9Rpsmkdug6KPdKnCqC5Q0QNd7m7zgKe2B
5CK+r6A8M2TaC87Nxm707q1ng41GmNVI1CJiUrxu0sIRI+sNAboKWvx5COD0UqksNrmQLh0DCmRW
YxLsdZF4tbI3wJTzcaeA4Y7kTMItWQCH2IC/9FMlDqgzkbVhnlb9hr7StxILhOg982FRiG/L6IYY
RuQQJv0huFGovJQO+0qsEREVXWobZO2T55DS37rKfmIgYvSKASVgVJA45KSS4zbzProX2ggaNhfI
IW6ayODrFtx4N0/bPN9rn22+oGmeSj8NZ5JHqLB65QbLt7Yhvu2SiNRso3ED1NKhDUNVs5Zvqo6q
m6LUz0yRvVzl7R3+Y3HRAeuMhjsz18zlYBqEyuvcXFc5KMZTcoGZbrsnUZOlsTIqKDlb4os9xVm5
6ng7bW1EJWChXXh+shP8bQ58vB3sMTdYSpXKSFcOMEBz+F4fL32GR74QRcHsD2kHxRtNBXOf3o+K
XB1o8dcD28LryEJu9sPknjjEhEp5ZeQ0t/NrIJzh0HKo4kXbxhO63CWwdIXb/wwG7PBqqamj0lU3
lLcNhWe0WvMxMYPuCHv+meIPGpxS82yRvf6ypj7XkFqfLgylnLbTp0ZBi9uh7lK+j9SvwBOomrgH
3yW+mhF8R15tavy3p0Wt1OkuLKS62ciXA/jrxv0PWCcZltfmLlIppSRPUcuoKER8qeeSkL1Ejp1R
VM3BxLs2UutycXQm8rVI04bTTOPeQSS4MvZEGX5Ylxab3IFisMs/BSxZ0geO7OZLii0EWJq3KEOo
3zWSZTmuREHldH52Mg4IjXKxHb5QD9XfbelHy7QAPO0ngOFkSzyMTk/B6vOVSfDO5B9wrLSpBdRG
9WuzFC56RIVZknHBBO+Do01WYg4EmuyMJEzuih2sKhn9KIcfI74w78iUU3aJpXmdbX4k41/jd8tV
BhCC5AyLZQKDXpaBLKc63OgyQgp/oCl5EYAMmNmB7kdcPbHRubPmlJTSIsLeMU8eeoAjSvpRaF6U
jmE9TR+pSutH21p84tQgWvmDuvuiSti3Q7qA81pmzlFEn9kldgSpJAxx4kcF1ePQcfEXWaVU+JvS
3KwIvsmersQUYybOI1JonKs6LX1FUogD8eyTuoDaUphdXdJawTPcYkYUg57iv3U9PV7ULwchpSWz
RrfshTQcZjbgNEWcl7JkbylYFEHdrah82A+kVHb37dw9Ba+6gsjyFMGeY+yW6ekXcNRhSYklw0Cm
/RpmcUu88VdGazab80ig3qw5rYs9jHbp4WfrSOGdDrKuiiKzwsg+4heL/KNjhyIoA5Dod38QLUQJ
KzOWFDgWF76fA7prl1oGMMioACXZoiln+1s8w8D6PGUxKFpiLnC7X3z6QKW/ryKi3LjJBgEyr2mG
OHilFhTFMfbrvzFTt7PtFT87Spd3yQ3/so3EaKt7ze9p8SX1o2opaiPSv6jU+yaTXZa+5pLcYred
knT5cCMFoJTKsziurlUOI8noU/rsUUJVCDJ/skDyPtn3fGfE/uzO85nkckwTt/JrE92rrUmMR2Bv
widO4d3qjHvMrNny6TTr0009nizsAMRKrMKdzS+SFUU68DFXRjTtIXqpG+SmRakx/xXFC+1hIsrw
y8KVtWP6g2jAz1RJdik/lqFvgV/hF5QDjOsE0vDO2hU7kknU2Gq8hCwHuog9r4B1Sl49DGt3bJLF
7l9feNzZxQXORcndIPTunXyWkbuckoRzGPvvbmAAEagHRYttpe7c1lvK+ksMCxPAcaBBl6uwOi5b
QDAPRl8ahtfcIyARdloHEp4VMsG/y9cFqPNfd+Z8Cs5ZC2NtnCgI5zLBv9Snjqp70JAzWiZ6vjhs
0BTVNFCHm+AV3C0/bfkkkMezcK7BkLHmfgAoJqCz1r92rFn3tUcWebbPyyEoK2qHFD5cuRwncO+a
iWKKv6lkg8wQ5phP9VWSfOqFyymkDZYq4sAUo+oX4IXCF/N6/gF22uKa+HzNbdph1NbXjI2AB6lK
z7/AqWakpJV5PuIzqb+w6UHAt0ECutQcL/tpQj3f5hScEFoputsyUfdm2v1qAbW0iElp8DbwcTD9
mzyidtoB0OfwOR3fhlU3c+BhgdgE03ilgwxrMEP1oeR0qMlumsg9Wx6yZqUUjuT/vSbtvMrMOMMf
OCrv9JqnlBlBJblCCJU63MF5v00j0Srlb+3KbFdaxR5wk6WRfRCbC99/AA1GOmysnXbCHL7kXvIQ
yoe3pmJTv3LcLFLpM20Al3N8thINpidrYJIamK/4vZujMO58C5G1aCCtEi8HiEfmi6pcnB4qWkjM
rhKiIRbHpm9B8DXcgFMUql3TcpPVV+I9l3897dKhF3pnoVOef16BzZxkr2rY5CiKVruVoMM7SgR5
6IE/2qtdL/KPgfWP5r5EjThQz9R8bKY5aL4h3g3aSZc3ctr7FvGFuYfk3f/plhWVMG0J+B4Oy0wc
mtA3eXRyhUs1ED4lYAjsIW9VfPZ0ONImSGDsAZH4RAdzUfn0j590vd5WLWFjMvrN7jEd7mVmqrxu
r1VEERJdO7Of5n0WROxP7lbtkLGfFXnAKeeT0oxs+Ox9N24UrFG9ucLW7qaVyicf+PqeYXqhOXCT
x8XSHPHgxrUE7Z53QtLGfbyT8woIOtA9YpRZM472hnIB+YQCWarTqTv7kio7FEMQcC6ruT4amRGZ
mMxlk3lQ10ASUMntguV8nTTnQ021FAiqbYAAJcH0to5+V+9Xq0lKhGECEp1Q3Hwdj1HKFe4E68aT
vZaZDVT+IR1uB1y8BnLGJg65BBGKL3Wa7ve7r0kenRm776DxOhhMvKnmWjkp7o4bbcaoISo+UYq3
T19/e24XdfkFTcakCtiHp2ZVXLAJHPLOoOZZkUwEdaZcTrCwluQOLJWbuHsK1Q5Xye0q2+GSJivw
uQuva9XEKP0Tlpv2nE7IHHQKwJGQE2mD5qER6JPyBpDKJPAr+eqBH8ioZ4hSmxHcVbBlcW2n+Wk/
KSrbnx1iqD9FNrDkVBRuvCwElVV9uBtlXJ/uEQ9TkJtk+wDkMlHQ5Lt55vSDRuapXz8Ifgn07srJ
I0BUfOiwAGR6sKvaKPC2TuRKo3AUrieqB+vG+lS4JN/4Rg9lcXDNNkjsCU2gLcYYjFkbb3u1QVaW
bGxrCrSZmN/2cU2L+jceohm7UHK14axdRyasTdDi04A8l3bijrhHZ+hoMjZmPiQ6H2iKua80nnpz
EUSzdLeoq9SVDnnnMe8tI/G4F696hfH/1T0z7D5iOyPKS3QJju6gkMR1FwXsg5OdKA+ua92GsLet
6q9mOWfIvLeD8FKjQDs4i4rbuxzY2mONBaM3gzScgKpcGy/XdPk78xnRGrCD8Kd7g9bSzSoqeL8E
hBckmb833IKsJcOryy+4B5rDwQnz1esou8yKE7CQbeeXcqYyD3Leda1j9VYvBWBnjsOjX6QmAgyW
Vhw4aX6NJ4Uvz2g/3Rq8RpB+J7mFc0MevXicZ+3x9xvfLmpWzLkgfR2mdraSNhs7c7W5ijbv8oOu
GgGeu4QzfD0gYBRRyt288RFOw3Qx0FW28FenGPM94LxN0itaAnydKwXybYA+PIIgocHA5GVJ4maf
znJudZMt3CVew1XsmKJZ3dRrmu5cPis1Ub/9tbjf6zI9ooEU0m1MzqiRkjFj94PaVXqIhIagkA6b
u7OWP0BmTfV7O1RWXUq/jLFTM2CIg2K86P2jymzu9Cywih5BVpQ3JpW04IAJguC415oVhaHeECmZ
iXv2CnsXi+PYD5j9ALmW32lIuSyXpeMF3JTkq+HR/rst5/sTNTd8auHobhVd0dpdA3qqh4bhwqhs
g21cOHiyigogfMhua4MEyvHiEjsChLsQjYtSuZihoyFExaz+E4aJmp5mgyOtD988Zx7ijne9kw5Q
HUPU50JjbftZzzDuf5cLkmjxKuKmRRMZ/UtG0q3tpEETqm0OA3R9tHmqKo2lJP7M1WoFR6zAorWP
DOd47aZPRGnn62yj/AZd8lJ+122nXwBy7xT7SeOxWAKn0UL7RiVNjnJLUiEyiw8qD+KWe59qr2By
Wd6fExKzv2f3f9ZhCdulyOCnR0M3XnOxhDYGcROGlHvW70x2mDoQfQmrKoyIg+VbL0vsFLtEiw7C
ui8WlmPXBm1wk9tWlPp8/qZ9G3Y8DDyNUMPXGsmdhyPzlb81BCyOiaoE5r2hIv+1EOAnK3qKG/M9
fygEvKjrgikUx+O7vo73pG3slwZnQrJBCEMHEkWqI0X2I1UXWmLQ+H3K1omOT30XWO/bshcXFJq5
ch3sOZAf2te4Zrp6wFtT4u8IwRnt8icePFcLrIjIjhI8piuZwALE9S9csm1kByHOLUZn9QcoigC/
mC4yh57phlkidMXUU96g4nFj/XIxMMfaUJ7D3npUredKhhMw3VxHUj+t50Ecg9zzu2cOY6x7JJpe
uqOwI622wqKIubDS+hJdHPKxEvELhs+7FsGbX9QKY9Oi1/wsE31ge/YnMGI2n7T4Ty4ZndhptCOS
X6m5LlfI2HS0r9CVSksQ+dCSNLdG3gk/hIklTMLtRJ9EqeDd1V9NdswXRWWa6mYgOZa0XhJUaeWu
HLp6Sjfx7c3IidmloU8pmR2kgAzlt1uaBV4ZB+jFaNkUfkeSkiw/McNnigSAtcjQ3jWlF52wAUb6
yE6DbBMSTgfkF53y4gU5UjlDSSVOAOu+cRUnqk1p+0zS/hQ/FMR4kX4P5VTisddcakRCjK0F8VkU
IVDYU00r7YcfJ9Dqbf6TDc5r1RQHRoBHzOiiE5U4H1/7nFF2PMwSA/LWYrJUhRUYQp9rd6Vemi1S
fC02cRnyb9aSykglV8caAdlb1jqJUNexiXK4nP4H5wuMXx2SBK1eUEu4C8DpjPJqxYGMV3ZU4wPc
aRVWlcTkjbOpyMT8/3jFjCsOs0/NZAI7AT554QNhyFWlq/9u5M676ae4pPPXbw5VqBspa5VfFtPk
c8JM2UZPjatvCUSGLGiZaJ+3NiWanRK38NV1ipHPXp5pVPfOPTyJHaH6KtMQFHdHayUHu76h4Ywr
IXO8g9laHea2eMaijxiYJMtIbbcpXqMOL2pxc1nBxN1GBrHlRBI34L5o1z5icjzlN3EAPORdrFV0
SKb3ah7ir8LifdXL46BFdsveLcuvlcO33M3WWpl/dSG7TcEQY7HcKa+OWbCq8sWzQlAU+OuN31bV
A8y3nkz8EeSr/lesucMJs5krBB9kRTUcpddZ7yX2WqW0FeW5m1OyxkrYEpaXIsaeAYzlQyuH/KTH
DOcTk4FfLI9WipwPpqzt3ZdGWWMbrgwVOtVyVlkGypnPLWTrLb3RotceVlJHf7Cw/MIwL3WalBc3
vpY4y0jA0eFUM8v8cLYpwAD02YAlaJZz0Z4Oi080f3xCbpB+pPSSv6rSsVgCAak7Y7IEiscCEzz8
W1UMab1BLZc6c30GYGPLXV3NOtmU8hbcu7tkJstOIxah94a6s8mGs1noK6ANlc92Hd6f1W8EG5hw
XcqJy1KIbFqPlkyVGssMxaXgeRwutT72WFPeoXBU9GvsqcFVeMuJvOMAGuc0NK0q32ANeaHOo6cQ
CcZZCM7y3K7puBR8IFROcBoPFUC7Udc0PUFSAnI7SufvMVeKhFGbBrmgBVJ9XoXAMDhfFXPHGB8y
vqiKAdpZi33PVaO6tywOs1WcOZ2Fnj3nLRqdtEQF08tuydcvTVvtr1WQH5dhZZJu8adzfxA7RhvC
tNKhN/BEpTjj6pkihbZciFwHdLcvfkZNQzEWwwk6Nbj1fTnx4fKOcOUSZLLmqyPnOdrUMOlcbQeg
SIiNKcVYI4npJMSww6HxWbGGcRfPFZ5iYI8ZoT6RZQR5x0RIKCkLpsMAzLJgphk7HIsoMN8qcykw
VGnwlBOaGxE9SF6T5/E67Wjz30SGQK0DifKTBHrKsYFNVL6pwuK/ILjF/j2yy+rmxtRo+CveirGU
OUOorcMKdyXTCUMhhNkXdtwzdaVoXp1SVF3D+Db556jG3f8jT7uvVv3/rg80ACPquZOkmRHKGw36
MI2CU/e3/+fgydCJ7jShYTkHyxiHSWyWPttpNwx+YsFXrtos79tWoDQqDqTovhM7Qx2FZ56P/zN4
cDN3vVEAFEP38YUplO0oc8KW3B+ZVeNKAyUGov2ho1VNYLM/sC+Zwe45gBcb3HII/ZgLYn+Irfqw
3vOwSe1daB9y3XBfFPl9/CiEuybvUQL+9NjFZgud16Qe70tLPVRw/hFJfcjTOCRBKj8d15C/ZbJg
P6v5fSQSLA3w9VSwNLnz0cjlXd6Tdzyff0sMhQ81KZlhTa1l+iQm6cuL06O3S83OZuGssCBfzfri
E+23EFTEoMT3M5mnut3v0Tp1Fm3x3J07skuuUxVnNE0U/si5Xo389gfQWp68njoguC8d5Q3UjYlI
C62woAGaAB8a7MLumo1chmv6Mq7rvpJyNLXYKIiW9ySHwz3SvD06KjRUCpLYkY5TAfPnwkxKXhXC
W+WMSXDQrXfeOCQbhxF1rjma72x1mUNdxy7OMDVavRushR9sck6GgG7OY/eLN2XMELVqpQZuBA6m
mrFv4cpUF5ZkvOwRywbXOndKwzryP7KF/WKImxgK4p+Od/eVSaa+ToAoxSdnS+wYWoL4sKCuHdQf
m2oBgrKRQ9laudVHxQojSFddljVCLNteNYpk/Pl4qF+bhbJj3fl0WwytSEGH4XczVyYaz17kk4sn
8+7QNl4Uj9lgwlWZ1sXmQMeDz7pFJ/4YWAQ2jDEVjDgDUqNK30SDpQPPp5MoxL124F9LoXmRaRfT
X44P+EbzM66m9oQvh9r1WTNWqxDh4l9xDeE3Kt/h3ighbP97OIRwOFG/vnZdb9Jp5T97HtO9Q6ID
H4mmSKK4gOKvPcwjlamnZY2rXHVIkszFyBCJpFE+elG/QtSYsoH1QPWBk3ltfvDZNNdwiBOB6a44
gwE0LYcqx8Mg/qTOsSU5F7HMkNVi8D+4a1yYeZNl2NfWXlyG1je3l7ZNOZKqSpIOdD871p4sVRnF
3hNTSZtQiL95oEcTy0jQPNo+0J/hzMylQPBjOskhW2EJIhmwnSrMad3GGmzy20fdJrojly7zelZE
s9teDcEXuBFZwOw6xTDZoMOQz9CMUPinb0Kv5Li3yJMuWgOn4ZY+aEzCnTMwRAI8eKx87MKpWn+D
m2phjt6WJYpAE555u/t1WlMStmNjnyP7P6lmy1E6ee8V6szLvot7wDhFPDKLTxUP7f3T9PFONEgn
8U1zOCq2BW6bjcYM/uDWtEdqC5xfG+dEaP716yUlqNNeO9jIDUXSnEt0FVK9X/gChCfBg+E2knkS
ED/mgBlk71LVa4nbvacbHRxqovY8fiXwf7Y94umjdKyYo1tV4qW+OvrOpzN1hVjt18ucuzdjp+6x
zGuX1/qdjWySCctsAe1mYu38m5mMHymC5H72N29TB7SoVuecpQf3856RfgkelY5eCUNiW3uJBAan
Gnn+Ee/U/ouH8NeNou+TrnD0kAu18qgE8xuc60sWIh9SubvFl9KW0FDq8ycXQm0ZV60AN3IyoE5o
16aKu0h+/orirknOH0ublC+d24LXWSli3LvPnakXaiKPnAodrMrgXdlT0+jKtrsOQcsb+LINrnm3
CiWX6tGibGrqZWsFnLSOiIvWo9pdzxK36xkAARigYd7YvrQdtYNHiKM9KRVrrY+Y5gN6XV8F3iRm
YSyO+6jM2uYpLFUT3KIg0h+VFBU5+vQAQG0L/MhO1O9TfkZGB0oIIqrqBu26bR5fdWPbIz2c9hHz
zbtGiS8yYjVK45U7NukDgjc9Q2riN+cfr47zqDh4sFqU1ZsA/hLiNU1iKMm3wGAYgJbwOfLbZbNc
8YcFEfhCra4J4cUzyF1kpYNoX1DH+XPcpiTH7ZsLUZ42gCdVJSRrZNgmLSrJ411ifseFEuvFiNl8
gb7amx0mMazoGuxPZgeCiyOrAaw+FKOFS3Tt4KONLwgylZDiNOFGtqAbQgBJIjv8JsfSfmlIY/VG
GOyE9BZHrvcihEB8HVbrL6ScT/QoVkYhDZ6lLGewNps7MburgTZuR5ofPBXAAquDc5i24bhdb6vT
L0VutGxOJTbpWlcouOlf1OsJckqcjrhCzLVQL+PPIRR3kgc2jkDdf7cuj1vt9bWcTDTPop209xRb
Q9MN3cU3xG/DX4zPwLssgFf4BVCYRFBZDTsLB3aLyZteS57u8v8th9ltC1H0+C5Y8k1WzINA/b0v
SRK6i1Ek4ZHxJpt/RSihmo0RZRWc3rc6A0Vqk3qlIJFSbs/Ix7DbzSWsgEqCAC/FDSsuaVjAIkQ3
0S1Co4A0MLQpw2ilerONmMf65KsgctF29Gaeym5BrydDtn5/lcmsDhiEXoBBKc0Rn3npplgEt3qo
w/5U0P9TxUZPnSxNsd5jz/+S4i3k/v+1+wPgv5UUC3YD1Le7v4oXTZyt/ErLS68gp+CSaDmmchnu
f14EQg60F3gbW0iFHSTGADmgLAAPPGxcjQa/LR1cIib3U5uN1Vkfep5PX1m7F/9eEhIoiAET89Aw
Ms4cqUurYRxQ+OVNb6IPjA4NXB1o7mSWd6rt59bqP9FlpUNPVUg/YsI8ar2LvnYplfAm3qMXxo2Y
y5CION7GuGqwy3yvcl8h/tmrdyR5O9hxUqv1X0vmlQ8hrOGHoq7pAYOjX3bQqehtZ8yLka5qheYh
uIXnMc19L/vwLvTqT6f5LEaVM5wJKRlItVQRgrE2syy4E7M8Eeci5TjbJ+FaMyx9Mcvjko7S9qgf
dt4Tmu+LWR8gq24gPnVZ59AqiXr+yQCCxp1fJnFlxzqmcvMTVU1gSwKuui17GS9mFVvLKX5gmmCX
aZXe/7MRoc2w1VCaV6uf6t1/dThz65A0CbKdgLuvGIJ6wicMuAXIA0X+MJ8M6hNZ/K48rINKdgX8
T3piQK/wPBSl6hVzkrainWz0FAHYuvZQdgpMj+nDtpd6WF3H46DWkQo27BdB3QpmR3F4DxL0vpb3
sLfJGlyYC+HPtV3O5y0x33L1metyHk1kb8hO3u5XwSVzlSUBtWE+8wVp1fVycenMc/s0m42rowwa
DUEs4fbnT9TqNQQ0OkzlP3hknystN0BxkoSa4tAGw9B61lblL/DORS0mmi4+hI5lldjkZkbOQ0Cj
GHsQa+I0LPYSMI1bisk6VuATgwIZuQ7vZC4/1IVpm/6ABwh/VDdIX0lVCTWwYcoKq2wcjKcvUFzf
7kUgFn72sq4LDu7Y/t9YJX2MdenPzPETDm8gFK7LeRYqFXfPisgACIvSlROFhiQ+zxZ/+DE1nCQA
WV/jEIMMCFt6hmWFThdnf2C/l6T9brZ+4LCEtxTiI0Doq8u9cXdJPRa1wS5oHZ6IQhBnq10t1czc
MKUcKSNOmFBNbIjlz5XgsD+TTiL91h2Sq6Mbl6I+P6rdpFAumLzLNBJ0sC7Ml/e3rmnbd0BFoMKi
EgMeaS6YVGu6dvz8EEn6GGe6AHQeOndCMLdsi+uHXKbU4ad6D4GFwcEDsDAjB5xQPS4KBZzQSP2q
JuXPM7IenLf18DxiutFKHUNaQgL2Sn40WtmmmlvOAvUsz4F+Z0aroel5btOkmjG1Rpwq8bd0J2Rw
bJsfcPuPt94PXskpmkSP5WAN6L4ynXwDQwb9sa+Kig1CoW33A8RhcYO/s2cqge+GOlr5ytBJAfmg
kaTrnqiAr4olClKaiYiv0a1k574iqgRk3qHJKvRX1ppbVahdGQiQoSWhF30DzMmLUCc7SlMIyoeA
numU9Gr/gpRmOimq5Q05hBCGGsUbkvlvxCTewa79uxz0YknyhivMAKp7YurkUHo+zTAEWixNHEDa
CeESqYFK7Vdd2W+OUQDvRgYO98Nynp6SIQbHp5QZXuzzQZ/JGnDUJfShVjVFao6q+bf2fGhQCAWJ
ym7YIwcjEGjNJXCrVicGzxOtB2t8IEGefJQIIQbGivfkL7huJ/3mOniqNAthFFBnuQhVpTQcy0gj
PcnVurzU5rjcYoRckB+XMg4L5tchDUIKL22B/goNeIeQy4OnMWTCqEnvk7MUvNICgcXVvS31urX4
8auQv0qSvO12w2n8lDQ3BM3vliWu6jY63gDOR/0FyvSz6JM88NGlK+PTKC57KI1vqyMpdQCFRQs5
XrUbG664tcRcI5XoCBYXquf8iTPUu6dSpENfHlCPaPQ5znj6MC+SO5LDvS3mVkcsewsbuXI7SoTH
O3MJ83Tph9BfYRa1CX5GxXlHmSoNf1mr0yJ32BgQNWCRuMmEUnuiAM7zKQ1lq0tZZRLSYQMEUCr9
9NBNCiLzM2OzH3ySxif0meuLvoIJC+kWaAjTFQCoPiu4dhIJc4x4gk1X/fq2lkTIikVK5f6Tadna
XO18JHeICdCpgdxkilQDuNDR0XWIPQI4hzE/lyERWM3YZOFFJa5Ujbl0JmxZx/i/HS8zDTyFB0sQ
dI77XBxjKGl7WjnEW39jh7OxxjD0IG2fhNne0b2kGK9ITE5BHR16QADU94cDn8eQMubsBhyog1Qp
NqPHWZPkHgbxH8lzMoFI7VFrBat8qEeCCTyLIKsjDDtBXqUKxf0Fln0vW9fdU8CoQfLh1lN7zYIy
p6rwU90KqrwxJiyPFwvslZo7MYDNio8YGL/xt4KBALY3Pxv+yJyxVmYy4Cl6ZhAzLl/lhZgg5HQU
rkVjMidkMk/JgK1ecR/8Ija5L70yMsKkuxPxU5wkydyyRSBgqhnUEu2o3+QwZeGqoczGh6wSCRE8
6N9IVsej98tyqLka6+lCbQLWFK/XgGvZRV6rrv8g09GEib1tSAo9qi7dOykLdUF3rwbbBSmDYJJe
KJsH5z7U7JDr7Y7esH2IQ4+BbeF4dC4d8+XPaixNoEx0if6wTMC3Q9qjbrdEum6RKAIyCi3BOK2/
k9xRI+cR45wLT9b39XdfZjQNiQphdimkMzH4rrkHDa9//rzU2p13OrQ2jPE15CCJla9Qo3VlAMoJ
to3dajWUzDT5wbBekPn6/1M3YCsQAu7+ruD1VdFLbr1P8qg9VaUwmc/w170zznFbzk2WUFJ4V/RY
mnLxtUBnWtS+YfTiSS2Ite18wXNLb26G6DH5m1pLLHsZonieqnTFMaUwJb94QAdZS43uql9Icsdz
80DPpSUh0jdW6tLySzMT2nPMyapqzpB0/z/6DNqgid/1vaeBAzfa+lixHwTxPnYXjQi5Vpw4HG+g
4me1h0k/Cz7Tlls948WaSMLxdJNX/6qEkljN6YdvEnDwvXUINBSUR5689eUS+V28bTck2MDXQ948
ajGtlKV3fHbo7kPCLmZcfuaRbGVtbkDxroObVyZjtF+DcXwezvebZ8U90T1fpE9b8iL+bVibJqXP
wW78CB72x7NAHCNR6jH9C/Z4xVY0JYSifAknq2BggoqCKio6HzWNcHb/ZOGoArcY4ceuHWSaB+wA
iW7sd2QS8wTC7T+w2fCbreBo/cpHTqWYnDD82Yv7g/uGB55Exn8zCdpK/O0xfAO/w5P3hmJDPvIS
ehN6cshQF6qdWvQCc9LH+a3cik26bfxWdTWfE26T8bqwnFdaAByJSql+aV9M+6SwBh3WXF4KEQ3m
vd2QdRQTfRL7BKdvC6piTJiSF+q7sdExksmu6/yfvXFftbWJkW8ID5t6BZe7xVyR2C+ElnG0c5ti
EDVqcwpu3FoiR3krA2Ru2Qwqs0QgObeNeeL8IcQsDvwHOgV+rXNUkWMY8G+7c/cdhj0wv6gu6oMb
6/RUAshezxa1GhWRqdiNHh7wLb0xadskkYNtx3mtOO9Cw/aLB0YcBQZ4+tAKeyMVeOxfkkstouzr
w/gIjHuEVIUh/tIfUPdCtnGY+GEF9FJijmhL+lxu4eTGUmsTe936yYM78ICMzHsK9QtFeQ4iLAAK
ucqvj/V9t494s/NfKUnUUJd/d+SQsb5IJHuSwalYZP/xhG09bnTv1vJZ1i/AOgb4dNWqKjwo9XC4
x4MQLUdxvvAPY0p9OAGfy4lRIzlBB4aB/ypck1lcepddqC+qEPW/2JVArrrzm0dkvqLho+7nqjxW
/L9uptBif4utDMmvPRtJCj2kSmaOBfv6KRJhGWF1jm8u+MO3lNwBbGV60aJlIqIdvkRIT9xmhHRL
NFP0tylj4GUD54POFUwF/UnioffnRnpLtXx8RZYtUvb72YcW83wiqNB4cB9yjz9UtwFUtiu0X6D+
b/5kflUkDOfE22f0dUIzxXbkuX0yNddR/yP6/5teZHGojxCzf3+bmkn1NvN18AINGHbcVGnvKYvM
dWME7abQqIHWPhXneEOME48LwQHtUN450Y1qCdK0u5ngpsfxl7kri680pLq979bxAYmm9Y9dI2b7
tvlyMQrEYyB18reT25cVWzUwGXzDgZ5lMhJTdUDjzKobNNE1fCfO/DDLK6wxsl7zXLfDtsbtaGbu
fIVf08tM/zvv+/4xV7yk2h3edyUf6b+PGHS40OQShiRckcfiFt23+pM/xDjisIEKuB4NVvuZdtaY
CjlRZz+q2gwuisMvZptNgoV6pDM97B5KM+HeJmkk+/svb53PjpiUAZMyiPPO7b38hOheq9IiVAWj
ED8MA0Kps7EY1RykAT6GC53LvsLZnaCVaEVLTJzB9zT42ZIwWW4U0pM63peHQIGR5D5PIIBUFIjM
19qUCd+z0Me3i31iArEkF6qnBnrTI9T6i5OuJYYafQAEdgZ4SPHxA/IM55Vsfg4I5oaZjanwxSSe
PTo4GO/dIv4B8XtV3VGU0GYnRm71t9wRknAai+xzqAIVvQK4V3PdbHGa88HHuKOLgrpJJGnXzSVt
L3t+J6R19zcWoryznAwAKs/DwXow0BMiG25uF+yECMXWhMWAiX/5IMblEabKE1E7pj7wL0JS8tau
XKnZveVAH37hTzpuQO4IvX/SC3YQqK174UXvzP1EY6au57gZryhXoKS/8y3Sqxb5bt4pivqEd4Zy
FplgtzgLM2h1fLN6PBQedNcNvbpaNutRv9PJdzq1Rdi4qKQTGwJttKPf0fCrkXBNrEZpk49VIN+y
NKkTxBVDkuH2Mgfq6lnxe68JfFdu6Ty4s8YsXVJ01NvKhWlyAZsnk4tacBznOf5pnZ1WPdKM3rdw
EQj4VRFJiVV5jvEmmtNe76uTnG9Rh5Vk5MYyQ1Xe402Ivu2Wcbx5hq2jUWASUXxagdUfg6xc3dUP
A1jxWN1kUxrzQ2U3BnLhTCiLEb90Yzma6u7VYit3cFa11awHfYig/dZbeh+ICxV5MV+7suI/7+pu
gcFrybAj4bb5wugpCTmFLu1FDf+YSBhHPQ1n2PxVLwtytuMYbNy7Un8txJZ715A2BiGJmOa92Kq7
plPHkXqDceHo/b/NYE4otSNohwDAmPnzs836o/TPgGkxZPqGEYtxFEu+T8oXBhiA7ZYdhQ6GrTsH
LpKd+Q9EJHjVJFq/qaW6pRahforA604ukkay47J6oUtpJR0Sfuf50vr8LG52EOvIGZ69FaV6h492
8nWhpE7m3s6vRQiFZK5otwT/AoiwzOqYU+yi8ehqSoxFPGk4MvbeEF6vUsXCc4BEvdEiQF/Tv8PC
F1/BXbjeXDDTZFbKu8FAXSSNwBXjQXmRiSe2jekAhZDY0wip3JIjQxXiTv2IfYZxsskfO9vRnVg/
PwUDaNx+LAB/ysKDrD9kBY6L9s45H5fioN4ZkfC0f993lAehbBWccV6ktd64MiT+AxE/s0qGmkeu
6S3O1ggnRt5D4FNdbB9y/jb8VdyJ9W0W2NW9biMiJ/uK82cgWEn6exL4Sii+IAA0nKbocwVz37uh
v+wnWwWBQvbnDbx6JnWj0/lisuQkpFl/GsDuDN9Y71zf2lR8175C3PdmUu7en2f5/JICiF5yTOVy
my5FsNSXfEYTjkg/fkGQlY1w8PGD+RmzgatgZlJijkYmZlKJEzWc3bYe8jzAAp71IhgtxYNb69yh
KwZCBP9Fb4WQ2emg5uCcSEpGEvXsgpbtuzXSv9A+OzeDrPCGXPdEmwpCyOZyw9+ZaCEQ8wcm9wu8
q8dIneEZD1CqXJhRULmpLhVL0gGB9Le3hpULM+PVAKHxVdMFPIAq2QTKA6lWoby8kyy4jPHPxx2q
vFTkN4cX2073WcQzwsd1urNsZN3dUWWgmn09FU3pmS03lbgr2cEf1rz1BTuQWH+nc7kI+CYXcDGs
6Tv7/XmeE7reFa630cYgRby337sk9J8IIGWO9PqznEWCDl/qVdiIgVKvRM3s8ctyzLoDE25h/ths
vKjfvnXfYwbOiNFPC93c98Ld7uauBe6BKB5QF3tbvgKzyrfFz98vreKOZKtRc+p2idOfVIdFmQk6
y06GtznfT/PNJaBJIv6i1r14DZJMf70+65j4iulJjwjbfN8yMrIduLFLVeSOCtBXYiOR4hbwAPEH
PrxmdqruBQA2WviCVsyVbKXB8PCdgSaMdeIC1dDfOXwTcyukNkX6AihymXOZLPfbMUZ7JiXLpl8O
VeCPq4t0i91JhHoOMjN/87Cb/yr7kzQ/kheDsnTdwPYC3v0E8XoVMbo41GViFPtKSCAyqctFjC7d
HUaZtzkURsnq3avOhf6vrxruawDhRtn/FXWLpuiR5LaaaqrQ74AfVWAOAfIOSdj84RIkLk/WIy/+
A1wxJ5yDcUELGoX3uDWqLnPNlxxX1of0Lamo2M12UYIWt+EsGc1AQPAk0PCF0VqvEWpGhzWrkSOv
0319cZfh/EPL/POXXylkMzqQ/XlXyAixq+XfSVwz2OdZtFTXTFpFdO1SBi1g+ElqJYllBO5Bgi1C
1dX5PVIw9inMDsKNqc5Yysu8Ro4t0DZaa4M5sHx5W742yhc5Ug394Ue1TNFxWq7JeCUTnwLWDDa+
Sx+J5eJAQEKAGhg911QIBDFil80fvNkC+yuFkzvLRYOKbaBBkF10XSevwizTN+CijhLmyaHlzvWj
PB8A/pGrZvIcPBX0fJqOhVoZhN/llZbz/qdWc1E8sVH8bh7NNN+IjxcRBGLTTbA8MWfUyT8iVfaY
gIwdPsM1HzFjrAtTyH83V8yPeeQTWLjo6GnpqcmXlHPfNgOS8l8wDQvtNSK6OJhWUEObSMcNJse+
REk87lvz1Ku1rHoDeHGnbZ+wfk57DndJtOC+CuOtI1iQJQLm3zeZsTrClW/8RlsbqcIIbCgYNn18
UVbmjLlJwPdBdfMQF+ZQ4FBEpErZjWNVZ9ScrvBI2IFQJodpyzTtu6JzDa4y5l9kugBvrf6ifhFS
agCjMcQxo9z2/qaFxacEue8Rd28YvPAdDqF/shmOq0OwBu8+dmcNjsP8TMAVG7s+35pwPu1Ep5+b
9H4f5lvAn4MIhi1wqdUwOwqt8Xs/y66Cm/qGZdmrbKooeH/chnFrUbXn5NpkzGFZG5ZXK3XHzxRI
WiMglE/84EtKQMqOVF6VYcxcZkxatSj8SdIOUlr/D3AWO3lltsoHeHGk4scr//EtdBfURvq3qsSJ
TnBVOvwfZDbYkQe5Q1DnZR9+53vEhXyOxkKNTlzQS3Niiv1K6e+od1I6MSs5JE5Q7pu7QVkmeJuv
36VkohGiIgY/sq++Nx3mEDjKNAuBUA7S9vT0d7OymXEc6GIby3X/s4J+M/kXdAXf0O/a1FPxRkVF
ro3ZhqOD6Ija5w+1/XUuF4qW6vHPujhFYbtwiamUNIPgaMiH2FCn00IkxFUV7rUOd44Fs1HSQUG6
XAY7SpYYPr/6/tTK/yGtdl6AHyEWz3zDDNHcfC27SKZcUVyBBARoDpUso9Q8qFIWwxqh1CKZDNb+
E55pHhiEbPkM2itAXKvOV3RvLevoEw0LoaTKiF7JpCoR0CGT6t6w53Mck6XrPUQ4WdskGvj2KwiY
tFZk9tovA4Jj6+EZcgjdTNqKbr7McMQU5H39zzXxIrBPmujIfx+k0O+Mlzu44jrpFEq1cN1eaRf8
yte4+BKKgaubX3XY2pBTSRwoKgzLzL76XdwA6ZBbCQUCfYrT4oXl+arQM6e6HPN3IdGs9IUUkEKj
xVcgzT3ohxLkGivmD1fqd3emAS5Nls7VOiLw+I7La5S5UftzrKMIZxUxKFsJQb2qGdel93xOf2qt
dhxfqVdQmBsn67R9wUtj6357DlOvlpSfDk2h3Yl1DqKyzo1YivXiEJ/r+VenxfaZpwm0DlAWrE+k
8cvXqIXDjrZpj9F9p0wtkxWHKZ9bhsNHbASf4k2tY6QlwrnCqXl+3xcyEUKlVDLXPB8gVlbnrKWY
XVcM63VSDZHwn3kBMpyX3mVqExpXrMPvK7IAfiGI8xn9ukrCjrkXlmRQX87qod9Yth5V8PpwO72D
ZcQBXJoWOvsehne46SlnDN3P6mDV8dXigdRxq2xD3R3Jdb/B2fXMKMqVIpEkBofUTxkonqeGe5e1
pwKZ20bQQ5bzzlR0l6iMEC72LSa/Ar556mxp1GZWv6Ku7Aa4k1el2nIMw0HASfpstUCdhRhgTU2i
7i3Pj7N5xLBgcfc6sBSZms/ZIwNcrtEkaiJeZREWvx+LreQhsP77HpB+VBnOtFMbpeOSwSjLfv0y
VwESUOWQJ5Oj10zEamxWS6lUMXnyUZW4+l+y0qs5eMFJ5g9VtST2aF98sx1rcSyG1YtWPr9I5cSA
UhzcIhbwwEkiXtZ4BeF1CVz0oQe4+OeNOeukLIvJMxH7E3iCjCstGIIOPUqR/ul/wYELqVLVtuzK
kBRVqHuGWsBiv6baEdKisecoBCozwnClmZUu5D2xSYB+s9EV4w4klmqdqnk+HyCW8dewI/u37WVl
0Eq9E45CvKDCh+YT/EmDvD5fNtGD1WEZsEI592Pl6V0nqdM7fMilH7GWu5E9dSnFWv1qDhmu9igO
/Ul4dkl9ufPG1D2LHp1lBUL5KccpRIedxIicnLOfGLoSZASgzSTeTS5BZSNsBDRBgM+z5u37NXdL
iVTCuF9s3CKnOBEbjUdSJlAS+sIwKO/0lqoutuSh0oEoFIk/zVAZhjwtKMKvD7Rq6IGzPTkZFEkR
/13+P1oMYeAhJF2Q+3YXnalBiMxalURSNUjXuXY3XtulaocUcGwI1m6GWblSXkOPY1z3zYW4lN2+
FN6PXIGX8WqWgnq6+HrFHO/1YpCU99CSuIwinETO+qcgL5DnhsjSSg5667c2krvIPsFpeQcGtnOU
2exjTilLSILJhioGRtDqEdLRl47T2FJDkHWvaXN4/XgRpIE8sCkW3fPo4vMEiofzYItx2SrDU3vE
NS4g2ASCW+gJRAbEYKPpZqRoVBE1MRbLdw1N3qVxPz3+VkA2GQSwYLx4aqu3pFsfR80nryOi9voT
W/btbEKnv+mblUnZUSVGwIWmT9NULbUmYLmjCO/zWXD7hXwa5De5f0QIjDvtsOMhdI5fylfCHWGq
UgqMvNnlcgOTu2v/o/kMUGRUvvYaIDUBv0fgUTE3nXq3YdQhanZcFzsiqIuP7d3rwa+06G/qkaN0
o63fM0N9s3SY6YL+2bisRbPoYuHBxgaMXPyMd7sxmEXuqxdrAhDmlZXGhxdASQluMyjdRK1pQCDz
ZxRQIcdAmzjHc+AKpb5cv4xkwT4Pyjhn856s+R3d+/OEmPRLkSMkJhe9j8+U+thDb2YKcj+R1Hwq
Xl3Bh1mfTmgCYWvSd/csCkYKYrrXVMngsIJXFpl6OSdP2FBK3ndwtLEQfvH6QtaEkxFn6ukcYiWp
0cMxdGip1fqsUWZsL9QxcKDuRCkpWPyNQHlgHG5odgwYT5U/MatolVD/EMJuKCN0R1qsSOYCnZQx
u1gBlVTD+fUpaM5g7BcTk40ooqqBTcreUWiCf/5ua7sHJTXJDWa8IcdkNDIUvuMWbxBT0RXfGP7S
RHf70NlajbAi2xaxsA+ShBeRJWSxgscp4OjppqsKDq0thGQzwhA9uxoUttsij589BoQYmlGRpkwn
e5EqKJ1m/QbAsaiEOd4XGQ48IROP0aFOQI5UJ2Fog2BLMcRULTTYLeXyyi38bF9kxijQ4Zfyk0cU
h4Z6cIAKKCRQ0EwNc/rxp6SBc3VsFJSLvqWS1d4vXUlPO/XI4UVZER8ZqddEVE8xxFacyue43Uwb
uRHV8WvmPsfIHXu2pJrI9DDtgthRBdEKcGJc/9zQLnTxCx3bXAOHXbKFHdrZyjBOiMHTeRd10fTi
wP3eyf3A+STuwFgRtKLR0DUYA2cuGOjf3guewbqIOyxYsdIs42z99CeO9rOAW2LFD/AFNOl+6s+i
0O28NwiIJmgMshHB2wuimzDIaLcoNsQHbiuAGC44Vt+gdpcojXHcIWcRIWYpt0qdcPga03SYcv8z
h7/OWDuiqxVSGDK46gBDsKk0SnnymO2bWavJyMKUplYef5lwxz4zQzJ2dBJ2DUGVp7MDnLi5IzbJ
E3gDeLp3bf68PuZrQd2NwfREawrpAljhkqhywZ3R43j60mU3U+RiaHj06pQWEsQlXMLYgxPf8zBl
F+7qTawUrgrl/typpLn5LeQVeAXdXuGJCoo5zNTxATaDQl7IqSZTk/aAktZWtcyXKSj0280hD/jf
v/+kYLWsGIVQFbHKTb9878zEHTrD9AQRBpUnGPWenl+A+wnnoHTZIoH8VIq4c3tCv+smzuG0DgHC
IlkmQEhFvt8fSW/R5r2uXLnT6UCZ42B8O1lgdtY1TmrCgROCCGVaF927kYus5gz5skmrDbarO8dg
rjc0or0JHV5Z9+L9BYpQ3+CvjvVjKQEM2abWs2hb/yWCQScZsPFMJMZM02U3j4fTe1yD/tVz6P2g
yBSK85LeE7ekAugFIb+neUqxqc/xScD68q19VYat+wiEsOdT8KDEC+1L7nDRcDiOI567OTB7oEMS
2kxGt+h09ZdexgtVv4lr7ngEYXh6ACcshwOYhQBmcFMRkIUhycFyonY1RXEjIUSWGe9vk6IPNfTT
JWql4VdLzLJfCHqw3yJ6x4OdUmU1I0EtYWlZN/VTdyR3i91PyeLGcEJe07/nGP7u0xIDU8BhD8WP
Iso6WlyD5Uc2UQkPS4Mt+TDqFhsjZLsuu3MJ6S3TfZ0QkrEkeeSrZOLcDqZCRXUnSeLmcrHwlyQB
T8WNcTpXYbG7S97LHNXxBnkl/uQYuF+9Qy1lttODS77rFFhwDIPZbZexth6CGvRHH9Ih29ufvQMR
k8Xs6t2rY5XZ7ysUoE2hgFLfsf1BqIZHy+tQsyCZ8wc8YHSuChO0PtWAmjbMOXqPYvW8BD/OtHko
uVKSqeQpY8FO+dOh7ucjKbRB+rWPDCpmlJNqB9V9CmUD6dsVv4an2s+CUwI3wR3xfWdz5UNIZbFY
5bj5r7fl6GccZg7dih4oi33ug5d1bQnrL4HtB2Mt28WJvNxaUUC+zH5JGKxSaU1ZD4aFDg6sn6P3
eUiLJWvGpz2OWR9V38jiDY4avFyF0I7+Ef6OBqebaVTESSwPdoHEBN6mEXbb+OgFK2Z4ps19oUiV
vVWKSeKeMqDsMtRghVi/ScYNphwwjBIAlQl7FUt03C5QsLTgntUfqi2sFbc+vTMQ/Ijc/CjMCMWc
znXVD0LoWFgHszzhwhJpKxpDi5nFYWPajLpi7kzZorbdibB3dasU6g9gwiA9G7e8cVmgdXMGOx1v
F721ADj2ifUUwGj6q/+wT0pvYKCqYM7cQA/F8REbHAT8+1GFw8EukKtVTHGTSJF+YG5CuzLWC3SV
7sEV0jdKZMwjv+5U1PMW/nuwIrR2k1DLsFb+oZ/GOFXyV2yge2mz/oy7ezbXJMvYaEMvluwRY8rI
ABkip5xgzxXgpbMT2Ga99HSuO127+oMbb1MJIBljJpo5+5GYPqfRIIJjS8FBCX92e7MfOYvsx26f
EPTYixVbgC0ytd41giCGMTsGaUQ1+L8tYVnfnbyiUhj8lufV4BkA8b54QRC2Ms42m+wvwj0gseij
loCY/tWpZ9lOMtBnKcouFEU64m2CgLPhL2u+cyms7tVbkchckkunTDChE+y4/A9cxLOt/G1MUQPT
CvGbOV8ilbu4B3YA67/QsWOfCFa+yBj+AuIjoGUY8DRIMLZIDL7jTNG7WXsLHuM8SiYCNWogqhaj
LsTUTmlfusbOTh5Ce6BbCqg4nXWmUYR1Pj9mbDI/Yzo9EiEc13nODwhaNF+B4KyHfD0M2Zq0gnaw
p71bhFZBfJZ3Vif7jLcaGeOqNgorriGiAejpm/mUZG3P4pPkp4tYA5Z6egqh80PPVv6PSZhO87WY
wFGfObFj971YFxQmKm56xaoOY/GqsxWtVWZfX4QBxEGerZxgPE2LxC8jwmwI4upfw41Gt+uP88AK
fR+gFBmpSvqxacyc5nk21/wCiwE84iFDOj+OfkXmBSK0S5743S46ja8+jOmUWaYT9/GCCjm9yw7l
aHM+hHYfx4XWJRw3hzPlrW/QzTXt5EYV3nNya+k3qG0ig3YUXt7RheSWlBLlXv3/IpFErt3A4OV7
p4TYMUVxVZwSg3z7So7mWPzRmzx1OpBELqX/hHGsiBeBCqklwTlISNXHoSq+IvC/TXMUeih419A6
NHkq59jkv7dCT40yNQXuiORnn3wx8o4flwAYGUpx2UWF465xjy6xyP9pdrtkZCpvZdS5fWYrrtqZ
FWkBtG6yFK7rBkTwys5Ju3WcKfTI5Cw1frYbWEOYpq16SZi15Ge/hogZiXKhe0/+RZr9SJYdoRf9
McfEwSq//NMzB4F2+qA/o0NgRWC3Y7mnYiElnAROJh2j+1G1gEADtoAXRkDti0SP/PfkE+Yz7PwC
z9EmepcouTdWP/l5Bxu0umrdRR73MmQNVHuS8xxE2X/y2M00Ru1xFwEdbp+vUVfqbXMW7cEG5fC1
I3jYJT+fproF6bt0wG82UdRpr0O6TSRtSoEoREFQAp2/U5HVSCSlahN5uPbHcL2YRTocL13wrghS
Fz7xx70FNWizH6xEqs/oTfCJramx01VSrTQ/ZHWzN8HZbWWEqpaV5f1SCXZfe05+2QcVsWOztkbo
JeAK+O9/VqdXHmDCLGF2hj2p5pKgaq3fIVr5eL9BxE7ntOnekconFX737nMDFsbNLQZiK9lSD/Q3
W2Amd0F5z0GXnsmRs9zOaDCvTM8NJQaLqlWZz2gkxO3PgLqJL3GTLhLROoRvslcp/DmquagAnGJJ
7K8oybvLa6jcVMMAJx6gH4r92DFTuTejn+yGm9msSkd84yMwzaZUyzDdAJ6IW+JDgM0Zx7eNzwNo
dIPDIlgWqyFdjwnDJ/ZheaunJY7k7VcXX2hlgLzpBnurmAbdPJaxx8bb70N6WJ1YTfbcvCFRxYgV
9GYUxA7+gjrY+YVfwbHvzfJd1yXht1fLJ9wdvIMKgzAjw5pVGvVWIm61DtguISf4C/63s3VXfgiB
LBGkXXAndlmLYAmVskGWAS7wVag6vDaREYCw0KyOmk8DmbV/JsFj6qkl+XcmtLcIN/W3UOIzIxcd
Ybve7Tb6jUlb3RFpyEXds/I2m+3OOGl2ZzvEFlZk637lZJlm6tzjUiYAaApoJqnfKJpf4L/TdAuA
DoPlnDG7FZO6rFoov9CywKKpSrv8wPYPMEkpTV6cSlC+5kDmGnXFUbQPAKmrJDrQbyVcaKa+Ys8h
6zWBWw8Br8wOiBjPzlgWLKaI0fFnJAEwvVv13KLMf3XG70lXBjobEdEjZxhN8l9LxSCYSeKMBNlo
sgWB+ro0sxgY1V9lwS9tjqoA/+xyrd5LSBJ+kME7A9sva94mcGae/VxfLzqeqG62xBy3MdlmKEjr
ojv13ukCXK0nkCHXyq4f5pjazfTlGOrWRHwXsVm6K9N1KaUXJF1MTeFArETwCleGlnFczBaWovQo
N0swpwpm1qqXAnQPi4KBcDk0EGEatxOvfeCYcUisqmfDgXJkD185CkXJi0Cjum6viCccNxsSrTOi
SXwMvMHWYx3tlRU8LXbLCtcydn8X09nZw2N51dqwACRN0sHkHT5g3fJpnc7zkPhcScM4ecIRhSrL
zcLUhKk0+pZ2G55AYu3ELwwTb6mKXfHBJF9ElnaLjIqvX2Px56t/eYK5X4t1encn78sTnylU/kM/
DqJUC0btkxT/LdWSXoW4RYDuBrLuDSKbEDfLp4pkaSkBonYpQIE15Wq7z0IUI4Lxitqf/5a0NQp3
9dg8/RKudlKCbR0sACtBsUAPcST+Xy/IoRPXALnZTf6hFpt7/Y+jNdUyD5MRLZ+IAqmsSsg62VSt
xgExtuEpJUeRiQ2ut8xI2vmJcNhSJtfqj7TZEqkXEX2GziLOQcw8Gm9OD4+SDwVqO5S/MWMjZjLW
AI+BpTsVd+INYyO2i+5XOBQ13jYuqyKCVdMjUIG5iN4t+2tjcoyUFs/oxnf7P8i5bE2ziEHoIc94
uXcOgKzE210XsQZNLY5xXJJWuwec8wYxCFK9z5Ob9x/ssAScUbdCureR5EIpoPSZxLcrhYX29k4E
yxfP6htIQ/Oq1frL9vu7eahozwMaN2ty09f5KSrIOKRiDdurhPjWUvhqDN0DRv55ck5PUddyVN+W
tUB7lqJX9RR89XH3xlLB4sNohztsn4B80TsU4nXeAYHSoqQ1LGz02l6ESbICnfoTbuwiMVT46dWC
OXkmrZ4TJEinu6Zo+I8lYLVWWox6LML0WsrSWZ6qdiwzE+QTwcJ/21xgN9j02X04F/qix1dA9l+7
RLhyAvuvRdwnnfmN/uxmI1SRKhp0IeSNWwxv80g/P5HfzPAyp/erFWH/5kWRccSpP0N3hwjppaA7
5DriOtC5tqIyaodGHE5Hv3JDtfQQ4jOS20ZEXboXCuE5ALds6dipL7SaMN5G49/3NstLOWK41ONb
5oBNSW33wbMlOJnJBNDr6Y8fvaFrW1KJPYLXNhgeuTwPcXGbndYUZWLOei0fVO+ECRXflf+pBDs4
VJIAORW3ew6XicBKbW/hDhi0JbAkS7MtNsExySFDA9rILsq9qfNQXBHj+vNf41R1OM2NDweWbf9k
3GDAArf73QlorDaUc4LyVWaO75rS3cznAC0Mm7RdMBRflvFo6kQwMntFN1LivcLkjrkfFhdHGNWY
l1micQm9tbmvagH78RPNg78OgVRfCRBdaLk0GBCErvloZSfgGntSpHAdM6n1CoRJX7x4wdLL2Ofr
aiWU38tjf0r/blXIeI/liBwlsuOKnBMxccuZmT4j9t79JkHOUqRilMQ6ma4WaRuLNExdeeFbpVSF
N1Av1fRls9pwehYu9xIslsqlRfXHKNPb8Ub2ywdPufzA8ttEnbgLkk+EAgKTLOydd8MXd/ADJb/q
4VqQMBlNwP5dhTSo/7YgKvuJRCqBmd3nvAbNSgP/eVhN4Q3rXoAqEonuw9+4h2+BV9y7T9PQqzG1
0ADBjvyqhUNJtNnkUxdplrcO2EsE3evjA23Db6w2Ez2IHfPyoaKFnJRQj3BH9+tJpfmnPZKE60Sq
h+j0xYsgnnJBZiqiQNyKzNm24NUncbHMHMryO+LObtVTwCZ9FcGKiXxU3o02KyVx8NtDVl2nYlPp
ouyvBIgK2P47jEwIha5WhXDrDgZHEn8DmoZTDrdpZhvDuKWCMIhmlWMx2ZSeTGQB8xwV839Jr9Lp
LDkG6xiubqv72AjBYoAKw159oUoCii9GUkgoT487OLpT4WkgEr2zj10lficef8WGT+UlCHPgCmlF
Y7RcXyDR6nj239nho6pfRDPpaJ+uQ+ELx42P2rCgTfNIYHRxbrDf1ylAUtSAiRUwc5QCu45nT2Nw
OAvqt0qGjB9irLPjSFEruZ2F0s0FokGxQPlBVZQcWv2qvILqYV6q1ppLCW8lOITswfRwPB1bbONm
uyiUMLB+tbszxJQV68KFP8MVs3awM/DMvmmzDj7wFR93L9dSmEftlB5RACsadTMmcpYAO1bKCaFq
bSQVvR0wKH2K5GjrJ8SvWfqpzI21peibh7k87ajHFa/CBNsy/mI6VDNfNgHL4lB/yBmyj2GwVNAX
iAPWU10coImbtKzB8XaCVJcKpswivKnMmGy1gW15d85hPlhj9T7bk3fTBWkbx13l7cbD4eosau02
llZ7H5UJ1+YVDSVDpEvvoNMJOEzQeizgWrXUkv1jgIM2xZTEyw6doKcHVxdGWa4H9DVTDK3Ka973
DK0HTDO9aWZqPg8JpVDsGA3O/5GSCUWZnAxrE6kIAwaVy82C3leujmMEbi+nFUpO7KiHRSf3VqsG
KBsvwh9RZorjo8ltpA/WMb6lqPFvvcq9E8ZK2Qvtsi62t1gvs8t+gTk/P8xWEN3Es725V2sukS06
pZB54EiqbxDIQV4srRLSkD2wEFdET50EgzICeOaL+ZuNfJukZ2SgJVe434YmjPz3LXHsJrK9NE42
bc7HuROILw60Pbjg/S0g2bW/iswKyw848I0gfgD3JSARCeZGuekf3QVIHeC1lZ8NSupNtJDVl3ST
TlzKNTC1B9D/IsjmBQX1ySQxXGz6yA5TLb7ehgVm9yx+x4GSLeJwA36rJpKv0MdkWsFxvU3Ljn6z
Ya0oTLWBCJoL4/QFY2x4UPMjm6Ykj8Kj4QTioNkY8cvSvcx+srpAGGK5zp79oIJri2AQaKA5fCif
QlHGXbH9uyvtVcWcjv6DLeKXe2Y82e+DQZSqlj8SAu6tj/ATFHC3PkPaPSoVsUAtno7dr6Gdis4+
kjD9K9orQUaPYjFRP/oJ+nWR0ytQcpuCd+7BBwI6McUWdAoppVTuzO/U+TkaVRWVxV/qVnLD08NH
WkSZfaND8XjhzFCjyjk85Dv2sDe0qjor51cfaeQ4RfoPLHgp15SrHPeHxL0f5MoBuJvDlFzBThkg
X7toBvuYUras/mIyOcvHN4f17/NHomYdxSkhNGjPK+1qK1Us5t3HNk+Yv+BC5mBus5Dz9Q9t4suC
uzsahcPLtogXwSao7aatcAXAsIyJ/5er6dsKSKOJjiBHss2GvNS0KFXQXb11z2Tt2H1bTR2a9sQk
UZ4oAxS4CnnkbrnoPbgTKI8sGfGOw9YKQOXLDLOcyJWoEYzobC9tGPGNMWB0cUynZpiikIkur3nb
EVUxYmMlqKy0SKqNV2ER5pab2ueS6hROPNdZXlpSXAVWK8z6CnvS6+v0iHZoh803q/yHY7q0+ct/
uVvTo8qKu06agd96P4W/qwZvN5Pnd8P2bg6eoA5WJraTWFZg4CCaXhDuNuH4nopbV42t3BoP6+tE
MEaAJ5Ke9ZksMecNJ7MM+Ah509D/IOKNejSAVnYvwr4AgAK2qMi4moP5witXzSEOX9C/pWJkZx7u
7Zal9WUIP7fz4hGb+/WXdgyCVtkdIbaZIqNpxtKH9SzH52L52wC6lyFThueT5TgmwFGcZ382/Ix+
FBImw/budIxCU2iOhw2qyuVFzuj6C9qahR0aSdLD6lXFy0kz9hcwewgGW/fswAvdlP7pr6bCTw5s
bm8E9JEJsly/wawixxkcaAziXHHBt4qk260hSvZ9IFMpd5IHpkefhQGQt4ajc3PEKyqicXq9gOMK
iG5xVq+s5UbrB1AyayKUzp/L7z4AnA68qfAp1LFPqj3v/UQ7OVgB+nv2bk8EsuGLhma82Z1B+hkX
G1do2oWpTmAwzFSeVxMHKO/vn0mnpopcqXRUbFjZB/m1hmi4BL9VCEkHYCCqeUzc5dnGaYlr2VOb
WmLGsWF8btuoGDpk/q4IKGsp84NvprtfP+TQKqpAMnS+pySzuAatnKD/x1/DYRSXTTM2nJhdiacV
4Q/naJAqptL+u59TS2iTGoBNxEQnJSlv3mgWl5DVJCEgJ+xzErUCjjSMiLw/zvq4UtmK2q+GS0oj
olCyalVLAnznqxz9sH0NDN4jwH11t7zaTTn9D+L+6s6J21D+k3tJhRW4DUIcU/T03VHkCfT9AW2x
Hk24Tfx/tU4U2syen2QAC/qFPMx5x2jpuhlMJn9mM0EaAQg1xuCfNz1fSXWGZjmIME2jjWUgJ0DH
PBIjyT6csbDIssSCAfpWWIenQb9NS/9q1anowr8fl1crQMLAeMVa82rmDxhhruHppOOE5QkLXjaV
2mCE1d8g8tNnC9eFkqUo7+u3uNC3EITLpLXD698eumxX3xaLc9sC/GbypknTqqeTh/VWTB/7jnMe
X0LNUZXD9p8ZHQX83yIG8Z5LmE0mCbbbQXnk1KEUQlVA+wLY7oUlVnnDG/ipYaXa3aH6v+XA69Rc
1Nf3mRUVXyFd068Ze4M0LnWLzMY1/K/rzFFb3dkMqIcDC1ANkkLRPkhrkmphJFO28uvYqYtjtJmn
VvhX9Wz8JZZgN9SuX4QkqQHLiEOpn0VSX+v5BR6XuGMs4HpOIzutxmntsmnriTFY7X553CfJEsiI
ak6b1JiaIxlVMdPFEUKKH4ebom7xtgpJGDqyAWqJo+zM6aW1ObFHMFXdzWCOQrZW/VVikeMTOGLS
+YXWRhL/GqS1Q/TNI/uOWX753Fwzc/5L9JelvvAX5dxUNIT5CW2EQl9KBAsdDNlNDYAPnVw95Exm
WbfeTzhTmOEWSxEti2rQu6ljeM6NXRE+nBO5bNQphdU2+sYVp9MAGKVxszgG0CXcC3rB92wRMMQC
rXF3Gfx21z8TE0gJde2ZJ2JxKo5Jpb3CXaytCjmqI4N+paSB7ZE6bGSH3nJC91+7YbAzKW70dHiR
bgSPYcWdiNyIdZEDWB2XarcwYtaxNVekNB0PesJ2s0PYlADFEfKTXFHQTqnUdGFVBhNQoA5KgsHY
/aOsTGXVEDK1MfqBPK4Lkkhgmlez07fBFkVjnYOCqCp9qYv/WAejddPEx0p3x79++7VZLeLZ5P8N
LzeYigCF4tyWDF1mhWanRT5xkAVO4k37acQanDDAp3xj9cFG5vMZa4lCKYtnynuep5lp7l1zTfHT
J1/AWtuddxADay20q9MQHLBoTGE4okHZaZEi18GUiHXGJ34S3vve8hrwXVR43ZvZmrM2t0LJg7rr
HGZF4Utv1pbZx0jUFKtIEbIJf7ejNp7TbEZ6Kd8NgI+Dj8s15vIXi+5nqVrNL2i6FT6ZoTrYn+6I
QpDSYWMLi/XQU6XVcsX//BNpnsN9Ta/+CEchrrjWvaOg3G//6PBZONGjDN3kfE/nLEzSrqWCCXo9
Vi8UJY9BZJCTzIzfuyVQmXxuNzbExllvmTwiTmp6yhu42sX8KPAjOsX2sBP+KG9NAALcXBqTAH2r
y6yg+fGjsWxiGEsJdnPEeiwlTmxTKzSOy/gOSvf0hYNK6Bahr0nCC3opwDQK6jOjQvgsyWnWHfiO
nr99cl1Rju3oWmmfcFu5Qm6X+NS0ZyfdERHFVSBkziqyHMlirSnzI5pgc60DtxdSDKIvOmP+3xzV
ycZ6uOGigTSlbQMWvGzsjQ4+H1lFG/zwbapLELEQnHjXXYDz0zRTXYZLxys36Ki+mdWOLi2LaKra
t3Rqtsi/NXlgBaEW+qM0FcDlC0F79SvtRn9stWws+bburjb3qvuKA1VGV8ifYyLPYBs8MTJ1rNsz
LbJqcvuSaUl4Tl+wAq2+seEwVWBVoNyufOpRctPEIHA3C8QNNDS+PGbw74+QYNZ3ssc1bdlwQBO3
6Y8pxu47M2VjbTMG+TAdAuD6xHY8H5Je5Xqy6XQ/e5VKM4TUV2tj9gxVaKbG5VA1TrRxq2b6Zabe
ibE/0B/Tu+T9j0uYDgG3RdVqmCb7Ir6N8U8iKuuw44ATAEnnSajp0+RmcPRssOV082u7AF2lrfz3
pyEu2H2ivascz06mqfgTPQ/wmUjdV5Y4GRLDxkIhD9/r1DzmROdrl8CtZ8pnc7tmqKcArJUAxaBe
hjwbkTyzylPmWoOHlHSmdIiXu0qomPB++s+kYUh/oiQPR5sYibLnYKgKgIXnC+4/ROI2+xNRS/3B
M1bDTsxUJFbwbHypcnp8JNLDXzFWzn8iCHyDd1AuaDSIqOdiy4aLjglIVtb8BZM1w/+Yl87d6flG
jGR8N38vxfnYp0OdGmlwJz4Y9GNNZYTsAwkLHkWmT13KwD75QXYZth6571u1xs6Kpvs0vDyuWNCZ
AKcmolSL6eueYXCjl3frMrx9O8YQvi/zbx+UwAkFxL6qSsmBBOJWNcZJZ/rWQ1cRH2nGf5Ic/c7a
0zw9qthtFJM+K4h5/BGVOwtFTtCgEwxrq4WVEFKIilPwgOpBuIaDix1nbopwyLr6WjU3WyNxHQ3i
SqJ698Sj8OKgmjLpaVWYf17oZbWocYgeAW7FT0z6xAgf3KXU6TkvZI9/Pmtb2p+f17vHJYdRzB+G
VZag9wyJDbU0It/tIr3nuHOIiZvLRx2dE46Mx8c8NQNrYPJCbzwlWf2XKso7UH0w5XmlhagWvOPW
kgfU6mCYf5mz/vgH6wm7ELwWlPcNCzuFrCbVb9v98KY+lpPvzQrKtERiip+5MRAvcbkv/5mouAT7
6b/2vPH7aKHdH8dLD1hZ3YxMYUwECUh9XbO6ZixQBKVB/TyzG4LBzkXi5zYxGqvyx3bHIlKlLJKp
bDOk90q/L1D46d4SI7kAQsqKkvOALG2923mFKSvNSNBjsY0Dlh79Hx0Br5NqV61ZDWQTC7+zr0/Y
rlyLqbiFIYlTH7ntIQKX31yeBJVxf6EbUIIhYzSd5P+RtO/93g14AkztgzVv4smI8clwGXQ+CvMY
7NsYxA0MLNbpuy3R3npqnCogzweeqcuB8U4zuR5WnNS43oUhkX2S7w4MKVJBTs0KkGLTKAqNbKaP
ssfB78sCmgSM3avlBCiFxHGAKmWz2u+inUxzeioqf+JlomIFVA/wOESgSQHpO28SkaozfDyxoGw9
UKyK+UrI3E1Xjx8RFHBhAsLChfiC784D/AwzoI3Jw1Oazgeuitxwdqw7fGGdpG12h034Ac2zkU0R
ZIciAD2CZna8VzN/WdG9+xW3YdfNANhYYnToKZLGWe+OjWsikmYUOQnjUzQGBPH6XB6P5mefkBj9
teQzSX8ivMNOfX35eQ0B/iVcfHq4WHPITPOJ9HTx8g5iqrBsw4jm5jTzex5Wu436Np2vXEll23KZ
BRtrUJPKYyQ/+9zIJ7PDSgudVZ0QEWsxzksoNY1TbfVBPTxHlNAFbJx/HBA7CvY2j4TevgIZal/R
btWX8FGgUTMmJ+2KkOk53k7fqWaclFkzeC9d1Vrt5si4fZBNNfNorcR88FL9FsjcCeFfXesKCom/
p3EBz+DGLcXMdqMz8jaWwAXeZSxh+XVJdFTxOzkXkg/priU2LmQYuZw/hj4OtqTyBGZHz7yIJ7SL
4JTh21e3rc0onZ0w7Fru+zFd94+iqyY5mkF2MUhwchxZ6A2IaaS+YH4ozsro/lhxsG9eJB7IF4U7
udojey5EGWnybLdFmGiJAdhXJytEgZaJ+GTXmj3nJz3e182MyMDXeVUIzoANhJZunmKaw3ImvPSU
cP55esttvwjlSzmIeJ4mqdIi2utPyXw3AHrRe3LMRGQ24UijwoQmf4T2SEZP0KXNnggxkBxXap93
P/TYZYMcNox8wQsqQFHgfGaH0ItdgawEeDjlaMVn32RmdQCUabFT6WvXvGHVOKc1eM7+p0ZWWS4O
XSYfwGQR72h5Y1KBHP6SzUDnMfJaSvfHNsLSlgRf803cvmWdSLeVpSPfzZaDvkXwveXp/stX/eUt
h9pkwTHZgM7cVtuU2xHNT29FPDjnC66ztX331Is0FxZ4NRnRBWI6dYwQa2Zn9Ur9YfGQ7VCOBCVu
YzgzOGDgK1/TMa0gDXpAEyKhzVu9Z1FUAulttddE0Ba2l5ZWcWaA1JoJyUNTJAhq9sHbdpIn8NmG
qe16jlBcL2HFLSodGmsnH+P7V5wb5crwAulIEcTAd/eYapBYwwSCNadUCQ1BA+W9P3zXA05BDXWr
c4MLa1KrCapj4+DW6RfMy2LTazY42bKrjEWEjZte6JZKephx5ay/2n3UiNCAHlNaYLW2nrNznkfL
D2GLKMvsZg++t+BSg24QJzF8sI0H6OJ2L29/ZWqME2SYr3uDPQ2ZbllfpQ6s2c6pgPh4sDzQwz21
jrHbE9uVfK1su/R6seXkMWVCpQhcWZ7yIqzEeo9JA4W3SULkz3dUdyfP43YG/HyrilnYgag6Ct4C
W1Rk5oO8/8IXhLGSjsMqj3KThgFGwvphFhW4gvn4EX/tw4YWDcS5GDcPoKe1ev77Gtrdi37IItpJ
L+Q0XYiJfMIeA7XhBvKuusm7NbI0GR4TKLdXVH3VhFlqKtviPq38eaF0zZouh828CttJMvhXf7GO
kgxs+MvC0Nh8dKk58gfh8ak8Eaz4OWzxJ/f4iI+mfzZL8JleWfez6cbKBsMjwRh22ikaAyiUDWYg
rPw+GlUd8lNIJIKB+cOuIgV+zmk+El5VM61zQby03TjpGvgxWPiA3qd5KdMpc8a3ZhZ8MiHDcl1j
oHWNdMVTwW+52BvDtfGV2eB+fh903QsABu3JrSGqbLFeDT4qwE+3INDiF9s9dnMP+Ke4/JmRsdvP
SuNuGIJZDv5k+3NrjoMZ1knvXzwcSpDcY9P1qZr+fSssw3NLvCHaERTiM59/FMi4pJtQ4dwr7qYO
VwaxUpMZcvTCifGm/cbT9s91MyWzARee37ZQc0nxJUonBfZbbtWx1zPSWbHCFnK0tGmct1oE7lj3
6e7fjV8KbZQZMJk8DO88AlIBmAjH925TbeNcztqI2+0rmLhe/BH9QJCe2oOjJjEpCUSE1IywwlnI
MhOVbAXaBMHo0C+dLCUusJXZwT1jX7WMyKtLNnDn4NSOeVeJ8GU3ulgZOMgBzKW9o3KlGTenvKPb
KXZrcqOwnTxRbV4VUT8VJGL7Ac3snCei4YexzzL5iOsLmBLZBi2/DX52aeH0OfQaIV1VGcG4sb5T
4RkE2kuKuKxkQFFLLjzwy4+d7BVR1Le/LgocEhOSC4ZBV5yebLgZc8TBWqiuzg50sRxqu/D1e17g
neakHL2cgWhU2zXhbHrFNuT80A9JZe9ia5RI0V3NMQ1BixmX1cRs+4sjMd6DF+mJpp1IoIQ8mJ7y
RWEOM1H4Ga4qFpbG5YRAFe8lGleCa1aeQuStc5RlzPnzV86cP0v4PgpestvYnCJ9hqh333spWBpq
sf3QBlMxcbUr3IicnKmV5uiiRb323NtFJ455x32WBy71hoi7iMwIOjpbnYBwVQ8IBpBv5ezNPX51
CQERZxkQEZx6Liw8AftUci4Hn1TrbmM0EO4OcWckObothgsXAUWUG2LT+Mb/738QJNHEnMLHGT2K
QkQHMgk/WRLcn61i9l1zzu0O0ZQhZBMfIyw0kYIc3QulX0rn2C4CkQHoM366FFkoGKWGKvb2icUV
TwRLCxwcH3ey76rGaXTWYeZa9hoaDA4bmB7A4njzoou2trFaDfhWdLIjUMO9nIdrzJCMp1ECYHOr
1Je75J2UIg6O2Fa/gRJfX2/+SJp6R+lUyCqymv7mDhB7BEdHsDwdRedsWkrJPncX0LbvXvk+Kdix
hkJ0xyvyToxr9pxRJK2JV2FsL8GOZTFYXuFqz7WbRfUgL+Y17CSveXn6dMyrwtSnp3Pm87YN/+Fz
p1WroaXwaTLzBU6X9y5Qo3sY/r+EVpHU1BzXu6M/AuFL79Ed/qvOjsW+EeNH+3LDyo3CMOJWYBZz
P0LhEHMSc2zKEyEkGUBye/UGXhqOgVMmtQgSe6/bC7tVjKmlr9OMlYRJf5nAuw1zizaCPBArDZDR
hsOxw1SqAjwJd8jjmYOUUC/Zh73lCFCLeUlAsyjQzrjpxOIJKfm8sGKZI8IqBOjIaOwm60bUycOi
YMqq5t3D54Y+23fK1vMA0Q5QbMHh/bb6aYTzCjgqVYoFnabWGVhWs/RzCwMJ0bqZQw5z7YQ9bzvP
yrdXkSDH0AiumRB7zvL8WWc+dRTCeB012AZ4W8e+aNFC/q7VebAF3l7W8S+PIIFulOkcNRm3lR6o
mk4EAzszUsKOFTmuSBw31Fa4rIru+swqslwraAuCSa5J02UYDGkjG09zVbE6i/LEJM52t1DsiiTs
ZIJP7QaLNVqhMLacVgDP6YHeREH6EbajSYkjkgbL/lQlskrGZnmDxqp3sXWpBIKYFqOhyDL6kLB1
PLLu1SG0aatDXI/1yq6/oTZVp7dmxYT850bo0piLuonGiThtPMeYoowYSi7UZ93SHmm/Rof3SSwS
sp7PJNfQ5oouvhcRNsM25kfBVjLc1d832OMELTsLCpGVtc06VwujY52hFt9KFIOOJjPKaVtTun4m
zk83ulav6imsljGQPIJu0jrHXYbzvZ/VkoHiBunB2rQ9qj4MdmKZxDPumBT1erJp3GEtbZoQGcKJ
w0GVRJf2WEQL4IfjHJHA7SI/YQ4q4nN3k0fQv6cTshqN5JquZyYcr5Yun2JvvFN9BuvpWnvABOHP
1zbtGzBk9+JMag587ESecf6ttogvCHp3GDhZpKQxRzxuqmWbM5gJdBnHXSq4xBuqzIop1X2OHlK2
Heuk3iow8lTEQf2mVWBj4QfUPgd36F3z6qURKJbzfUOaBxeZoC9AnDrLh021dAIQLRVo4aEGXxHc
198dgmwidMfZe9EWdWfkplE80w8GsznQcY58EyL/s389sr6OR48yh7uapvuetGzUn5M4s4LLVsGo
O0VbNISnf6n6+xlYh+Y23SsYdEWqVfHRjrhV92jgQIAsU7sxx/BOBOy3GiuVAK1eIRGvJjqkmYVx
s/Xez2sOdEP7yFOEA2xqDTMYjOqNvn1MUJJiUeju2kdsrqZSvEzEvSeHmR1Wsm3k2J4YNWZJ/vTo
M9QJFBzYA/ZDSeuBbCdHC1CwIF7J2a8KAXLGz1uvJ3TZWf7Lx9zAX0uCdw2i2sYBtPoWiAG/Rv1D
QR8JYQwpyE5AYkLecw/URBY+Xo+pHN1kdw9a9SZDQMHZZ/n901fdrXODWrWh2+zIRAYUY0gYXRZe
TRXjh31Z4rqdDCfOei5+lrfV3x63z2pjdxosvQFCYqKkbCQ2fxdtRjXZvWiCakkVfTyIg/h0P5Nx
C1wFm62ZAupoEtmVliXihiSUzcnREyG1YiBBCYcaJ3fucBK4ojJ92cqXGE5jvfBpMfe0NkXRUME1
VJROgjuoLLv/w4+bIWBtjMLJpEYOgSlUtZTwz/JTf+gUM8lzQ2e+NgAeTHzLwKdMNhPKb+71SCiR
6prisixQogsKR0T7NSWyRTo+Nm4d7OzRwmvbBFNAJ3AXMdlSKg70pRSzE5R8H8MD561Jl0FdwKdi
WarGZlHboDlnHgHz32g1uikgHw8m1dscAcODNIPdSW7htvgPLFkFkdJvZ8xtORyYquysC382Tf41
OVmKe4VQR+Ozpai+ALHLrmduLHYTr02ZBTR+FAmI3NL94UHoh3BCABu8tWBO9gwxWCY1uNTBUA56
7esg3rJ6dl9RaoyVI57hDtoGJgmpf4KN8XeYrk9UTousNjxiS6MjReWR3p9kodAwiDHfDlnpOgc2
nr/O5gQyMResyHmhnQkLl3M/fYFVpW9ZgcxBc+DG3S/SVTpLg3aWwxwN1+Kr4OjMXrA0n8OZUext
rjJDyahHTCR6f6vXx1WOpt50Wdle5KlsdhMzav4RKiq9Ri/XBx/J+OWyfJlNKBIuz2F5I1wxUqhi
9dOkK+A25m+aeOFK24t95Ix+xTnqKI+rs9S1xWWe2BUZBrBIKf8drngbIHuddj4ldCV9mHumwL//
aqHHtChk4R+MbJYlfhpP7aqgh8hMILcLR6FQnlYJeT/5bP/KPk/RbwWH0QBVOxwndPLlEBvHBJYF
DQLGtYxrhgCHeSsJh6A6G8bw4m4AUE4EyHetkgLvRA/Bl7MfFpU0p8HeHJ/ueJ/y71An3jpDDwUf
U8Hwgz0X3w7yLA8jHRPVUraHUdDBmzlfcE6HjdmWQJ5ypwRQ0PveyWACeRT/AtKVxu+Ifqmc9k7n
XjP8v847Bjje4b59f1q9j6meGpyIt4o/uDyK2IzmLocPkHev9OYg1CvhGKjglcr6/W0EupsjarRK
2n34QzmiymVZzN5wHeVUGqB/FAM1cNj/qnEx7OKpNdQhqk8pF02QsERMq2pCqg27Hj9WrfZuUz2i
Nc28MlNFVUPXEvRVCJLo0svzGbTQR+jo6IucDmuCJIG/xKFlerqn38+ADjRMMHHus+dozB/NifeF
z01d3woYKM95vH4JI2UlwogJKj4OM5IjEReRBcodiupyu859fzyudGqM2pGSEkhVLfCMCOq+nh+8
LgXPs2WVytfkVp3sMJLVcGs4YISwYOYaA2FemhGHSz+iP28KT6nFUo2ji02H0sC/POQSarn1FuDi
Cv13qgxKA9AHnTtPxigw/CIsqn77G/QlcHLGBGHPVNNu/eTHY3peG9klG826AND8TaZdBZsyaf6P
tm+Wbq8dQBBvWZntVBq/igzUqKMTrSqYPFLkEL7HlMKVum1uNUwqOyCKF72VI1ObfUA4V/nf05Vk
oSNzKR3Dqb0yO0LMguvkRIC8gTdHjA4T5lq7Bg72JWKe9vah2KgqySaoBk9t4KmHbkyJzXWaYa2h
h/3OHVhNIX+74ML7pVIa4wWiKcf77O9rnsQaqQALJnfV+Jjo4pfOtIiLJxMMWUZZ+b97Edb86oE7
RywNZpKl1hRTsV2YlXXxK3G9Lx0dTBsc+FLWPnARf8wVVKXb9Ne2urIMy6A4onEzMc8DOQVkIGeS
NFGhQZViS9c09UyYIgNrp+3esASQHNmLY9Dy5hSqb/jgqH0nWq2Y7/qx5lz2j2F/BRScr72t26Kv
Prgng5UO8pS/mIuyExrucWu07Jri7waqA6lbsnKi7vstxh6WjVf7wqvj/44QXeN6JDhxLObxPKNX
GMOXQDA6IbV3enYikprq0BW6s9hhSBlUQV7aip1xWlPKqmuC9iyt82pKhy74MiLEdOcnGlNOGp6l
vsd6XV7s2Gwm7/CdB6NFFf0bvu82Bj/9ntMpBVJlVHBqgi2D6A85Lx1KP8gB0obvZc1KXcjaEter
FhOIRvOfsVPGY7CfSeCidbUYSkQKAmRUE+ULWlwnba4ArcUP10RRFBaAPY9Nv1oyv6lrmm7MRFNM
9v/t0ZP1JnZ2AiCn8lo2QtHmdN1bEzm9mWseo1hA24KPaghOEFGeYa7GIGMw+ek996qpLhhEobHg
vBaFO878F4Lv+bArCJtkHqznB7OD0EDteXTcbfXJOiiaADE70zJu8C+rAPuvlYQnVaVOaaZdi5G+
rL+yU23Ed/MX8gBI814b37L2IFE3icDWJilt4QKTth6yrKENg7OMitlvy2i1iTqt9EChmRiS/VOD
QxCJyGm2KYQBS8la+/0jTM8FG8zOFrw77Z7kM9siPzgElFQQVr28bzedO7qewVLBHRRDuzCXpgu0
knRHe7hqPA5mYbjKeAVK6aaMHTyuhxAuZUdJZ9R32eZMTyaHDn5t5fi5Msqn/PbWxW5WAMDzcIDQ
bcH5p82/AQ0nU1DoJk5ChM/Y5R6BadPSQBqHprRkTI8+sHTNECU8BEoE6sKVMkXggzJ3LMRUuKR3
gV3gxkgCHLKv5mJlv6PMHLkNwZHZnLCeJOAMF69//hJ78syBylfDY/PlOaLOLBiqdmqq9LkhzqZu
fcK4pQwdp8AIPTYwGSqF9VCMsJiGtbYA3aBvzpOLxv5RSjLSIKKAXMGggJcL+QRkS7dwDNUjTi68
Dy5iiWPv0cKGhYqc42XH3zCw6wFb2YjaIgjVlAwHPn4bIjkOdzN90aKub3glPkPdii9B4o0W1iUF
IaO3AcJXcC4BunzYz7HeOiscz3xEhuHohSvgZuqVv6mLN65+pMwtr+8UbkHD6pSHRKdxTG4Bzl80
EpZVUFzzlabcUfHQTaQZTfsLlFY0lUhUpBe7G/5Xzh0lf8OJZdSEdBlCtItbz6M6zCR7/8jEqedV
05whixirPIcYw1X7jW2SU2Fz+iWQpAyZC/jfaDSPeVIWxcZu4cdWZFAqmfGywUWM7ZVbf4SMui0P
o2Ycr9RLm7CbF1grspjvVO0I5OrMtZWbWJBsTuLVDgq+Re/WE5uGbhQdJcxWExyDviZnx5M/wfR8
qCJI2p6rkszcqcgTli6II4FpuSo5tGbEg916Yu0yZZxfsGvx/n4ws+1/V1Q1BfN+nOHGXw8XA6et
IZ4qnVkqVlUWBvieAYDCb4ATokXtzJgtB7/wimoO74XvjcN5qjdzA+tRxohlM0aIj56J8XXzQDu7
FGTXTWxClkH2m7jQ70wi7lwOIuslmg0w6b13FwlsNMGpgawy1Csqei+wFCGxcpbkESe4lgeSM0bu
NrwMawVsj6k9wUGxsOinPs6pHbycTe9SEVFHsvbhHOpBsjhcsM4rnuymIxcFzAhHJ1fmRGDD+e8h
s98wipZpm1icgxsBtzFp3uJQzG1l8jy85BdygFT4nvLwYwNVZELV7xs80lcaxLaI4sPmITndxs0T
gygy6ZOWG6mkE0NXh5djmORxNJis4z6I1GsEOK1ljib1pP1WGaIP2uF5AN/somRZACQlWfH3a0IP
idkPzlD9MSA1f6XetZwo6mHYCHyAM6wNgAKJXOiHU1wItfUTW8p/dZ88zyxfhJDwmM6zbaz7ATXU
pIvvu6s750RCHIV8WP2pHJpOE5UFaMZymc40ZREkjvLpGc1h701dpEJJJDxuX3onedFg9FmsDIpP
iLZ7+H0Dyt0OP8id2hCVLfEK87rjbj3pa20y99OHPRftV2pOeq8l4O/yqJw1L5NOo5K+J4fgNBJG
asx6vYkTpqSZN+Co+FDMFn6+Gma3PPgf6VBxPfo+JGizVFLABcMPyCFHfVuTamHTOyPSE6JD573e
nRu5CgYfYiCq3C1Adwg6u9MI7Hva/+br/Jcws8Z5D4SxjqKYZltbvS1ChrC280/hOLwFgVHZOi9e
L6/MEgeiVpmgL1iHR54DdnuDz6ra3QrVyz5M+u8tPnEZI00gAO0pIjlFWYzHE5/1PAE4f1h9niGF
lROaoXKR1NmOaQSNtfm6nYckD8dElBgSoAOWPk9iZzGg2Y9FPpT3R5cdrex+gnQozXUGBEdBfn8D
1WYUm3sv+g8hjcgvEvO5E19GIdQJtWlPtpCNQzyRfQDM+2xztIaSXIkOp+Kc3TEAt2O9XrwSzXAj
NqTHGdlrFcnW2Yo1cQ8fdZyj2wrZVQ8+nq7bD2BuRMzdYx1KeaRHVRM84PkVh6QrHn4Ob8eiFsfb
9oDgZSJi2Zeksrrex3gXXM8LKaXj0CKBO7gWfq2ms/7HSHh5SNkqN6hvxKC9iK6lgkK5oJjMmdXX
8xe7atCxSvLMwFQ2qnnFQCCEZp7g57o/24Z/ZerYycZ0JSpPxarwC1u9zFm5gpqQm06Nok8P9qPg
EfB86Wdj/1eqwUAwNgkX3IcGSZ5qgwxK+SwBPy/Vx9YnsE6358vSJWFx+9u3P2TzKKGW/6hSJtoY
L92zR8Jbhk3Dchu6HcD4n9OkSrobDEqB6NNs3A2AuhZVncI+lnCrBAkVKEKgMARHwM69Lzp5OQ4y
ZTZUCfF1oMpid0ZkSH52hSiztFRW4SaR3DcpgBiDhL17r7DRsIQRybPbxnhxU0f+8Wmh58GpOSZA
oWamymgzvUx5ip4FJ6FuIde08SMRweYmgfTNsf7fd0uLN9yHwyQDXqIzJ09do/ZWdqtYHg59dqMb
SuWrVFUKgpV+TlzlpfqwPx8UmjboFKqOqRa534L2amQGcenGIL0FyBGi4NNo7IQRzN4BWkpsOBin
487x5IvrlgUhydEUay+f9ivQUiN91ubzhkQKORJr67OHk1FgvBkreS1F9nNVfEllw83INXhmQcuk
sxm8qIwVVSrBx5nqfi2e33ZN5r5/xOZKW1scQKsHfIGgCORVjCjBnz+Jp8pKWiNQVT6FL6Sy3EW5
drBRrtYILxe+IiMeUKU6svmiI1pZSbvZYSpl28A5QwhslBiyrFJoOVL67dzrVKk+6Sy0dlQntecS
GhBo+wieOAuquNeURiRIGQrxaAHdgkudTuOLV/x4R03ind+RxbC0mKLgCz3XVLWa6DhKZQiMajak
QcsF80le5+DamesLgd6qMHjJnqwei3hCg95k9ac98CtSz3m+QeLzJR27NCrg5wEAZlFw6O0vIWoY
4Ga2H6uJJsOz7jF0agKSuID7CtSDiERCembZqdEmH6pt1dqwrfbEjXWbFou3P8Sj84JMmJLyqL+G
wrU6w1wC1/mBa6l/kRLOHQA/HIjCf/lDTJQXtm7JI6Ns1jDYmnkd9MDRJitLI4NdhWIalVj2KCW4
qiaMtq4Snm5bEc+7lsIrV8d4PQkdiaBllFhCYprMOFviR7cYXYkcwCMn2NenRavooGm8csAlrUC9
4nvGWVwNODBDOtPu8jQszvx8t4NBZ3FODYAllYP/n46pLeZrKfMug+jSkcn2a+VA4h/gujdF7LYK
iJOdJXQ9vXd3cEKzZvkj27ACBZmUwPLZF5BRlEPYgZzorgWTukrc/XX1lfZufJAamLonxudn5Zbv
+NZKssuBehJKmaaYwIE4ik7I9JzUuowlkV8dR9fXscnClq4lj5PlcO13UtknaOjx2mlXAKw3zZyO
fp8P6kPi9rAuEegeQaDO8Ju+xkhW65ceFef0ZJNe71+DeMs35B+kyxDAE8T1jSONHKuAQm2VxYtY
2V33vEf5mQ5s6csNnCJGrNucYo/Dav8NRd+6Oe4MD3KqGd5uLrwhzs2XiDGY0sQIWEdAk3QdG6Hi
OFIFMqh4GTcwBRDWUBxmSyIHeONTE50lWShMbgeqdJBwbUhAjylWrzd+KRbtH54zEHeu+tOOoNpO
THjKUhKetAktPlTK/3VlZx7rcREnsJbJy6GmoqLHtuEmN963GRYZ9kSyTNHQJ/2AXfIsxQbIHDIx
6aeWyfcnGJmTDQILXeeyolwJpWoG+wXvvLJN7aDyM9fX3rS2PTY/mlWPELlv9Iz0uuL7dYOoJR1U
CBiAw1SuPtPNR3Un4E1M0TWUuUyMvI/C6qZiqvuFavnQuSZ77EycnP8Uwy+dnMqFs+5+sggdHiuT
b33OzpdcyxwWKPMZ4FwMxDIpiCWa6xwL5AZcfnyHvjHVfA7YTB0rjRDJ3HrkL6iAVmrZhRTDcz3d
li/HEEyV5nMILlZefp2J0ZNnlGMD0GDfQBNHoGLXpA7lUO31FtpyAQI6b7IIcY3NS8sw8TR8nAZB
7lbrBRAJHJbYXqaawDh2UicPDOX8QveIM0UbmADTvPVjy22uHIJx2jh55PBRrVt1kslVWNT9a6OO
Gt+1RPrFDbHBc4w/adCIAZUCX9jIB4FsKnm4qmS26JuOve6GGATGm3HIxn3FbsaWJ36waEMXiIna
heTh8XhxVT2JQ1EG9z8Yx0LbTY2JsiUEPznuw8wOjHrRts4L1IkprWQVo6gEhXXrPFSb2G7LNiLk
JXLHt9bwvF77sp8tWWU0VIY2nctL6AzKC/gIwiRGrDwc1ZosI5F4WA+HxBaMIZSM+/iI9qsRLyow
zrkFa/eBLy7AE5ElXHrTaJ1qxuNWADDr3Gkl5uwM2U+K9iqEURS6lbeoskL9B30bj3L1Zi6rsAAO
k77bHVkgj3runeozsxBZPRFs/4RodMYyiA01KH+ffybYrX1Nlkyk/B8hOe59PniTpLZxge41zyV/
TLLu24QFdOM8eVizynNbliBcqfg+eRJoUx76hcehf8moMIJi5P17varJQQUzWo3lA35dqd7qyIkL
gsgy4K/3KAoQFhVP7sSEuymHawbcQ7mNuiIWrtAq7irxoKJ4v9YOsXpGQn9R9Ql2g3QjGuhlHcBU
TR7LrfMo+DrpWcm23Q5v6foXnoOmnG0WURRBYoAzin4Gw9OWddikoMqYzFhRzZcPwxPLTYtYQvtr
fMT/LFXGqbjVXo+69bMVjwZP2l8iFiPqP7cvHnrjf58kWFV/gFiDmNJwhDvAyDEc8d66lDcejPIf
dZsEhkLIP0W2Xwbw6ziKxQG2HnU/v7jSHpLKuzIcUnzZYi1hwIUlqnZImqtOSpXRBqon7K6l4NF1
C0NkmE8rzrsuAMaHAHMcCfSn231AX+xsvsXBg31F8uQ1xj3n3Zs7QzZ4QlcV9OPk4Vhh8cHvdCsc
OgWlbDyhPHvF9JuLN6QCx1T02zXe0AYUxsCdQNnQ/1dgH5HcfHYOBq3BEjmqQoNkN+pU8AFWcU1h
jeq4PH8SkMhVSx5ngAR6nXkUcfWrW9Qeisg7YaQae98Oynxy9Ju31LbMgvC/ff43WYbrYpq92kFj
iR5bY1uNJVzLC61fL/vsbuR4Us3wPQHBb8AprM3DwITz+dIXplZdcBEgK5+KpZDs+lDoOhkg1A3b
ru5nM6u16e9Ah2N92cmmAeSz8YQ8efaQ4M43MlCB7qusAPntqJk6dhjJzVk1gzNXfsDbsyKMBmqu
QayoJ2wkdcIaK6ZHIk5Feo8GHKu9563x+2KKajdP9ZPeynDmqGx9qZltl4uuiakyGlWdWprVrjAG
dJFvWcqM6VqE2h7qj1yjsGksycyHop5SFwkyFN5Klk3nVRlVju3SnNr+SZUqXLb2ka864EPr+8eG
HdJp4v06cNrsOiQnA7CodbRRNWPdCnOhnwPPoval2/6kKtB/ssVxskL7vIxCzJ9V9VYrp25uMbRy
0cpRU+OJbOMymlBq/9gA88474YwkJTCbqwvtnOVGOYq22gHRn45T9LHivhwCsR4j+XIL2ytub2ac
9VLtj+BziOHMnfHNDZPIg+OlT8iDjjKIiS/5VUw4alTYf13ozsd+/2iQxmMn0oDEuSdm1pSdaI7w
P9FwSSLMeIfQuFPpmwhMWzTxTgu5dnLMvqC8i3b49Ng0BE8E/WTSYHI77XV9vXlHxiFOL1qyFfHR
Pf5gAtPopYhAb4VZbU+Rnv/gJphzC3kPt13A2SVzVj+wAlSf8m2WAs4WagzmNOSi5nwQX8DHEQfM
e99bT5P1YDCexjFejMQyxCNN/36rsXj2ksWpad+j0CSKBZpfIQhDsClsXk3zDGO0q/BUkhqzSaNI
3yN49bscICgvjWmZF4OwLYqKU4GwUzOy6e5iUCBwVwWFyPq6lEp2HD1sY4dmszboTjN/oS7EnwQG
HEdj8eIoSE5T4ifvysJCFDyo/bioE4vIkwdQkO7chLVsYxadVvni5/SQNq1IndkzViP/hp/bhmpk
hoJy3ohZ102EsbZj8uN4oq0sG30928l4NhhM+ZJtmuu0WI5EaYaoUJPC0J9GJxSJrV/sX4exQQZ+
7aNy57013RWKYrkFuhA9jHQvCqjYb9VtQwhMUahrehgyEoq9GpXlUTe1Zi/7GLqO2BBnDgP56yZS
y1mJ8xXBJSqLudc20ZN2kLRMc7sa7Z5gn7CDl1OMUbGXUTngi4SiVDcDxvbKZKi03SlHUR4nPt3V
NuUBy9mDksJptm2Tz7y7jgczfsJ5Jn3UE6KxcrdKYBMq0rdeeq0qXLn8PWmAm74SNU8gOLYgSI5N
FBZTJyH5swb9UtsA/0wHgXvIBH2lEVwRKYblXdEi9sUhmY2NQkKnmKr67eUjabU4VeDLukQPKvu8
I1rtFso0bnyt6C1TwYxbDxes7kUHh2l5XyZOPdzLJrfE0JAfd1puYu9qMgCnAUZ/EDJfBPQPag/k
9VmejH9pXO6mTNlIbl9tmcVhcyPqnMTyYkdOL1ou8a7OqVHe8YDwaBbiMyuFUmTfTmMJl3HEj7gV
wc/LlyOjkBWgGL9ff2lwR+nTlEgHRYeNJWA1jhFXZhdFlMth2bzaghXGDmhuM09h5ISRrBneNysR
8n7SQxIcz0ElMGXjlq3YgPJdqfAoscXtXWEIilCmG56minHv3spOg6cLm2SAD9KfdSB+75ZHt1aD
B77xyLBdXUuKOPQ8EJhvg68pj4IyyB1+u7EpQLmjFvceLfCg/FvRW1NBDE9uUdJkO3yWHs5liZiE
eFyQkyc0RmwB45zmHuZSR2/HO/Qe9vVJbu86EoaXJbM0kFgRAhWiR4D2lqc+siiRXRXcBN8UEnIw
SZIVj+/9nd59Jyq6nbJaAJWHFwOY9MP/TlE9fbRSiW9KgPfadnGkf61+b/P9VdVff3A7whqU8pAV
0FmcWrE5xmthASsw05/W6XcTQc6Oq+DufuSAvD6sWsMjuPWbJi79qN6gVXCQmec18hw43XjTpx/6
jTCWSn5/xfx+RKk6Q44T5PS1796UkhrqbPyfZTQnwHNzgKg7iUTPhA2dXe5bfihoagCTu2TX02Yn
6uxI9BHySaj2OwWXaAdtU6EEcPD8TLtkh7e4mWmEkTWZHqpNle2qNGZ4wgMRqy5Ts/nXg/+y+EoK
Pg1mw+YRzbqpzEs00j7igd6l0O9HJqFSpcIUaVzqG//yUVc5rSfdZgl2QJGevXEk0CkWbfzm6PQ7
2949FODn7AXyKcwehm34QEaxM5eG8ned2kLfJzqfwaOvzUmjnfkRH4TrMZNg68ZHN0mSXJQS/gIQ
X5fdyN/sqbSW0pS7v10aoeqDZEsVyD75aetlXjPWuOb6+nLVflWvEY19c7STOBrIsH3Syo+0Nu9O
RNQz0QIOVPUF/kqyLhHq7n/jJzf9A/FfJPCYPT+UG/8M8SDno0qBffTVKmTBt366Jzaks5t3aUpW
XFMiqB9hxWNQ60UDp7yQezIKTOFizgVCCnQ9c+zs4ce3PfA4mztOGmI2wOmk6/nQZ/PCf8sdFFpN
l/CEiIP/637yZyWNWp5QtBMTjjHAv+Vnq0vw/TCNjKpdY5uizkwzaLOnBFq69kprFvWUHtyZ5zX5
jy9NZktxZj7RXC0cgALik7sfBxIKQ9FbdZbhRqGoEi+6YIQ842s1S9rniSXF42OrgUCTai1mIARS
VwAzhLyAyLYE/SQYt/y1CS3zz1r2iJbQFVzvCBMUEaEpDXBgC0U3nQ5wDRd7AZpfYRPEK5nxdYSA
m5tG2x2zb22agJDs9TfIENoF0+v4t12c/eFktmKVx46bJG/Femj+QgdWKc0OQKJP4f5rggJBSlF/
otVx458CYi+i+L42j4AzRwATTu6r/h95KAn0dgxkzMHM34WvHfns4I+KuDkVXLoHOI5QVnhXxgjL
6QQJm7Oqel01f5gFR8eWss8lZB+BQtuVxOIwb9DjhAjVyE9l9Oy28x27cFtDOgvp9uHWuWnyo8oV
PH+F2PYUQSvc2vaOHegPSYCyLARsm9/XEZDK1Hai9acoNqhHIZtZNy3jW5qO98RYCsO0kLoff26D
H9nZFq7ZHYqChyuBz6vI3DP8SYxJa4i0Gn9qVWtLA27yzVlQ5b5uzTCdWnWe0jIJVv4wcqdsUOgg
jQPKtk4un65UkOrgYVkctoY773quodmC7iezedweprrabQcnEoWmRlQNPkgrHf+AeAOkyaWS68nC
BKlDiVPhnbXTk2cWZJnwgvNMnin8NEUL1/dlmo92SyyiqBvKmwVg0L0AGw/jaDGdaEJQnIVZ7bUA
H79OFMHXjfvno0ypqPtLgGiTVoh8/zb6grGXYPEnUd85XcO6i3uvyAi2BnL0e419cha2eDTfd7BU
do/EO3MplAb/CKXihCFp0KDEFPy2klVeIMFrvAfky6iDsYy/o/i1baJXhway5aXvF9ZUR/SFjsW2
r6ZOcDM24dUiHYCupiOQsxLGhR0IBZ0DrWqKMj43+AXA3Mn74pRYSoECGQwwzgkG1QaC3clultTV
jGvJ2nThAVBCNymDfWwYiZWcZs9VLnYgpZZw/4IUm4143MnNbfKuR9G72SHpjDMAbwldgiNwqn8Z
xSa99j2BPyt84VqlcO9YLxPyIDbcngJKN0qhi8PqVV4YZz+NbV3JpFMaaBRu+uvFPNE9IG2cZOlp
AD5c5sk+MOmlS/FnmXAK+nYQr1vMHQh5t3z0RToiCViCBd0dBHuYPM4bXgklS4IuG3/WgeUcPm9g
NkhPMVqdEBMBmPYP/nu09b9Nfca3RwtGXD9yREUb22+hFTBqL7BFsaHA7VPDO2Rtxk08eejrJLoA
B/limjs3C94O/4qrbBhbaCo5wmTcf7XZUlboGadb4TuZcIg/2pSMJVVsSyT29DLI+m7uKiIK0PJ/
M7Rw26u6rTTRsloz6Jo+lYDHXpPYe+GPQvaTdyDr5trp+MIaRkI2/kKjPDvUFA74EeiUcXlncx2N
xXcOpXhzJdQpFGZNGo2BCdz+h8Brz874q2TWFiUAfC99udJACjU3ME2rda1QHSNok/HsE0PwVOmk
Fu0WHY7nnS4jbH7rG4o00GSiRrgeUA6i4O6/soPx8qft5k6PQwEguk5NjniVQZvVj+yfQGJM0sL+
LEUghQgJ9dFBXOr2GKvUC05bmuDOQPJyv/85klAU5E1GJinkO6H+ccXkbTV4FeIyqq2ZXRDjPzIu
2fax5t/T/O2CeDuHYJHYaxau8gjCFYHup0N0ODCh7Goi8SV7CL1HcC1Fd89zHXynWQAMyGajXU4k
8m74KV9epSjgMC9LkvmFQuS1xgBNeuAhRu5/i6kAQshL792Nn9b7JSLwHEzZpBqY0f9R+Pvi6Yf9
OubgV7xZrKCWu1+JriVSRw++Fz/b+p3f2kUrRHpcT7Trwb//siwujnhLqkDhaNE5guYVihvL2fbU
aBgbegZaEL77lH+go/EHsuvsMB15VzWdFegCrSzZXDCWtmctRZS8QfYuiRfpIxEoOzyoKlm/iIGR
ASxuUyABWIt2eQQc7wCbDQodBiL1MujrMlHtcNuHtoWs4lqBSsojiz+q894gbkyMosv03YT1EeOH
jUGwvwTmDU+WbIhWWqLq2b6LnHY4+B0FmYzk2/0WSipyD/Y3vndKtCroJ3x8+srOn6Njq0RK8jFQ
l8Bp6JKThxbC+V3ucYZBFu7FmHeNP+a5nqiJjtnwCSIh5cRJHkkGBtEqfcrtsbrGLfLpaxbGv/r5
rW895X/Ukjbap0Fd0BNSK7n6qT33q6CPebNY6UPDfb6uhScCR2tVtSaWiCk+txhGH3mvCl/TFui2
JNmJN+shFq5mqBZTspHFf+QArhw5MbGvuu1ciYXE5WaqqHDazZQZoCLYrBfbzm9HGKVzYS7DohUZ
4SXgi2o+uBc8hwdLntYujNiOnU/hAZ6yKqjgMK4prcj52AkLzYoaGwV16mKmlFbceVCR+t0GL0nF
m/Fho6PkIY6bWi0EOKmxOxUCCfo+2e/btMQ+OADFOnHpbU/lXbaHKzzn7fvzL6obDr0Uehj55Z8K
wF49xsLowzYDas+og4erFZLoh2AjIcKp9NbYfRbu9uuFmeH9h0KE48ZkTaYIPLcwweVaUaWMZn7z
6XdEWj+92wzQBvN8bdDbZHLJP8DrTNeE3NgQZAPotSdMSiecXco++NPcZvzKYVmE6+pN6yF9hWtZ
QvW65kFpxCCsDyIax9SFUvwrzXj+7egO5uDdUT43VCqk08oJECGZgfPptkXHguKpPRHyYeEednZk
1sehZ+TAqVYT3dgv8jdknC89lJVqW5WIEuK0skETVChuK/fXCR7vq3CqfpXLyvkQC+e359hrjT46
c1QUr/RzPx9wBXR7W6euDq3XmomK643fcb/TaxCzLE12CAIAWY4r0bQbGHedhTxpQbgVYDTs0IV8
XK4PvVwYLpecoueBWZ8j7UdMNwHVefsXtXWIUtsun8dZ0PFDgl/+5GF5EcjS83cjwo9i7+W2ImfJ
+sT7iLkJi4+vLe/qYc3eKmp3HH5Xug1y+ABsIec18yis11fsgZCsE5LYXcft0r9L/hjM1SQC3vcq
rrRjYlOSDcCf3qxKpwTcX+Ap4+u19xavUz3g/RpkwOp+U1Y4J9JAaL5t4RejywYmtuDKo3wl5ES+
LYS/1jQ6XTkbYRYq4qKjMqatyfESVYqkwm1ql3L80lY6sqdSsZS8eWwRWKhjVEnvTn4Szg/bWSV5
88AzF6qiEX68cLYHtycylzkaSGiK4O1FKLLXLBmI2uwnqiZ4trSDyPu2sZR1nz112Wwz9pbdJMUf
1KZtfwlbAVj0D5F8yCtDBn0dK8m3IWRXFVRspwNm0kOw1y7JHYrUtkbvoobmaB4FeLolxmeni8oW
IXoGgvGLRPjz/EGl4V6kKYsdM38uskZZcqSkT3v8YVUBsFmWX9UVskVczZA+QH+16kW80D31uXK6
s9M+ea9PeEJ6OBeT4H/saEjI25gfcWx1TeCUJ9Bn4OQWYE6VsOGvW0fvhKuXVvQKhCEsb1MNES0A
lcEeb2Dx0lfkr59HotYuEyLb12SWJfBuHYdxZEZIkcFTTpQD0ggz3carLeZFimCK46u4bxR0VgCB
HhRMr7kWqWM+W0cEOhDg3zH+WhUINmFFbgOMxwHqk9xF/uLjkylnqwV0eJMqyi/46iWP9PfnFQ3O
BulNGPuWaTMLEth0s2y1sJKYg4u1zlPrsshFo4W8Wzwno/rBYmCQ186Hz4arkvQCXhWABTa9ojrq
nb19PAsDhdrNU6lrlOs/irkk/riac9LJFvF6kQ2MHoBr8hArJWuOJfKoYYGBMcLjGphWGjyNOosh
ZLe8X1ZRn8JMIEvMljB+1OFzJ1hsfeCvCJDcVLeXGJMcVnNLXIzHNCML9UnF88derYEjzRmmPk5N
McAsU3jc1uLopb+gmtRakze3kPM7++bd/q08DyU9TKPmdca+kwWfzOFGr6+imVfc8yUBSNlVeUto
10jwv/IgfClaH+RJZAL/qgHXC2Yqc5QsKOnvwfQy7xw/xDEJb2HgBLfpnMjC/gt7342vg747wtq/
+0w3JKWG8unOJ4UG8gCv5pKZT3QlhshWL88E3kMq5l0zfZgkK5tD7UyLaguop2xux82OrNttaUMN
NdKTJLtADUEOThrNbLdpPCbzabSlHE2cAy8GptPd52pH9RJWFVsAVLvDHAaoYAYbdvQtssHKce4B
eliXEaa/v0D4omX9dzJBFfZa7SaqWjQAg5fpX1dN38P2MAdQ0yKO4FPJ5HJD1IKmqgwK+QvDu7v2
czsn+3Afv8aJoMG5f0QlsGuZvo0iVFHnPftsOu8bpocFAhOMVbwvl2VeLtBnQ4FIuChvHma90Vwo
EIoI8WidGSiGS/I0LZ2Pkl7rK5pfv6OdRWOLgvrJiBY05EFVVvITM1ubZmYPDSNjxp/FTODriZ4N
GCXg0pM+Np/pXhJ7K4H9OGN/FxLVBn8BEvQ/wTkWx8ORO5QLuF2KMexgSOK8dQSfVMUf4Hq3CpC3
xEBSPZRX3fv4km+1POIuFfhXildO8My1AirXzReDTbrC8q484TlrxGjjrrqvWwxoiWThs5Jyn27m
yZttzLp3DSpP4f0pyj9o3rIa/uPAiBQh4ASupd1skJHrmthi22fjg24Y+6c650innOnyKHAbWuh8
GQuLNmwxi9MP4HRbvTktQ7VRZRKYDyo4JO412kN6abjHWjilO/4RShKXrA8k8umSLZKZFx6derPH
mn0f+fomAjizuSW4BY/cdf5V2hUxdItVSRvnuA+FePXQ/2U2ec8GN5UW8Hxd4rv2F3Pwe9WwNQL+
AVP0V9uZJb843wnfILR6lIiZw4zE1vY8ydlsTP3POsj5FfeuzduOcDyj+rwYJMrFLCkrYPyBJFB+
ANHKZh8/3CXzZurK1XeglEfrmyjPJMWiVaXcG5Zhfq7LjN+L+JXsYCiNsfo4djPstWB18wf7LBEr
KLfHZSwqLhrCILDbkbyS6THQ+9l/4xGnknAY1do7I+fiAx6j9aQb2/4Ubs0ZSvFgjxVH7J1cbRsq
UL7BdvPvvnLUCE4/Gly8b5xhWzhmCCi7WTsLD6G9VVJO/xubfWlzkTZPY//JgYTv6A2amUJyWfiE
Vy3YpUM9mxgW/B6JmrZvIe/bNB8cGyL9+/4lzSb0kw6w13slAi9PLVZaupyLe4p0cHqopC11NKBJ
L3xtC1ynPImffQ+LgKBAqwmpy+y2rRUnfmBWNkBmCHhX63XiJlfLcwCRagutwY1RzUjspWgM0ds3
8a6n/DEjlqEzJ/T5KPxEb9ZKXW32Bzy4Rz+zvYGrVkcEfbYKWjfHGqcLuS+kFhN2LutHsCUWFbIm
Ze5MNePHHb+JI3pzPHfZ3PR+FdPJWntH6Y4ZLbEMKZLQJ5AVu8k/kfqXcZUYkJQn7OC0iXUgkFKo
08ljLBothGOvw10lRfAvwGDZATdqMEq6i7EXyUmWkrQ14yPxt/FK7PahpSzUYHEi5+DjdCgBCMH5
z1MRoxRMw91B6+0E7x615pVqT+siCIpegTHF4bLdeODD0UILuLk41F66rdUF4dmGkQNW1sN0F25A
s85KuGqYbj1gPd96G0cT6++GEfG+ZctncgyxK9XcPXmpFheQlaKn5Jw/5suq/yCpDTDvrJQgJzzm
JVfvdo9qLhJuFBbUtvWvpCjo81FnFhpsBMyt1dot6ljhbf93bmcBeSneHNSi4IEbwxyRWV7MHFL6
V5rEKpGtgSDRnyEmv7OJ/3JM1swsWSp4DNlyZA0HCiclAkRI3k6DJTJsAUEEHbpR2B+h3ICkPDju
+aQHlVjHUKAtT2QFAYfrpwcZ9WSxmQH/632jBxO5FU72qlTLLgWSuo0Yuox91hRN43F0hRbKgB+u
btMVE5HJEzsP7wqhXUJgTGo5OHJPS8L/H/nLXUF/JibhGo8qaSu7NcUq0h0im09TB4Au5MymhvuZ
YMrycTlvvjXdoXlKx5/6sRXaLxKULFcKEUxXVbDsnKkkud/p7q80M8NYvoSeK/179PYTNivsBTHi
Lz9un/t/9FsQ4WNTpFvx+UQm3Oy7V9dzVsBu0FpyrAplM92MiXZIyl47ZYjBxkoYhNJuDFROXAna
PKX+jW4l9RGXG5lptQkgkzuFRc/XnnF3cTkltNkVajGmxe5EpIT6qnMl/1rtXIA1kpu8w3O+X4bH
5t17JnDsgLHUm+kAmOjjuZneKSUbK6I0ZBb09pdt8gyca58GRyHb1x0v7CmLB0dxdQHqNSixmoZw
yhkohsPXX0+51OGRYic3ZzVopstLsPfSsrP7Mq03b91DtYDbATe7l9LTl2YiR7DZm9c27XE6zt5i
JgghKh0ntmAcN92Rbcf1yVGhVgs5jIP+GlM6Z/rocf8CDngOuAgJmjAhuaLizq857Mskqh93KDfh
mvZECO6iUHT1cLndNKqkQY+SszuF0Cf5RQRL+QV9r5/RUxr0j4KxK0JJb+gG7Dw+JP1Ld2Ez1nNm
CGYnUKAoMzkRcSwLQOxZgGDDzldLFivfjve/fXw1WNUtnh0mzWCtVqf8LUTl4NDu7T1blUToKuSX
n6vymvugBnMZZZqZweoJbxt62qoEiwAcECHVhBZHxrJAiODdNeoEMmuZURT6oLwNoYQWFaC72avt
8KRZTvGj2DokWcYLdHqm2nU8uZsNj1zSxZEH1jcaZayT/uNpwdesNQOgzJcbLRe58jYpCJ2X7Ldx
b7FuRslJUwtG8iECt0sPhrxYaW2gOt7eSQUomzPkofRpAHh3dsdGP3P0u/rn21G4LtU31WUOicG0
jNddp4KKmHoDoP79aKHsbk0mhWbowQ1G29OImA4Q9KgJddPN+qEuxIClHSOgGpyxZ/ZGv/YmXoMn
XcXiT5d8D2CpQOSbOhm9m6eCS3eB9jI6F0gSmTpoG3QcE++I+axdUA99HRPdhLjLSgtctsCP8SqC
XCdFMD2VrSgd6mFi7abiXL5D1cnrQ8jXetYPJP8ocloICQ4Z1mEx1aZAQca/Y/7Ljno1tU+r2D2B
jhGaBiOdze38ryfWW73aF0e/46sKaiGPBikw3gjdYXIyossHpMgPiaDc2YD5nbabAXfAquYaLRtT
ZT8R4G0/J0Po48j3ci25Q0eZ83nvUrMgtz+y3PIwWjJy4XTV8JSSIwThGWxINDRX33AninUgvO3e
HdgrGAZ5yjFqdGacnTPy2J3oTtx0eKlpEN7dMgczm2Ae0SknfM5+J2Vy+vdPp+frS4e2A5FqP7A0
orHOJ0cdcrt3AbNOACLp2U0jBJ29kWBP7XP+BPPWqWk0LSNs+8BvVTzhNqrNd4XFFIXNiETOjwPS
7jzSPIDz9J+OYCQpPI2RNBdJDpZf35xMo1vCyA1CwPYzysP7jWMkeGynQM0vfyVNi19OvcaRqpUU
j5DUpuqRvaMJoY5NCsNmpITXz5/YRBSsm2EdzNJkCmruR7ow3Z6r95X6TPHlW/yfFf6KfUbC+V5d
hGrshRUsVCjvKLDyMcbyb693OfwW4pnbxt/n8iCQcf1fCtNoEDSNtmG2GUHxS6O/ZBFnZ1+oqHyd
+4Pq1tlsj6mBMyMsM9rA3nO0kzch4GzjrIjOLeMefbKLnD+NrTcjxpGoctOVgUi16ixth2VoX8Yj
N/x37WioKTuoHepp3azc1HC4NBuYBmal0S5k5taDI0JIKVWfd3k6wQ7bH3U/ixVkHmmL6TKfWlfX
WdOinp4YNG/Rl24qSPMxgbSuBqKjS/1r3lBYN/Q8GXzl/AXF1+Cuxok1LWSY3Zhri8XmZlLoEbX0
7dLotjqgNmOPp1RGGx1ACVFiuvVimUnKyiAK7OOFlt6t3JebN8gYsHfynOpIQD5yZezFWIpc0Vcs
y30uW75uN9pyQn4EgQS4y9mYvQLWwLhwlf60lSbqfCLHlLa1md6koRehJQewEkOX69zP3yFGeIYq
c3RqVkDRooKoziMsvABnpEwjflz5YKuXKQrR1VJ97kTaI6ELfPe5klpddTUKp06GE0UA+DFcYkgz
y9LnvbPeAbM4jz3CAHFx2uWi7MBdwd81VSzuE7QYJiW2dOUWjxrN3hBUwJt75lLY5m+VxPjzMDMQ
mTxc6afmTkHdUNE7ITrOXKMmpBHmPfk/XnGwGS8t+UHm/2R1iRUQ97IchSEzPQD5cyX1L0aJZWQ5
oNkvLoKw4JwmiHYUGbkwy0vpsN1e5zxEIFIyNrkhueu2Q84f3QxIq+5NAT5W1dVWMH3PLGkTshHC
/+rp99Mnfo+mamc2LkEAwtTngwH8ROwLevXb2gVIndvLyp6GJC5DCVb0pHiouvxcbFdVli0zJcjp
MZAvvpw8S8nhJSE2R/yiDtxyOuzDFhfNCrSrNDzaUZcN50VqiHg+t243wo7+BxPjQDSgDcoYiIIq
iuhAOHp5vzHL3bgq+w9S8OF7PiMor1SsCpJLP/WNE0wVe1/q5ykwc7kJS2BB0pmEB+xwgW9BPQj1
OQOB+4Ef6qR43nKYX81ipfDcdJdgCMfXXito75Zu064Mug7Auys828oxWEKwnFQC4T7l/IWu/5xl
9z2Ag38gPgTy528BIyA3FtkNydSLN7w4KtfLxk0/1/WZ1kb4OEV8DYnHoEVAe2ix7XU3+C2PkaRQ
wyXELsellqpavIE9Ug+vRMDD/6+KrkSSZ94s46Bgzz1+03TkinpJZnyvAjp9xBn+Wi/2a8/uuPjR
r7EsSWu514dH2ygjZg4cg0IWwCBhirj4mBqPZsJ94T1cqD0FS/6MyoRYvkyVrxaM6lEwJU2aOJa4
EMpEAys9BzUED9cOENir7AKroJjR1mrxFQBJkC8/0dHHO9KOQUroMKMlZpi874S65x76GdyVjw94
QqTIeMUfjCK2K4h1+pEgWu62XJFXUUDMGI/Nyk33uDxhy/R8gLlhXfVykjkNPN17+xVaIpU/g2ei
ZlmBAhusLFiBWafKPiYlXfEMsFpL8FqUDIghjDnLUgfEV0hVqfd6J7SQUecGwgoQnDJZXZoP3NjC
alGkJGfQB1Qg0ZPfeJlpXw3Qd9ppm8cNLt8JCsm972UVAHD+hN8G7VRLurineKG+WLk8gKVIFgfN
DZby2T3Zh+3hfaH7yEvNhn6o1/Jh0ShS3GZzXXnDpvHUO5PtX0OTIc+b9J2ykRfzG/8uxVOsaWfT
2a+OGm3YV0UkTjHOFYA8RHGSlu6phfJBlH0ySU/MbigR+aeZHYiwHZUca4oBpoqq7DKy1VgUgtPG
OWUbHWWNfwOZgmp49A453OAR3CfeZbLH2XbTRTEMtlDvObUhhb1Dl+lM6UV5VJxWIOfnUq2tPZYo
sLZBENzC1mcAgqZpMIUmnkFY7PWLyLCXzPLGGrqytdCz0uDBZxELoCc3Qcv3wUb8DQticFzjz7Mc
cL2UP67p0TTVoisA4YtmDwyslG0daJNBGIJ1hgu9K6xRNyiahGg5pEfCyEz10YowiBlCLL2WtyEv
lYSuNjLXFxpqLivhOiOaaxEZXZVURrnFxIlnjkh7Z+nZrTR/McCJbdd5w7KXNC70aJkynzBqVW6e
XY7nIt7D/yiYs+QeBjNbAvdZcWb/MQaKX4Jbwk0BdOBKmFcgIzcAri17yixSsi08tLjTejcB8Ehl
pUlxsV3eqmhFrp4zyPPvQZJ14FpmbZvOQiG6n1SZmChcMF9K5e90Pqi9jXO4y9p/LKRe4l9Qsqgq
WwB3iZtJvfvT/9hyYQL2YEJhe7Rtf324CRKqXki+Acx5aonFHBMUoB+5QnkBn6uYW9aSO1CVBW/b
GetxzBbjUK5w3SF+oiUGm/Paza+xGj/SAvsViY6nCItKHQLfuM0lsHu/rW1Ia3MDIlN3AGAZSm/v
TeEzeKgLTubLTMypdoC8Q4idajnTYVeCH00+54CLVooNok4rSNczZx4Mvb0p2oCdXLuXwJpABIqs
2/Wpr2vEymphcBHTLPXxJfia4EJX5290vqx50wNRv5IwtUCKxviJv4g+5+SViDSN/E5NKCOr+gnB
bWxX6GzXnkbfY6LGS5AwgFeIw794v/JRtuJjsFlCr3FZ/Lst5PDMI5oMl5vFVGyflOuKDRkCjYPv
Fu0eqEDvr9YxAZHGwz7CiOF7yaFJ1KBxOXRkFVrLnvzqbM9IMxU0rdbmw4IKmzLqVr81iCgOOC3w
IJUN22RrvNo23mhaPOd647fHsNYIRxvEGVJh9w5f9rxCe8GYZWgMD2Y7ZA26+y1Ms9ZupTe1Jn8B
hC1R6tLgd66BtB+iCaQZWJ1VFF4rOt7CzJJLBCylMofgDDcTwUXhNpNDhQEmOEKL/60mGv9f+EQp
ePHFEQNBiC9Egy4xE20NzXy5AwcW8LbTSG2wpzeecnTos+T+ybHs9FfUeDCYNEEjIi5/b3cU8Mn/
ZvmrNFylUsA4upf2Bqdp3R5RAQEg3zmY+Wp1DKJwLJ/sXQVI0sacl3lBTlW4eQl2khSItq00lYPq
RIDB0kCwBbtDBaOz3JWHt37wz1YDHXKsoflKIKEk9AVi2ZeAUtxVOa3JnJftDd+Rq5LQYk+pYPrn
MhQw4t2HP7HRAMA/cjLhEKubewiKM5px9sX7+CWV0peXChdnYQ4GfrNqG9xNDODtMY0ILU0kzKsV
LmgnH+wErknQzxSIb/i9AXH3rk/f1BEtYQY0qXb9XR/BosjtxUyIQcvYkcPNooB6MKIUasOMkeTB
m5/Z9IUItEw8BHNB9risvrijnzjSPYOoAZqTi7/f5iFyD+71HeACyGXjxSu85WzA74PCLr//2NRv
aOynLN6TKJeqxZ15wmwqb3RnLpnXS1D6GvIu6dRn/k3T6cqTxCgWY/ktXWv5vu//LVD6/1FzEm0+
WWy1wMO2puSKSFIyR2NxcWKihA4gK08xm7HtG6uBStz6Tfd2ca9xKDEEEbg7yjVV4fiKdK9yneFp
GlRlYzSPnCtDMFdvhMUnD88aHTMrhPzK6Q7ZbaItaITNQZjRHUeUgYjILMhOcM2+c0xeM67/ko1v
ERUCKWEeZXXuBlzl2MA8xk5TchhLR7J2JVq3PCBiVMHQwNEveInnndTl8ULLiINT6BzET//MpRbX
UUNgX+FtAAHfC9SlJejU0Q9QrIOWo5+dNyGbq4oWC2DvSJE1TvKPRJX2TssdjSUtYvjF7eiyNkDp
5eKcGFCB2hqQsjy1RjSyOBNBk153if5mCZA578AKrNU+mFzAJEA6wBRwjF/LBMnsJEaID0zAjAN0
7JoX9Gy4fnwiEYC1c9Buu0+ZZKtDiq6LVXRpgxpEC2fYkanrqogjMvqCx1nyfM2BV0cLqYqKHrMY
T1IhjZ11lKutYxXTnZ5dtARvY6glPOHVz+BpbCMZeKXvJTNx5K3hxM1O5hzxL1GKk8G7cm/L2KKL
eGV0JjR9BCHvkjBQXb25FwzaIFBRCgo4R4bmG0gU6LN3QjRF1szWNFb2BXp6cU0eCedGux/l8w08
6UCXBJd2e5/xDeYRyfmFYMXqc7aiOr0FhKDcM36tSf4BgDOOJp0IStXnRsisJ97vL4l4RdsMTZlE
+WmeO0O6hLVsdtsf8fggIjcBlzsVrlO8O1n4F+VCWf/WkYKQ082XTSgpeMCaTM9CH6vxHXv3gG1g
ezfcpu8eznx2eq0Kiw6oWMUO2AZku72GjBOrHOYZrjzAaZCbwQ7vkhbhqIB2UCIlqwEwMX2NEDyq
6jXQYXvOCXJoVMeT44VIge70ohRw+j3c6JFaHhltYNwgE4NF1bPbe1YUS+vpIkvtqhayQM28vKVd
lMS08fq0gwdVOR9jcIZTTD8wD6njoH6qORHDuzN/JTBrprkpedkkBRaPoyMYO1YmHYk0U9lI0eix
H1wl7jA6+2Z3ORF/lb4fs5nnm10EH/8goX6WxpKo909yD8EKH8FIa3awu75RqpOi6kaw4cZf7FAR
UbDWf3MhjLuqlZtjNhQmMOMgR1caZ/eAKHhIE7olOzQ3nhReigu5in00MVJ0GJ3FhaFhtwVuRbWn
sw0v5n8e8MY534z/1i3IEyCKrRLXKVk+hlf58Lhg7E1A0twKtJbKiIxxMuEp761piwRGDH1vFV3o
IzvKbvbTSwX5YtwA8p0ZTGZjbNwU5HqVT6q+P4TFpNHTROno/iNFUPzmfCKQ+MS+8HdNvq4a0HdC
VJ6sQ9/nRtDJK/wHQbmiz3D6vyAff3Zu0XyiGBX34/oIT3kEmFHWVNb9UquciFFEgEfIQyubCsQC
ZbSrPvStTPQCmcPr8Fj/ujtz5XX02FROUFi/d5k71ueXj9MZcS4Cshw+uW60+eicldRCL8nkTOAG
58rvR6juSpCETrcpseA1MV2Hi6sMcqbbpLtZ+KDhm2v2of85aVULWV/4ldrPrtdlrc2qQg0roq/n
59dg28AUmyEDVxroPyhBe1CSmjm/369VGH7lFY9SDTvFhC0/XME9kdA87KBGWzJEGZwQWN6IV+7N
tN5r5jIrGHPDzCmG3tyFaJTpWihEj/AReoH+M6djqgFUT9UZYK4d8wC0Co7F9XQR6zN8W/t0Qx0n
NNXnBF7pv9F80KVCcXbxpl8YTOFjZigmAEjvrVCfz63Fm1ZgM+5UmsJ5hQzIGQiCKrYofw1j3C7S
/zL+mkAG2RCQvnB3W3K0wvYk46aFX5wmrr7kd1EwackGw6TIF69QevqEqK/qumVD2KLsu62NN1Om
GvMjWO80//WVe51x8y73DaKwFX3dBVO2ebX0Jn3g0dToClRpKCyUThJ6Dg9prhTNagfSkgmhiQmE
/Zt+yeGMwOqQFdY/5T1huc2u6IIVixiCPIsRes7uXX2qeWzsi3ScqT34H4QuORm/PEXPUF9+P5nQ
sjp4xdx5K+lBzVTLIw1HzQtF5dgdkDxOEjrezradIV4Y9N05kRUdI5Ha5fLPsbH/kvF/IyNEBxyM
9XHPGK21LUaEpReeY+r9EEHc8KUZxokjh2rqp/GHshai6hRedaSAAKiY0tq5uUBDKObLMBLQtCRf
0rIvVgkpwMVabQB6H4Y1i5RwaZaU6QWnxxiS+m2kUOsds3Z3dAL4O4jdkPbdTf86bwkoz8uV+csx
DwWsKsKJE6NRikGkHjzE7NgIgPe143B1H9NyzP4f4zJy7m/XkZhWmzsgw45RPURTRlFdDr7XLJjs
WtbRzZe0EvoUNN0oHYJbRtB5jBjiDGGQh2r6bcZ/RcIUeUveXSnTQZh/0lAr8CVYxAeI9BMLK9uS
Zbtc+XeyXI/IXoOueUg7qFfcH3N6vD62j0uKzwPdfjvofKGO4XvjjNEEfgHXt40vV0eKdRBwRlCe
xvaXwJDeMA7tKnsB/6QgMLd4tXphjJniOnHKExQkLmZTRgrt8du0efktE/IJTpI0caYOqV7gocKR
UWWTkvjtMSGqCu1EHBa9hKeQOVg4cTPjvFCeNCyERngGreBLHhQA6KLXg5vXHm7hYa4Qy1xBEza/
rWhArPI9KzSMe7IPr9BElj9RU7TvKGwncfWVYbAIlQ5u/zwgqIwpb3Z9O1AN7ZLYczHYkGjwYjpB
po52FYR/fDMAqO311l17mVM75mxq+T+cT2HKNoszn9/Pwkwsswp3oMbJuqZ4uxOYalBby7m9Q3cT
yYxXz6wJW+lmPktRJky8AFrLLGQwmOagPYYuMbYNSbqMFexntgtJDGUqnrt4Kgb+HSdZezsyhq3r
g9bggwfnP5Oxq5xQP3KLv2bFuJ80ke/YmxXEm/UiYrjR6aX1MxkGRs9ohAPysq02IIZ5zhu+WwdU
q1Yv4kds5zcXnKQ7y93VBr0a/mJPL7xB9eQZ5WV2j5L/+QDHGnnzEI0gI1VOqoHVE32Nu8Zz6Hnq
3FNY7c+exu5//ATZFdgK78x7Vc1ti4IA46KV8n9gAsAAyUOgjcK/IxQX0I0j7aGcqFq8LPVSkMT/
SG/inUqy3F/xcslJVnhBnsxGzSxTlgq+n0yTUqWvaZpZhhNGCxfLk5vRBnkaQozjUeOSgysK+ra9
B7UfxnWocrf3H2x5IDn8es2rRqmzqbTpYY1VahN/hchriSPF0+wMnJBjB7+G2eSCHr9vJCZvh9V8
ED8MxR7cLScQf8mkoJ0W6LDORFxgUfg1LHSZJ2d5vHq0lxS2pUqmhmpLitYqoPggWCm0XO/UQ/UB
WKCvImYgYH/zHV7iaiB/8v3stNddDdLfjfkt4fhXHebhe94MbmxnLymLyGxwuWh1Vv78hFxvwCkK
3zop9W1K4im6bHKiYHeHStkeMi2atW4m4BZXhlPU4h2OY2aL36pCDnQJxUpvFnoUEpi3pdnbr2Co
lYyrkK/CqMEffLnkwAbRm4WTlCk5LbciKpopc7irOVBKRrtrk8Z71fQ49Yl1YYF206A1saZ+ppYU
slb7S9jHLxHOgEevpmIzT3EszXqnsZeYQmu7IDUqPzUavuiBK5YmtI18aDj+b1qUHnQPwoNa0yoA
zcnOEtWF3bfFkbyvBa2yzHXGZgs63VJaoZXmnS+0CGyrOCpIjynmKj3t+XwrU5SOxvUdlR0C1ZaJ
wRmaG1HgRq6bP1kseVjMy8S3oKeLRpuIa1bZ2Ev8p8TkIT5ifhY2nKf/VSTIokV+fOCiobNQjSLX
Wm1/TMfXwBWHJ3OW1KiHyGMESPImCJvZlT8Z+pi6/ys4+FfbQRDHTn620u832O/VvjAEoPBTUzVY
Urp0yzJlIoA5fExX/6ESaBdkShfUJq6SsRcQBtscLm5GzvnLaTfudcbZqBKeBekv89XzmZhi/wck
2jF6WkYkAHRA5eQeofjbX7bHaxGiaZLZwaKnkt13wnavlcn5Zso657r+eZxceDxvIDv1Sd5R1AKc
Ky2cYXO1u1Gp+gPwlb6cpb9Qp0GDUN5ulbQr0TUEm3wJp1FKfz6DsQnNNQShR7/Qf0iVdig57gkn
BW9t6unMoWjm6nROXozlMzUlNkvb6VAzlAv79vhdZxnTNqhps75PT8R0xgRhJHI3KoVriuQ9/wxE
GZA31GpZ4uMccoTqHCjxqStcEY/fbfTYqelmLHm0Ao5geVNfvL+jKOY1LoVsKVZyui8i4yEcehja
aeCxn/fuOJgL9SZS/x8Wz0m6FsOCRO9FrNe26WPpL4itJ+OyRPsjWa5j87DwAsF99KgUEeStTJKL
Ha3BuK35wPtGGZMkK2Mgciiqjxc0L9UTD5y54Sf+yZSOFfD56xz3J3tk2gJjuzmjGLGypcPD0CH6
f+bIL+TstYQHf6HBmZIgFRzssXksSeqOLXST5/a+aVVzPbURIkeuxzJtPaz3KNDj1RtD1hmRsaXJ
U7b9Bxi6NPqSLrXACxiz3OQRfJKj6+G+ue/GFvoVhJlULt6PPYh/iUM2UlS3pPWFp8JPEKPdbXh3
tEoIotqbCqYwTMJEzgA0sBc4Y5FV+ENi2ttIPBLY+r7XECf6nd+JuDHjO7f/oXMXfbeEHLxrK8jL
xupWagKzdPdk73pC3z41W9eD8xFoYRuZYk8FvWUnylEh89bIY2z9wrqHwHcjQHDJGgglsrxrZ1UV
3rbkBtJmp/SDCjcTBP+gR+KU5lygQYLU1HTRPXsDfM8mNV7G4Tc9bfy5hJBSDNj8nTteWaMsfd6W
IhYIWhxf0sGQTUmRi8f/rJnkZX58Y0FsVxtPrmRTvQX7P8H2yM9FKuH+/coqB5IUZfA4X+h7XLby
PNadO4PD+w31xY3vUHKA5C4ZyyaBkSOtVhEUEQsYmsozdf/JneQnKRXZkl7Xu0U5sS019Cpqo2Lb
ZU8G7xPchF5b5Lfh+jJoRpicamnQDY6lD6vidf9Y2EZjazqwp3Jc4DBcAQAcIhvFesZgMJvBARkv
/9dzLtsktPXT5s8Y3o2MrFYCWGSi51ujxUpsUbl3xlFKJD6a9f5mYfTt/iPYu6MjNzj/pjSlxuA6
7tSz7EItWp3HRfFQkTR+mYyMxOgjJoOt/TS8JY76jQS3SEbBj0AmL60ce1EQD8QAaTnlf+Kmrk6Q
1/3sG0/beZZ0TSFn6K61zZKIt79CXLybszGLYobbvsaVpkZtXVPMF9d03wlyKpWHJ05mbZf7m3wh
nsIX0AjX4NzLWyTAr2Ntyi1ZRVCDb6i6QSpKduahA1gj3xT1J3pDsr/NO+MoXfZhRlElAwBOG2/3
sm6pJfvAOS7cPhHc2pGUdIjMaLjt5bdVnsQFQ17dSkAMANEdkWwjKOTKKm/UGcMUNx7obGq5Uokc
YSi2l4RWvbsHReKowqbujlVtaWDbDVNAkYby0fUenJLa2LjbePwwB9QmCTtDEEfbF+hpvXTT8DEO
yGeGgsc75sJc7N8WlXLh5C8nuHeQEuvpzru4mMDH5qHQTYsb//c/i63m+Xp9FE1jaqPIsElYq2Uy
G2KZ4urvv9Gmu397zLu2hmS28BcQ6vo+L0Nmba0TAD/WWr6SLWQknqTN2Wxn1URwxuvNQxtQqnUq
eRCtxT3FoioP6Z5Af7avABgFJ8pi/PFnLu4DslyLTEaPqjBBXlSYnhcJ9CFCyhuXM7e0NQeTt8+u
SGd1IBV+BhNXRUHa+ZrEsm1xzlsOjcNMRmZsov5rVFjOutyShPamuhWzdc/5Y8Dg1nNAdWkopcqq
9Jn5HhvJBntNNeNHndaanQFJFizol9lKW0KLXXCyDhRD4IZjxLdF/UYPlhvZ2hxnpyw/JiqsAEi8
daaRjExLUXD8Jva3R5DW3bokMe4TJolOa5BG0PH+YSTuaOoLHewBVo18GPLJS/zmTOjimS9779Qf
cxlbr1QGVbwNZB+A07IGYe0NX4jTya6V7evxdOEfA0tB7LO8edhZPeQwyhD4EP672gXhIf507wig
6qjmG+GyM15XhT+klrSC64bwqvLAU8rlfbqa1+6kVCDLAlNUTGitwFIJ4kY4OcrAVTELYtka7t8U
0u+BTN17hEuL1YkSZEgEtYj+k3oNPW8Z2CWKQP0tqK85Q+tOGTd3kdw5Xn/rTzescHrfpiZ/C145
J5kS38RVGrOb5ehyTAR9rRVrbjEvry8Ku2gCaYeRNtgahI8HOBQMRqnG948nzgZgoidW5fz+w3tZ
cAsLu6unzyEw5bpR+bXubQtS5mh/6BkWsJu09DttC8KI4aNhR4WpqIU2bRClS1y9wACbFWG7M+qF
+3rJT9bKVP1X2rGELzDmYh/u7Y6xmDUzfWQUEpUHnyjqv9pVja2VdBxFRxbSLAbWEn6+XDOPlYvO
hMj3uu4vo08CeLb292OyF6gWHLjV/Cu1EhYqB5FLomwHWa1q2gd+uW4xs0Bsd6skCpC7DB4nzS3B
R6CIZUbKNPyWPrkUhzqSSp9l7XRz2DxgfDe7XwAjqsDwes07PAWdC40BbAqh3NGkuzV6A5VMJYM+
RwI9AQVufG4azjdFmKaD86WnTewiC/mc01X5SwC6Y33o1fC085kRLqkSciD0mooQ2+DsEMR021mr
GxOa/JYoOEapxZlekpJ9Y0kBkzXZFQ0fjzpwrLAUUFyPyqd+to4T9AAfGBOtyX1hjYlxXTq8eU/D
s82nRllWYOVthZcsxmmJ2KdeMEw7Jgsb7HbTHbbQN2xeCQG7GcQIn3u8t8CUT4euu2UaplxK/Msr
9RGh/LAahI1oWeLorBxCIgUxvtzEnD8F7mjvsFQiRezLz/+Sfe6eJDySEtS4Bb4e2FK/0a2JRYMf
+Nu2h6AWw6HArRruLj1M5g2ptegiGirAY7CzS2xTyUFpV5QyVLrO3ywRxnJb0RvY1HfDCs6PMNoP
Em+1RlTjDVmBMBDygnkQZFGgb27fQiuw3A6uXVxINHXqUyxmTTGg0ObPmwXLBL1LV3qTw4div5xh
khq++2sHTMAa71qxnhR7ZTUaLjLTbMsD71Sttpk7H/ZZdO/m5L5zjSZNGpukCZhJ38Y70qjI+yV9
VivDtJAQr0Io0R1QO/vzdsuSA1RG2dlljMNnRPapSvsx9yquri3VwSrk0vrHO2MYV9Cvr+bX1Gfr
tOo1kx21ShtCY8xBX41/CliLRV2W59COkQGvO81WM0cF/f07Cf3oGUx2KIPwYXFD5R7/46UJJRz2
0feaSNF8MGGV8KmlkxIvesM6LLasjrFR/bwDoBmLim0j2J7PobhsHfXXLt68GRZl1noLmiGfI1UJ
QUczJpWHau+WlrxX0rZP7xmZBh016r8I9NvYvqIDSUrFNpKupPVLZkF7d1ZHEu0gZ0Q8mt1S3ONf
q7fHcAtfHkpm5AvatBk1mB7bnUFfIyBcH0gDQszsTvFkCyWuCpQ8tkZmRYnS4Dd2Th1YNPvkbSng
Thw1asrs+eMF8ubQ59omwNdhtj3WWlp816P6z6cnBtvIcVwO7YVFvz7H98Akqc5IE0TwP6m8N3QU
ypPuHovSpj2X6i2pySmi+mZEDucJZSN2xB35YRxKQb1ibunD2jxJ91enJ2dzvmoUg1fdlVUg4ozl
TNLtMmXyJYTvYSfNpnK5f0t0fZ2f49WzwkrqK8gSd1bAbmKevTwZHSJ/cQ8veqKZCs7afzHtgjJK
e74LW+9kCsF5+3+EPf4QXLo28NydTJFlL/XQdF+OVyTTvAOsvSOVhGaoonoK6IP79gDH+PTanMiO
DgTWz5jGfpGJJF9jjBY5w1xV61yBR+3aHPENBYhuNl1H1FGCgLO+KV7iiJ0rmE7Me/YB8KA4Z4cg
a9xrvhMvGPauoSvmC6p148sSQBQoRklbIH9rm6E3p7JtbN1v7HnTVYXHY1HZhHMSNuUqu8tOGFTu
S0uictKt5+bsTwXJaPjgzRuR62Pm6L+RCEqYPIf/HpVHiKOxuAVk5evsw2qmIrIValwIEofBDmKn
cb6UpiBNGoCR+Lbz+hIzBDXJPjfGBWxgn8OrQ7L4mv9tCEEGR+9/FnVhT1rsshaExZtV9cokcqXO
WNRVV0jvXiw/wAYUhaQrtggWk2Q0SjHDomTbJ2X5Wa0k010+gMLSxH5433mN5/yQdODh1T2MWlhB
txWjY+BLvS/+SbCjV3TYhOrQow8rzpNIwL3Gu2516LreT7e8SIl8ha6DfbWbhNiX6n3YfTqUTEzm
xdZxc0qi7e2cytBvfkQ4cl3iuhnzqLwryfP6AyqzdHZWUqBXb6wiU7EmVp4RUTDrj7sHD6G2O4H2
NUgJRbkVi5qj4Z8FG/h+wyo0rzUymQZM3PtqVFSaO7T9pSycX/Tlwv5S4DmYbAdOSM1Bux4TtaeG
wZd0mZjW4oHIgImBwm9Mf8zA+NL2m4l6gJBKXHixaFfJdyxBe7kps6U6QVcYHb/AJTcjQrHmCdnM
mL3+rmckqAs6/t2rrATx7LO9nfXSgMR+Ai8jTAQDacUIExdl0VKZZUUombLTQ+xrh3k8Njkc+2aA
OnmR5IJZMAKAszPVlnsEeXMP8rXrRg6PZ2JjaypW49X5igRm9zLfo5W7FabOC/IiI/9srreSZNhM
DeWuYYLKt7jaugMrUwx1aofOqs51W0zYEqXF0ke/n6V0ufjyq9rgPrK1XsQPgBiFl16AXQFeKYTj
beYUkcQfVBfSfK0LgEvGugXl/JPYdMxGEi/zte0NwdytMf8lhxOwP17ZovcY/wB0Tc4sm5SG6m68
XGE9OlQIkELdQ5ZS+xMDQ5tH0yC/2AFFj6yNyvpmovxRjEOKwbl9zCv2skn6JBGazfei8iXPqYgN
8uwMr9wToqsICeGn6RWbwbsbn5y95Isyo2Icb39OfIGS+7FNYmfnzif3opo29eevnmPOUmubX6Dx
HJTxciPiWjieDfZpnlQfqBTaQyS5CGFqFJrP6KAOfIRwxxc5ZmlK9AwNbHzcAbqlUs3MEmG5/0Pu
T56c4Ttu4zgqqT3jJdlj/eWNGn2DZwJta8GuAOf+NHY5lboaSYmlquuctaH/3Yh0NnPj6QsivQKd
bfExwkSdVz8eM6mpdEumLukb/CwrdBeoa2SYEkZTlt3exxFXNUbqZr2/7AN45gN62wqJKVMv8zzC
Q3ca6j5EuAWSKoMC6tf6+3QE7NN2EHR6c8IZC53qRmpnDqyJOsf6mHl+sv768iDjBmO17WsCIsbj
lGQFvEj08PCIg7/S7PJQp/OWT7VkY9PGfIZ4uHoAAK1erhAdlHWgXaVO0JmH0hdy9npbzmJxaMl5
4FgnmnIhU9BLAZdeIe5ZpCiEYUH/B214fMjCA5xa+0BMKJmQvvIwZvGz4aRZ67wL6x32R4oK+kI0
wegQI9eCJjAh0DqeNNYltXvL4BhgWQhoOv1+XPwSxvpsb4FIeIDk6rsLAzxQp/diazIb5SPaJj31
ku2gbMEEmr3efUtxCA8ULiR6n4oVerWyLEgeVnNCyBx6IaNurjwpKVPMtLhw0QQmzr/tUqlD5KE/
ldEvcr3f26yak9A0xXQb/e7Mmr5Q111PNjzzT4bkFVOqF7+KD/9zCIAWKLo4aBI2RytDNuKv58GA
Zm+wIVGFL7Biy3EJUiiUBlUIon9wP7i9HEngpSNAgGKYotDiDC/CbuC/m3wIyzyDrW9O70lkgCHP
EvGtMf6BhQ+GjeMukuCfId1j7SNX/I4dtSwBKL+4qJg2KrKbTSvOigoAtKn4R8oYzDpacb4qSaqF
qWR7LqrFxlADckxr2RrPnwzn9W3g5kvPxcCcjSqAF6FDHhHwyUh3mU0XH1XxoXmRddoz0k4PC9Lh
/Oj1/Rc1DUwuIDY4C6NJahtmdOjmA+t4JvukAqGvhHPxqXKjIHVeMiY9mstV8MeP6cYuKDPd5dzi
ZUSW2bGX+CO09PrTf/mg/uDXOziCxKJINNmbBr6EjNFPUxxlsFClKvMI8jCSMhgdHP8LI8uTFB50
2Ak966agwJtqObb5pgbcYjFrrugiIaGVrsL1QRGdEvq+tj/E4BVB1iiQD0SXE7SzvM0WrWHa1Ew0
sRBW9xh2EKUYZftO0WPRBy4+FSjBavr8TJWIUBEjllhSw7PNcyY0A/cvvuiEDvkIAoA3GrhX7dhl
PiAk/Li1qDrx5TRbnTSMW1JHD/ZPzs3wBCXLzWRTX9vIhV611FXg3oDJgVvlAjTZzA9YswrdaQo7
pVohl8GDCsU221f2gXHdLpCURasGY/FOFf5D/+vmDAo2WsQ5Z0vB92mehEgiUxS2oer+L6kL0Fah
BF7OW3rgdzxxXk0Yfb23i5EAqgi6agpcdG+y6t1Rd/RTu23mOIFCsFZOxQIHPznU/HRSnO8FZVS3
ksrSh/LwQJy6CC8euB0UPE0OstgdgL0UeaY/aPYzcR+uj3FJuMXcVKY4dm5/3w8uoIxsA8x8/Sdr
U2jZ2kjDIxemzPVhtiRLu14qH778/HmAErPHSi74CnLZKgy8Gob8LQltcSoOkpCkhjI4CdvafZJW
6B8zjgnRBskdkfmcPOpUwpDhjnrKCE8OgjM56HZ3H+GsLvmCmT5UJ188faeKvB1Gf8lF0xd5UHVg
LEkIRpXZm4PJZFsZ6FbbJFsoJDk/sJWxRgWsQHh2usJm5qFLo789P9zTkSAfJpdi6otTrzA5e4ra
oT3IMjcDCzWLqRcF5cs7zNUsqAIyKXheO5SN05o1XfSsSnIy9HnVC+sKz37i6jpRcrG/tPRMS7tI
r5gJxvTeT8KtsqAH+wbCQ99w0R43E9uQ69VKh5Q+uzKBsal1aKznEtdjq9gM2fg4pXiU6lO15AfI
Nm6JT0F6mqaFkD0VrpmkBCY4rlXPQtDXS7RbQjV/43SeoW6kqddDzzHH28fckSHavKMsEu61NVjs
K0heQmFYNynWoDF+5R7opysJSGYF6+bRSLIOKfwFVx0ySI/VLctbmHEmIORs7JlZqzfMdAla3NhW
UL+D4rUvftfQit7tQ0k656DTfeFL9DSPiPjBEtX7Q8WSWvHnmweKVmI1Fw2V6MB0jjeM2yhxPZuo
gkvaZ0fLonke0Z1ENiEB17QA35aviLz9D68SDgagt+OqhGIVBz5UMrLGNFOWXm50WBWr/cv3xk+y
MDkOe2czzGHsghOz4wvWSZ+e8ChHe3DtnhB6U5eJKaIPXGJIabiMrX1kr0Oy9Bwy3ni8tkkx5cKe
DmLAwcHtMPSZq9uXRmYw9IM0JxG4z6VhaIcy+hqGOVWGSPM5A/5ejA5gYPP3wwaY3/eBzlF0NcOg
q/2TQVuFs5oqLN2qN4Vnam0CcK9cOTd6bOJzyQoItR6XFd23yXcacxEjfDX1+diM+4mNZMDY3hUb
+PZy0BhYmZKUKY6885X9MsjUIwu2XGEyQgu5puzHCj1JQHZl6ORaSifDyR3V+yIJZNnm+fQdb8sm
1Z27w2ejdT2Ee/w6N3JAJLIHxTVuElpAwFpmfe0LuVQzAkZobdK8y4G944983KLL2TsnG5LpGyHQ
rSnu1kv+d0JBP6iB38CKgdQ6yk98wlcYO+G6Kf0tpKKeqB2EdMgKrPBJ4+6ZvM/MOc6/bq1PMV4A
d3T5o2LeB5NRg1Oi16+vBTuXv3T58V1vTlWiTI0zhJMNfgVZ1cnqExop5i5sldS8Qww2h8PmWoMx
k0ScRLJQsg7gU0U9+LdjWl60xCyL6Vz6BrNIec3nsNaHEfXO5TagMfEJvDA1bLmLnvSwUlb4OvKl
npz6AY+vv0FvyIYcQhr5+1gLxZ3bMeekYtpF9hlXcGImElXbnjQ32/T4s+wwLkOVgcbCHiIqhoU7
rF1N8uCz+BEe98iL1aNfbwsyhBXc10MfEPCj/bTv0/n2Qfc1AHdLa1/aDCcveE3QZZanAUprxI5A
7vwTx5ghgAzKtTdPv2LQRsOVEkfIV23dILBh6W2+o11Di5TgI36/+RNzLWjtqGDPJg1qssWzEAxg
UC+9mywZqzGsFgY5TmNMFXDkuO4da0YSlaFcCIDYp+RXWCuA/FuQ+Q+f3KwZOIpL0qzqv72+T1vM
ahP3xRwcluVQgRFgLV8OIwWUtc49VRgNPnz4khr8p8hulxcr1V7V4e5e4lJWS5Um8GUrPpijGutU
03payuWDTvOWpGGwmnbRGK5hbvA9rP05L3wNlD1f/ckpNDBiD290q0r4gK2hELWXPcdbqHsHOLXK
Fluf1GgFxdUqbcT8H0hz32u0c1ahqevSgT8mBJb4mlSoLqRrkU2IN4yIXp2iiXbFg3aE6Gk0xLgb
waVhU/x/2pAUTivWDhjuaxEpiEyPyW2YpIYtE58B+9W0IPQLG4pfVX9J7bFeYnzErKF4VaXvRcja
KzJkJAsHjW8QTl9SKDuLtLmU8GCQIur//nFg4stedSiQyUcab1WcFtUTkhAtmX9TOqxgY9s1huJh
xEPcg/x6KSRCGFibic3/RDBPBD1zTcM6NygVgxBI6Lx3CT9ZVgZCuf8W49GkAHb9DOg2qLH+DKuh
zj6YHSafpon9N1SZ7w/MRL7EqBCxg4E3DZLmiV9BQZj+nvdaEA9n2b7QLCmQZ9PYbo12Av6UMoCD
BlZUxk8w7BGlR3Rw4bLxgG2ptM2TWUvNi0Wz2r0z3aIyJysOSgGtWCso9LJR1jEpiv/7QpTEjhNc
lSwqia3nBcnTcHGmD9Zzead78clP+nURjGVPluT0yCJh8l1DiKRSHuIpGsDUrV5Ht7lHa2GSSsIx
jcjSTgdhRwRQYmj9JRsUkrsBvBDjjg+XlAqymP74ViHE5a/mL5YKW230frv+c3IVX7Y4CM65TzCx
jqOi7MXE6ihugZn88lzNS0k/PGplDAc5uq1lz8ts/Yb2C6yDl2NUTJ3jsUV2LPKOMs/2/wXtbGE6
SxXF8yzDko+eYz8vTqNm/c8DqkzxvcezUY+7ryHezCyv9p1GMR6DCyBLpjPK5g4k6fY33G6SeA8d
fk+jGW3p/PZP0QkZuscUViZxJuhbTrihi+SHJzXVwpiAJ6DXS9MxCl8/rL7V/z/YrrgO/16UOeJs
DAXElXqJAH+oYEGTf6ZKnU+EESsrZ/cuatED89F4obAfZL282fzdL2hb0dHGRer1Nedc5yaLitsh
yLUz+XhZyCwdNgVofuSjuc8+54DlWkZpbJtgmoIj6Hd7daCo8q1RWzzDqLQtjc6J/LXzJ+81hJDt
0joMNmRDRs1XtQp7JROo9ceu+cQKUB4+QtxqbHYkVBJn2pchjV/fEGZhG8y9EKy0i5Cjepvxo/If
WxSfNGP0GC+J8uVcb3WH78lGyJpuLe7QpnW52iXROf4Ok91sXCiYgGmRxVEJpUqWTp+smpwZsfxk
crxhcUqpkW4GXiYPq9r6wDwV5irZdZmT76cIS0JV2g9NftuzFo79zPthyprH1HGbT6axKPxyePy6
QkySYZDE2icrxHM+at/TUcRy6vHRoUU8700PefP8NO2xhust5KIPIyYcoxV/tHshEKIdnjAIe8ec
pKKeFioQu9PPvLAyCg2hWweTpLrzkza5Ts+XHwqcVQjPg3J82Nh6q2ii7z2La03X0ags8ritnxgR
5YHiPydFeZRw9XHYuCyqGudpmxxQVg6omfNi1Zq8nXovbeAR7khfVuF85zDoFTqplWmctI7a1aG/
9ny2JuXCa5sdMHA2v58yjZz2Ti3bpyeNUstwbi2tNr/Z0P7wCxOMOAT6WLL3oXLTabrRs4JBA3KL
worXCDHzymqEM11Fjt2eNW0OTnil/cjhdpgZfKqKVGhPUElgVyU0oUgDTH47+HPSlxEVfyB/1P99
NBFryqQ4s2xJ4JiHABhpAw3TT6A5LpFqcObN77OOE9VOAGd+JPCA7/H/TCmFn2HkEfVmibvareQV
XCi5TgHXNI2gK3PukRyyyriUe1RqmOnJCbJWfALHZXhufUqPRItVHMSVhZc+fmhS9fg6oIKCXTBE
LsDUs7oMJkNy1Q8juKHUNNWjSkzYXf/SbY6dVbbrhfg+3li4kdiVztQmhtq+KRmEauf8hFUcsCE2
vqZXGSibXKhN0ZM0+T7FLhYQUrlG1u18ITktOd3fGcuSw/DKR5DJ5EJMPsWhGGMY/J2SWILRIwG9
dBVSi2ipQ5xJ2f/WuHtBo8bWnkiscNEP4d/qqt87FkyM5zH3DBtHqQKpJnFq4T9bvMQ/WoDsr83d
sDYngq79/0DP1OFqNCg/nTK/P6/l/qV18+OUuS+8qa6vKJ/mwpQVoZ48gy67lustrzuaw9vJ6BCV
NiydFw/vWXPQm5ZoQQhNpYnJ2FCLsRmWdpQfrfUjQTbhuzkERTKngLPjPqeR7GpcY8HnllYnqt1Z
zEYR7haMB4fNj3zcUkhUel3m9H66J6VV9KkJHLKgFlY4zkk3EacJq6AYt4jNU4bSeNbnKDCqlbh7
UOMDkF/efVV26EtsoEwT9G6ckLQ4MvAcdNjdsPXY7QIQpHlS4QCAorfiZGlBxBxlzowGrC6Qn7ph
LZsyFvExV9ZDCfUOkDJYkj8PqWrLgPLNM0M4y9iMvJ4SLMwgWV002hmLAswL8E9tA8ncpR4b+gyt
HHPRN9bm+NS6Gd+uLjkbfV31pKwTo011gPHaSdljc4alzLfhFSrLI/o098HzQVxFAP7nkb6ri5U7
MsK1uUjRcNZZMoZ4gfyqVAkWS3F/9sEwFFi+qxFy7ArFBftXt/fVJDGtp/sG9oBa4j9brqGISMRZ
6yOzxP07AaNR67kzZAna+JSlMQuhmB9ohwEVcgv0tr5JImmMLPGzibzXcZvLjjPKdgFyGL/UmJtc
7h/e6HBSHEfH4WwHaT/2ezUsjqRqQsQHNNE2xJWTOiUZu/a9slv6tQ3wYTHlqa7fS5Qlf4hNbQTT
JyFSMfXfnhAIwgn1ed48I5euV2Z8km8+o9cenxv+YgL8KF7gM4lgAzTjxQKWnJwWpznHD1MS2nc1
mA2z5JfpNGGdvpgQy4RCgAkAHByI9i7FjeiWlNKBuHmVFdcwliYZF+jdZtJQPZghEy8NuntD0aCI
WBrsk62Fs3rZdoalZ8DlkVRhc8+pgeXqhr5NOM+B5cLYArBVz18v6mzGtExQFVoXiv+PJwqu0vWG
3ggok6MvHFsfORRYzvv2MgPB52KxlJfpmz8cCbelerI0kA5J+5mXSP5DmD6bGxRH+kR2LXzbLE8R
ho/KBuSKPxTL+2yLO1yqHfnh+MwPdRqdVuYgYa1WW3nzwye8t8jyo84gl2d0t220gbkI2IU2VN0T
h8ulXIyrGDkHhEFkBbOkBHhgFa/Kw3ahuWdcSAnydLegBdggg/LKVX9CWohlDxO9xjpBcr6otwy3
iEAGX6BemdP49eu+kfJm32afegU05guNWB5dvrdnVMQXLuUJwNrHwe0iHk/+00/+vRaVNEAiaaTY
mayJabPxM+ESm+gNIa+yVS93If2cviREUzD0jTG4TKYSDjgSkzg490QmaENccB5UCSPf6tox7qJn
MXzaMxA1rGdeQLho2p2DkBaONhy1/2x2CkHylQRZEhEMAkBr1sCw9eG1iHD/wKr6u+jubF4QINZu
r2E24n+uazeY/5etmatq4TEwinRIoOK3U4CnhD62Jnccfi1CCF5fjDzUWKIc3xRVN41fzIyQnPMa
6Q+tToY605GnBU3nXER5hx1FRzrxvp0F3S9+6KLvlmGGaB/h7uB1uu+4xGKMb0Yhp9JFFGGXrPhx
wLPRhJB/Qq8+I9Wq/nxn36qoKmO0ezp73OeqV++dC5CwN32ezxd4kNwHsG/6aC1B1yeD/bvBYNT5
mTPJPGjVtBWCmU0gwkZ38nBuvcRQmrHO/FzVr3Xda22t5iQ35NXGlVdAIlLczFNrciUqHCDdOb37
hGaPJPTonPT2e6kXFCAumsLKQxNV6kQsea976Hxnsvw4p417TMQ07xAexUaAI1mjHVL6Wd8RpLyv
U4KJEpGdGbPFBn2OkObMtK9MPeNGtMaSlujXqgeINoL1Fg7/xIq3NpKYQq9S/0rPgGufFhc2wMTi
dsaMtbs3sSNnG8umpTuHKNrnFioVTeO1aF3dHS3BgIQkvPRdScwZcTwl468hV6wB0QkLSwJ/MlXd
E2SwclrtAvfq5qKAuZ7juwZOsJbX3VjddHkqTLuy0QyC9bfH/xInvqS9achOrkK2bRZYTwtY/J+e
5qgAIi1ERk4ksYF0tEOhbFldqHPKKpVL+nzLPOrauk4BNle6c5IHvBqd9SVmaDpoHGa5JOUsucPV
kSYhjbr7jvwYjJaEOvkoBiWx2r3j4zOz3eRAInKrBhtkLDRVnL+ZUlz61Y5+De8/8hXP9kSur6YI
/dwWFgBGt+XSz3OgQp8/bKZgneGj6qb/rQ7u20ZFsCdhR5C/CZz7Uh5PEHDTbXLXrxV96pK2K10u
DcfMq4BgJlfiA1i7sdzj9ArR9z2ALQNRGInLrqCQ57MqWnfqU490fq1yCqIB0N9Y4uvs0eXRy57j
b16sF/V+J2xIsfnrYBV06WIhL9vF95+PHCmqttVv17E67+cQ8W66KBCJrH4eVfMyigj8trthqqHA
XYVP99rG5xSPHU1dKNOj+nrb1Wtwp+srsO0axu1P/XgtFUSpLkZ1vLDb8a1KwkyPqXUruZHCsxtZ
IPVrX6KOmXAHSSjAbeQGcOV2h6W/RXjArQJVuT9U6xKM9DIDDvQ87Wfl9DhgCIC3W7tvrUh+mVjP
vc2/Ip4i/EypcBfsZc9OrAqotmTuk0aJf1med0FKHRBxWRsrdOm85ef43mhSOyMzzGXyLO9yA0FD
RBmvcSUOrbpqruPqA2uhV46JRQ+PlZxPyoI4XfU9O4/YvaL+gs6+NdZAcu9HuSwhyIToIUPNz46i
mk+75fcvXQG2LCCb9KQVzcGV29mGKfQE76UpEqnbrXDN4KC4KbxG4cl1/F6N3cDPX+6cKIlLsPRF
OAzuij3c266tlSxcfLyMEn0VuGes1yEyViBam3Zm+cI9iUlJdkU+oEeBS+CbO/ffMBVxiXPS/LIV
aZN51ZtYd9k8jd/ERJgGn1KJCYVJHMlrhhEi6y/PNx4wbF9HN/HvlXMx01aEZVhSdNADquknKmLk
nxOYiFjhxToaE1Oes7vmBOYaYykH1lx6zSCr42oEqMxoX3sl2mBVE+SYQI5OEXVtXhP/AFN3C7QJ
16SOPDdX9W2tH7GTTKX4V01bzBqzBZ9KGqg3NPt52OMzAi8UF3scHeFKwmXsyGvus+QqClSfuddR
exvx4spg140CHhNlRtK47wWOqcuaffGDEhDauN4Kh6fGMfvU2Xiwj9sQOD5q3y3xKdXvvgrZhjis
IyvP4BQEFLC9JbV4eLA0gzs75Qgpk7nalM4ogFkeT50qE2Xvios5CYAkZfvCU4vIh2wgc2KTIyLm
carQGyLCNhHE6K7N1IChAO5sWIfV7LhjBD5m/dJn/h1vnexA+jswrPe4Loxzlz4HwF2T1pfSOV+6
/SbdZLs1ykpz609VsnL0SRU7EGjSoYoRRl69b00DsvlxOIjB919ssjAFmAQHY/JOU/HYilSbw2gu
KRa+Z61GS+RV8/XoAPxiTS0HbuPgFajZEYHxJuSjN52IUM1zW9lP7oiaJdiIQddHRkZ9r2oOyrFL
sHVyl7x9qEFBnWkK1iNARSNVX+LC3Wx/kTgwzt0jiVIlU1gbeSEmE75snD1y2BlZczMiuo/3dFUg
5/zJSkLZWp8vtDnJ+6OZM+xKoEHRTggrzFlUZTWcGKDs4jsH5BrDcBNmwmpNoGaYany49XK4jufD
5FuEnjPK5q0ra+y4uHr60SGaklXLDRLQcLICDfpAYSuJMUCwSGgyVM9YF0EYyUITkdiSi7YTz+8R
qnw7Y6j0bngi7xV04XvgMDVk1Re0itZgf0SbRmX3J9NAwI9YWiLojIpw9q+gyWN58QBJzQZDdYzc
xfJmQ9CTBRLLEpCAPucNsMGMmfZn3BUFT4Ge7I9uwJDD41wjbgQG1+4VXz0kj1xlDT+svrV7p4hf
y/kbI6Ctb4nttKN7lU7NmS15agf7vV02TCX0dcWuSAqXe15B+vnqycP72gJLQWVb1JdCEaCk+d2+
OdmT8ReImvJSmPsp3dRxQIrJuwIPnbJgwicNjDuqdmFizRbGolOhijXT9YBqKMByESmKCei0zeQ3
bCmjHahHIgW1hy/FWOVnhaaYqVTVUWYzI7xDMrHT5woioUYGdBl56VRNnF5N8OrC/dy4ns1pUwXw
+4xfFEjjCsnFc4rBGtbD1sAW8AwWpFKt9wocNVgi5ROKNg7UCkDfYyFZfk/3BlziKAnRxK16tKu3
nPFFJlu8bzyVr2NMeaMCKX6oZKZJko1dfo9emZ7L7x5uce4O5XBXicucS0lN9yDO+LRxFz/fOsgt
kyZ4PDjzE/AzpoS9PRho3iNfMvt0mVCdLsQcgW0DP9mcndAahToQTDSJtrsvTtcZQz82gx+nOrDm
Z/F96cU5TeSb+1HmENU4n6Dj6pRMVZKcGuCUmhJ2kWdE7QWg1GUUWcVHZ7KO5WfnD2Z/fagrrP/k
/NzHsSXyVOfXh/9+HSA/tuwA+8GAvunlbfEkVUbjy8Kh9EoERjqsTwY/yIc5PJJK4hN80y3yvOqK
RfZjcN4UT7HzJ0B2L10GcvEQuCvGlKMSFt2qz0v8XpPKydVBzGSRyQRERlNyd9X88gWYdjyY6xsX
g2cCPvaI5U0nHfrH5VT8XnqJcFNd4ixomFA58EPSfVnazfv8VYX4/fVdbofXzNpy4bmt+McRRpg9
jyGLzxZAXay8TDDlHk1d87HLb8CWzGFBJNSPMDUJZQ6bDomAscnfXeZQAw3vS/YIXv4LXNIHfMdB
hZSk4njbHoZs3bU6yt/e2nc0wuw0Pft3cjupBfOAdR+jkZdk8cyacRiuQDP42y9EnVGZSIj88aoR
T25yll978BML7Vl5tEiskeuxzq1iWuGvWQYJnjZN1vEsgFaP3ganDE9/N1iws7KWfkCypoM0XWkn
bIdT9ytTHzOmgbojtuq9ovqrLvwXBlhLHSXFi9Y+u0650oTg5kjUBe1m8phl5+hKTmes4qCWB9iL
+jtd+27oyupAZ7pCSlN29G+n7ZwpMofV2w1o6YmDX7jfXuKYQJH+RplWmxMqlmNyRAKgkbkpbn3d
gr1ljhY11oNVp8HqvaFYg2BIDRyyboMFPkZfZOZeJ58r7znYbSKmW37SiexOrPGHT8VwaZusJslk
loavPpBSoCjZ1zVJcQ2bKpMcOYaavMJiUs/iBhYV436HDwkWYPyanCctpd+QbGqUNrI9NuvNWZDY
+G+7XC66upm6PkExVMFRTmLeeLYHq+yXhmxDGegVlR9tonEr9s5hWraNuOhgGsYRM1tPX1NdeBZx
yHdjXXdrpKC65K7AS5k/O1cOEw0UT77uOYThr+ibMb4oWuykFpIoVCV9hJt9ETti5NAAJvFx4hqv
Y2rLOPEz6gPxR/LvewIkktpbHFuKTst2CTqDnEXqy6+nYcEQlYFH3DIM6WFP61zC5bX+dEqw2XxT
tWBkcxBBEobh0AuTTUFMrX64DWTH82CMqAgPBtWFltUgWbmGKxedQDIuElw1ezn+EO4noD68+NPQ
h32zc1mihr6rkbeUeID4yYe0UW0JKnq265lM4jEBgoA28ZntS0noUFxNSgd6lbATquxajemc+RR8
E/CaYPirWleFK6CeDZ5F71NTzksFdOfDSNk+7pSyI3oQAzk5Q1TxNgzk1DA/s3MG/XO/A2kXm94B
CMQMKd2RDp6MsDbCQ0sVI81Se1rdc2ZJe2GQYnv5YIlraCyiJNnQZ3GZmRGhMGIbDiWDXGFY9AtB
Dk+NlAi5FxxSTHvN9F3CtsIRB2GiGgCnX76CnBDu1KRDJdQNL/aZUJ1/VYcwgFGVUnxVW481fXWO
IAa96XVsTf4cwmABFL3/uj7FBmegtpvbR8Y21t5QZjgUb4zOZBl1VsAXNSWCLQDEp21OO87nJppL
/IaWJYABmrq2RhrnxDXU638YseiUbCgEwDbVD6WYqY7wLLimJXwF2Qu1ybZCSddEqd9zeFyvXwrG
H+8831+XMLdevp1eRaau4XduR13mb0hkN5FjhZth+d8UOK3NINEBffaFWNZ8l57dKAE4b1jyZn9M
KNNFohUw8RcL5GlvUv+CVUVTCaYMUc4hFKbX9wX7PHN3qNY7ksiD8oOGK14D/tfK0i5pYenL8IuR
sVuBHC85amO9Nn/BEheNTp8uuzj4QGJfkXx7e68KmM0psCr6tGi745PBxxqQ8eaNQu1Wu+j3X/oy
ft1zjDjq6kWBRklHgvJ3hIosHjX1hDBKOxfyj6kk8OQFVjbyK8hMLB4nc8Cpvsdv5vHcONj3gNbb
+LpRRELyAvJRH+3sxedRXLlJIxbr0EgSMITDW93EiUGqH1V04G2Af1VzRSh5woNeCT/RVAqndAHR
m9B8diaqvSKNa0R13YVd1WqlrvKW+ftGJ8jLR/zEg3QkKtN2dBxrqjQplTfQ2Fd6TaFUnpdfylfC
BvldTQ4lg1SgKDC9cdf00PiRmy44SsI0QyFfn1zMOBO6AN0jrXYCKbJpT+QUCTnrb+0tfg/2dB/W
nsG9PbHF/iT6INgYLBGQgXc+GDtUY/qqkKTwNLg8sT0MdE5CzerKC8M10plcZCyaIt26p3N/AM6Z
hFj1pbGNsAsUVbQPebB1j5eBbC2T/+KGsrnVL7CMaHIAbNF6rL+XBqiwzJjPpOX2K/icaHjDvL0P
tUYkTONFxetGGlW8gFYlIQ/pDu4WJNSWFdEgWSUQJv72awg7CMU3MFxF1uawXxLCoBUrYZZF5kfo
nPJN0QnKgFmJeZVuWc6JUYwlpa/2UF8Iw3YuBvDwaH6G34OvrDTcsKkpgHx9Q6O1FK8euauYw53M
BX92H/RaF+DoHE34B66QwrVDpFQ3mXxHq8d/GEBQ1iNHE91aIZZ1LD5UuChJR1DePxX1/3IVSdLZ
nAysxwdwoh/7sZxp7UcTyeOM+dHX/YFtH4rvc8c4e+GbqYNKeyCUgMR4CbLo4XIUmFflr5CHt297
QJfg/eYEfFJnYjAaHGiJWEmjwu0Ic00GD8c9xrHYaqgUVSr6YPLrvE2loZgC0c5Tf9GM+2As8uLb
2r5A5HWSuHYtUc0BNTvT6i3jYMkEHQFnnEtBgpraawimYssBKjDNAlzApCZUmi2G6R8HQVtGEbG2
nGFLTUF5cm4WpyJSVVsY32oua5Eb/+CUGdT+AsLQQC5lyJQYRFpb6GS126ahDgC5/rqL/z9u3voc
knTn4MCSHEV6p8Ht2Xex73GVXfXpuSEoQ8eTLDzj/6eBNS/pb0OS93mshoCyiNBh8MmPAhGu4mJI
AElJoNAXelgqwq8QnHCLzQKvmbORwf/tiPkOKKy9JswwwX2GTUoOD96v30O1N5NCI+EvKKmYPiKe
kHS7ghotN+p2eEFnQgg3GSUR7UzyMUC9vAagMXGY8r5GFcITLNXSNCq+EH/RNSvSqDL5W/BEI+c9
dTi8Ecu9zFsNyrB3gDcRkzh4PgEbDdrBwuztAADeqKLX0HRJyrNGKeGbO7vgGTwWIc/K11wiyfF6
w1PdbFfXPYDUBAOUS2Lvb+RyRbWk/56WOEDBqo3PAK7KoBMV5w3UCMX5DTkM9NKpDdYxRYxqyC1W
OZ/2IALqBWrU87PkX5tBX8nGtURkLcSw9jt+ZOhoYVdAo52IK2DVOkGOgTUGp10ce5K188bDgkAT
9sPojmp+JMXau/R2Iy5jEjHLEzWZHzes2t7pvZwg1Gxq9xRYcC1c2Pj6nYyamPMGIyDS16PT8QcB
5+jj4w6npm5y21KPcJRvUvaAT5VmqR+2/Tv8FlfXMwtrv08Jg78iEnpeAdA15q5ukp33MoIHMLLT
SgPD6XWXusWhAUxhTJcipUdCvTYdediyPicw/+r6yfcNHsz08F3oE/MhOzr9B76pIH9kLc77bmb9
Njzzz8rJCECOXriPnH3CYInE+gvqSPIf9JcW0dbHD95otMn4iXAAXZy5S8q0AWlctephnWDwz8/J
GyyO72ATHEvxWSVl+bwKGH7Lph5ZJV5xV9ChBRu5WNdruLr0r6idCOLv8Xakcqxzc3/ie4zTs+lI
AYU9iCrtHbkNdMAxIUuEvY2FcatVcxaP7lsIpIaKgK9anOw6nJHui0KNCOKFBoE9uRvPYsM4GJ3C
Xrcdw6flcDMkihm3cmmpADax9BgoNAFyFzzlxqHAHD/iiKCE91M9jFw94X+x/ybU9g3K+hXZ4rky
D9pNO3NbN5G30mntO2YdBypLqgDZ4jGUJRxgYKn8Rwrcg4IXtg1ON6JzF3mPVm8F40UN0sotr2eR
kDmNtUn1LQQHDNv7cEVdg5/ly5MHmkWS6o2JJcrfVeqaH+dHRuX6OXYAiLGFG+XJsinKDo5gftqY
mCJGKdaYbcPk4nUTyHl0yIDqKgRQopCHdzjfyfPmPwuyq9JrSdzra3a/DBsLevKhI2o8eWrEzIEM
uhsztIg0VXy+KGI1sCxqbOPqI3A+mWZ1zIzdHdeSxAOHLAPLDdwO5LoVBfEoUlN4dJm++VGjE7Y7
M+DUnpQH5YAEV9skdlilO9EL+B6vDHJK4/OigKeYqNHj/NKQqQBLPGRJpTpWHDvdSMYmNwzJtkpx
YWDxf8LSoH7SeLkmDm++1vXHXuwR6AbQY2544Ev8bTR1+5gJYkE/zBGwO3cYrPMQUOs7fNiontsh
rB+4wZb7sf3ijqKail5pxwC7WA1DJhjKMlggY9cQGJ8qe1ol3pIaEztomcspdEmDKGZ9UhlYelaa
IwIPLNTXNdJarRdPDPrrRHLQd6VaQYhmeU2J9PNyKW3+wJOIrDEgXQeb/DqR8/7PLRTQWXvZStgH
CqVpHsSrg8uh/4fGkTRWLZh71E+Rb3mYAbywKpILSmwkJ/VuQHqHjRLjomNvAQB92vtaWcIuPQhg
e1vIYBb2jQdw1B/JBvE+xItdipJJs84Di7HHV89qvL4zSfeWDgrsKd1GHcQ7Q3spV23UVKz4qIZH
F8fv9YMAeBYvFBOWzoyyI2cr4pyFmQDI8T6I+yiiwD1/M00kZYB7Gi5tBu2q/2SUa3FIQwpAv9SA
secOC66CJNWQ8lofmfmYTjFY8PfDtRt5yDsir9y1cg1pgK2tRrSiz8Nw9rxiGpq5OCHor+FaW1Gs
Sff5zerYP14JxoYv4bdV8fdSPLalHRh/r1P/URYCwi0PiaAb8eMvl8SgkLupvIsjs4u8WeAgVOZo
TnhhBxZFyou8Twa3LG9NG2/HQMOH+MFhC1Bmxq7ZpATP48KoDhT0XyfB6bCtWY+01NDE1BxGtaJ1
SuSvBhpmr/wJZCzCtBg2gQ27KzlpPbI5a4bhqB5JLJHytYqIBOmzJ1wUuZNHchumEPfwoASsCtqR
Ppxwexlz8Je2sAMCBc3Xw9/xu+iekUdvCAgH5HefHPlh22HDJdUnGyA9DBhcrp/X8pWf/awmSHfJ
B0UuIOguNbsLjMNKmFKl3jK7957myOkET8sHyVcjuseH032xvko/yUPnx9Hijk4Q2CeG4wYe/qUY
CJ5Dv2fh16sTWMiDSg5B+BOGmFfMl1MtSuOs5O7nQ/2mVN62WrRCLBM0V8uOpnYU/Mthxf89pcSg
8UslcFUCES+QrcmJENrfZN4qK2Gg3rlbmyMNiTQQDCnytLAPlAaUeQyD05iQqn0faq2vFsfg7g5p
vAd4miMMJ1pd9s0n+0ereu6Y/xxlC9G7veQjeYu+5WhAqcmlZvtnFHbvNKZQ34EibtlxAB3mj8ig
HZje0LMrOhfms3ouvu2v/ZsJr9AJx9mlS1JV2gukh4bQhhDqIaTJXRMwLbbDlKTEzOtitYejHAro
2bI5dH1JBuDCi7E2lyhwqOpj65iP9fXJlbIiKpewniefF0O6DDfKJTkP9Ubz8o2b156Z5fmJh43s
Ik5k7mcROt9BAaVQ34Ksv2qh3ifZmRv3U1PMAPpmjWNCT+BErSZOQlDc4eUsnAbS0LnkGdlNZULH
R8JUbRPxCmC15gjA58dYY9JCU3RCfbBi0rkLJO1hSCpKxnCpvcd9zVvNKNQjPovESoxhzfQ5h+h4
Y7PYuKUcgCStEgfjDuQ8orP6S/n4zIbTeeYx+L+EdwRoC7MDgZmI73TkNdp34kS5BT/wTFjPStvY
+KXpcWcj6PTdC5pfA0ADuCNmIyDHnT9oq+cpJN3mUoAdhsDGIRj7beESajL8qczV24W+fovJ0XpJ
B3J1pVxoNOh835Frt4/SiiCSt/FslM2Krk00sRpK6XtRmp35W9Cz5tZYng3szg3tqfYRxOOK9Mj7
m4A1WKa89MGTkejVFRtIPtcjI+7uwPKAu7TDvufkqoVlYILwthTbAgu+fYVzkA3mIvFrRHXwK7Gq
uugyEvRt0JzEg3djoVSSBGPm4UQKemQY9IqqEI0lv3WraOHWxwuvKhATwJN4631afQYEb1fP3HLC
Vv894EnnQ4jI+J4atsT73O75WIVd1b2bZejaZrm7yT5RoZCGC9XAZGyIIIgozxRYxyWC056fFvOG
uMKGKgkf/QsiLUWRhLiYVlDQCNdgxL0IOHiUG+rE/et+bSdLKiB4hEvOsuqTSIwo+00C2ImCyvY4
BiTY9XNgM7AGJ6hSYGB2keO2w+U1vy/+cJROE+vkMzhDZvVviFWI76PIKC0j7669q7VCU4Ucr2xo
H4BURZGimtK8z4e27Ksdqj1AzjmX/ZApnAdDn5sSmv+jA3rdnmUAO/XYBKvpQrXj/pTzhoBYWXF9
pW+yFG/nzdEVdEgbV2B6vcZUJxB0XNHjLb+lRoMksEpAZ5EntxiUhAOx2NIYQjBf7Mvq326uIrmQ
DXtlyd9gqCbQeqlXH1s6PIaL28LtmZ+i3K/doPKZBGtTSs77aCBRFKQeQTsIrDTyXIj4FmgU58Op
nmtpoW39V7y4uMA8DDOsYKO4yi41e1CP9MA0jpc+FQVZuNRX9xB3MMXgcLS0FG4/7hRVi4IJZkn4
WW7DZfLvNnTsQ96UMh5mUUG0y4YQauNa8xRNofhQ8+KtPJuSXmTD0aJfn4s/3toutVvSnQRWcQCC
9qtq6aPOzQlupwTK9s8m7YbFzcXLzUqQUo2ExX+ZcetO/PnqKKdmVl8TxjA9iPhMF58IZzH7Nryu
8UeCAmxSS1UdJAKyh2B5QuXK6VdUJCd4zH47A6AM/EVSk5j3ZfHtr0CTncpZOZHNGNtlWYmZz1F1
luYJFEvGStiQenrk+mSCDnyApPi348yX9Dphgs5Cp4jZXArIiSPdFIbiN3gtPhq2N3b037tE0R5w
DUOl9QXntq8hDABHe3lWPCMzuzdSruwnDz1lh4Q1o1B5ng2tEuywupEeMTsT8jqB5Vj8kohq/QsW
OuOmGyW4V8eicziVwsFp9GPq0OCg6uYAVVnyc2lwHNoR8jSmNeqXSpvt74SpU5gzQJY4zMw/53hZ
Gqf9SYMYX8IJ1TLS+YMpvozKOFNfFH3qA0UwOsiaL9D/FSumGZ+WJRNMZ6BE4dgxwsbKps4PL9eG
qcGkxdoAKRaMf6KBmDExqx4Z+O8H5xdh5slA2cH+vnXGsXV0Ns0IidexGQE/ZpaS93ip8/vIYACm
tSEdoeyBWETYjGZvl0c9o58B3yraO3+nMowf66SV8XEIJBDXrcdfqPgjvUfcTA64TihHA/DBgG5G
gdmaRRwmtSMUxJeJmxlyIYw0b+V+G5pUZ7RzaPGXVdFSaaARX8BXY56GjmxPaXXYoebm0IKP2oIt
ssH728EFPHf5tyVitJxHT2wBjJHt4cvf8NTsY6npqLjicI0v6SSRiJkLEJc/eWKUJZowmfzxRaYw
2xp6gSLDjmOT+eUD/rJztmKxC5wLEGLFY+LYx/l9wozFbl4xMgVosh9Lf/OjL9G3VQTmrqe8G6PM
mgNm1Z6vFb1wEIVkncIMti20Xcr5bKOb1FzHesScKKC23jLL0SPyWnJRSVueRXtUr6/nn8+Sho7L
L5fJTaN4ikbLtwRqMKwbBQB/VLRpybUsnnI2dglUB4sU0FZzUEbM60T2Kne2p1Mblb0UN6rX9IID
CadnJS5j3KCquAHI0xEjdGr9nA4y2XW8fYwY7b6Exqgpq9wbV99ic+nLaEDA2Tjkn+/EdWClRJNz
QY3GRbfbKR7AeZPAYrbXbottXEF53BX6D1Y71gGiDJomxYArl0U70RK0aR3urXjB3nplzfrP6zdq
NdfOnQIYxfARKJSSc1dmJr2b7zLbj9AiwLjJ8hSwkNy1tpkSQuZf2WvSm9f68AoUIT5JLMPVx/eh
HvgkHILOIV40kssG13NzyHj9jjcmvhBhF8yDtzNmMzs3d/pvpD3V7CrA6sjYo1j6V4riRZBxVAqo
el+VUo96P60Fb4SZiknlJuPaCwb/mP2x8gRBXYiUoXxE4Q3EK+R31rog7AS/sIW2G+uchanT3gkt
rmWJlDLoZEA9wuJzc/ZXzSt3pV58982qpH9R036L4t+yNSXknYwCgEHb/inQUYGXCQwETrc0IMcH
ncfeEOGyk8c63WkNOd2TX6pHOv1P3mPDZCJbpCQQC4dJ/FlnTq2JFmP1E6kCohrQLfvQz4qK6kJA
dVnrNhn1Cvy4DHl8+JLhckxI1zARwzrQIU1YYaPzy2Y3RWqWVOwbP62akXZnER9WCHDpzUbBQFjj
/FIZBsCN5I4Fk8ujp31SSY1ERvaafxCpHCcDacV0kh4vmAL3qFLC/iOu1uJHyzXRvop3wvZFkOKA
07dhubpwsDnKWLx79z5zYBXXbuTKxviRpGNJQUZNB/jAk843utrb+oxRzePIxTbpvLDyv+JbYvNM
dmsSmOCT0b0PCEVW1voTZoP0rtQMjuv0njyAUpkX1Y9JgXIYrtXtfSR71fpC9BOVWu4TzwiU16/1
BD8ME1LXwkjwJ3OL3YhcDlEGrGYiRuTk2lAa53EjUMlsXvHwIaRqbQWo1AC0QjiDyh7Qw/wGofOV
vK2v4uW3HaTnbBCN/ZH2usFLYtefKt0M+NiDqNsoYBKomUsygOc8RWPQUjLV44dSBaMkwWooy6Vv
XFhoTzKdPPj4Pdx53FkTB193HQu9ljxWc9eWz2fro5zCvlpR4b6tN7e5w0tAwkoPkP+pykiUfzQh
y6Poqk1UAydevyk7LD4B6R8jmbOATZUiHhDhIfE/WzmFOVq0xiFPh/I1jZuAdu0yal5cOoDgR2Wi
1HHZvRsLuW/2gjYnDIAsgl/mKf8hQ9IifRYiCZHQ0wH47Jujtfz96bYunZ7qefkJ5RGCD+vd0czd
CtXqOgkMfZJ6RNLZksQS5cathsPALn+1LFVWXfdo4Pn8viT9e1TqFlbrU2/HEm/tWCLn75fzP9cN
DNTA53UGVxh9+CO3xFc0EXQCmJ+i2SGYWTdflTfmc99PzQVU0JZCxuguWEi9jFQRKLk4HnHNenpr
F8heZSI6JJ+HPMK/fvxlT74dJJ52eZU89Sk72bViGs7IMONZUGmeY04zZOjh7k4CqGthcitO3kgB
s7eLzprSx09IZECe6treX1Z2AiJxE4XrxvCWxwx2/6bXQ50RnSLFObZcDz8Bk+0sqNqgBlReT5dF
SYk+YdSvU4VDsk8nVKURr0eF04Mslj7iCYqVvfRzdhLVlmsGv+qyppmJGPHG0bUTTtvnCBPM8ISc
DunIaHO52pW8asWK87xc8w8a8Dl252UcbhmyelXyOKUkPQSVV58utt4VEOhGgkSDRG9abggjSNQf
2bsOPlZMgtWDArLvWdGIhZibQwAuh8sumwk5fBKkNyzKIsfEFPiSeDpFg9PEJjak5WE6NpGxUVzO
saDc+0m0ceCpuR3PKk2G90z9S2W83ojzFqzuQ+bu5RDg0R44d8mnKqv41LuPB75zTkMPsuKnLa5r
wO0zNtEx1abN3Ar7qmNyaeiJfFDgSQSAANpvEj4NfijW3GSm4IXaBUv4V5cEIKFXioEydJwlB8wh
Tn3x9GQ/AsjBAYv++Dq7Op8cShg6j/LfRowFEYRp8rpmYsaHN35pRNNjPntsi2dCtI1dSUK6YTcl
IToVhSTPIIbvctNAjCqVmiG5GWghH0yqa/ZbJk7xsQslfnlwb1rJNJEjRXiRnDm78mjSYGZ29RiV
VKH5dyaLuWAlqrqeilDetkKM9azrcBsQ6vZWr0yYYUbaEr60AaiFbhjNlBOKKHOgW+l+Y4xm+jGx
1pAztJ/L9KahclxFaFA89JwRzzwy2oarQVAb7RP+FH4kuPRByoJ166Ggc6QrZZbtkczYEO/o0WgY
wsH06eInCDdup0jFY5lK0kN0e6y3ZYwNqcKVB5oBHCmM83py8QrHfy4Xz1/CaeulWkiJxyuK+D3q
9mpjGdYfPVryiFXW/KudrLVtTS8SZTADn3QUHzPRDQgreM3nTFiRLA50tYITTFC7Uap6DEbPir6C
l1NvHGlF64mGNnzDW5HPUf+o5eEOavHKv2riVVbSSjBCGZD/jrEAFldqlxd4d6xb0t72rgoNZBGi
79Bz2x+dqtAyAmuWAJb6QH9KdYzdiLNCUpwg++Jc0/hFC7wq5Ll7uNM/gJq0J2v4ukf0m9mh8Lnx
HkZ0arTbbDVj96cEWr2lswQRthJfmpdicufiOuM84WZlb9Ox4Rl2gtuOoztuvuK9f/AB4O7neRPK
FXLGHR5K9InDji0qSTOInAXLrhXSsvnZV5FeYhdQkriY75fkSpBpwLc4HNtB4D7uyr7dfLV/fyQx
xmYOYuUY+1hAXFH3BGQ0Aq5JJ5iJZbiNbHq92ZL7EPTjGQUrxZllHOHsGCT4R+vIiiwDflOh8Ooq
zlWd1q+e0bI3oc52QowuUpVDg8ttG4gbyq2UmdWg/C/yWfEaLUunKJTBA0C2muDm3NNOoYBiFjyy
EJMm0aHu9/JTFhdJuF6F0mRpCAReguiK+CSQpercoo9GqfZ5Hmr+aivIm5Ub80JGtDfT19+is2nZ
QCX279hyJe/YNU3zfjAgYQ+byn5AXJXJk4NcX1WJlYrWPLJANTikzSS5U41fJ4KyDH+x8SeeGPXb
aYfk0VFxgjt2+cKCb4dnmkyL+DXH/8s+L/TsQwi+s/M7Ni5wBthNpHXk5ZEVsGJjHNC1fYLb+Gfl
eXONKkdcfIATd/egAYfgb+fP7HO1wSHwhqKvz+kl6VNp6VS1hHMsK0rpgxWfS7jRGcBE17xm8zk1
Rt3nx1xUaYWHrXL9+Cq0Iezr8LALD3PFG0ANOB+nQ5XMUs/8u/JTJDQYu/68PL5afqjcOBYBOzfM
HWx3ZT60o4GX2/ga1R/SE6rmoUd1sbGLBNUOUrMRv0UImkQh2hnN0Uz71WanxGe7cTt6gARSGti2
WihS2MQ6pAafczEwhn2YO07nqWyjpoh5CQVYlqPNyq2sZ8ZkvjMUbvAYdp2rpHqUymvYjfoV557A
T6t3myMly+tnefHvHFs/IHPDFeyz1ndcyyrDgqUjt7K0uMFFRPiA6oYYvT4wnNjwrsWjEAs9wLEO
RV5JTfkDjsKpucZlqwB1HQSFUZXCa8FyNOtNlYcCKTaQjVBQUmPHY7D6ky/9rBOjBTABUbTRQx6q
7D7Q/GmqFUal9jtX4bhj11/U8BJKaw54g05lreIosaollYsSAyyJ8okdjDOG91ByqqhqB/8GBLcG
651F4d7vebc5brWhypgwztSxsAWx60rCQtfrW1JhJg9Oym7kgGLQ6sGv8oBcQ47U9eTWdSHFZB2B
3kXzP3eeoj+nuQ+CPi3VPwNYJPfjV0m1+2N70Cf0YrFbqPLH3c3bohzf1d2n2uyaxMAT3s+ULi2e
IIdaortTYRdS0KckqhNKk8Ngl+A/CjlTZE9US0EaZ/99Z/B7NfpVqtcTXbMelFAyT5jTcNVy55yv
vOf7gx8vil17BFd0Jtct/yj9gdWstautnLFVRtqdzUNbbKDLBSVwrsW2ARTYLCWG1SVCAL37T+Pr
OFAwcVZqN3af19gRX0QbJO5RretMlyXZPhV+Soz+8NM9OtwN6yUFX/HwCOUbrmVPfMrUScNcYRHC
ESQaATiRo2aR7MZKWg+RY6tXvWx1bndR+JC/KfoUuzQSU2Iecwy7hUO+GCs0udpv+PJz06wSkLoc
7N12ERA35ZsRHJwd5fn96/NoJIiYxZI/NhSM6ckMb27ImQZFvUWvkdVP5CsGpv3P93D1MyEvmSAq
DkqEvyiEGHsfzDCQ99EdFqlmG4Hi2avnzJyeUnnXyNnZAW+21+CWvlFSiJPEJMws9ERn6EAHClQK
zDCOdx0xpL7epUe0adzvPr8QCB5RNy8f1Yf+9087sqZvrFuMm+c8yPxltMj7eYUhEqli+UgtXpdR
R0D8UGX0t4TG3lap19Xiys4evC1uONLH0k/3pMyjLK+U1oBNeeTzNKeFMV105f9LHRKJV+hdvmJz
hpIGIidpm3MVnBLk4PagoqpceGGQoFjZ3OtS2R1W7BUBbv8p/IwQ3GsIIO7RTtRP7v2jQPvQM2SR
8Ef61ICV5wyXNxM7JC4FNyW6IucWGgnzMertdCbZNd7eR2juDDZq0C2AvIYf4gvVd4u5iLIfUNUQ
aDzHgX8TUnGA+gptfzSmjSDT1FcAwff/IYkwcMJF/RT7VT/CTnSN/s7oWRzBNcRvj74jJVn3Hbk6
lg2MD3ioicZIFfpD1kuYIYvInBVzJi9jMxqTWgM9fQfZD7jwHTt5WTRAXA+V6N+/aU7VQyDmaLTx
Omn7FurJdnHRDSnG2HEbzD4Pu2qEPJjO31i3c81qZ6kBx+ByHVtXM8KxPLeT/nehtNz5i27j4b4u
BC7rn3BJVGIpw5TISo4oyk92S+jtBs97Ez8qpXIt9q5a9774pKRWpC7NToCPaAXiFxifKouGZ487
sgRgBzjhTnD6nmvUXj8OVShxfadzum1SJQ7VvJQyCdgpoiEWIagv2wzgwLm59Cj//2h+RPb84y2U
LjgZ2FT8/bNlDERpUix+IFkyXXwTWGS5rEOLrkYBJHXk8bEU27mnxPTitUmH+dPjF57XJJK1TOk1
ZuOJo7m+ayLW3H7p089Vhyf6SPQ0sx/i92n5Q2KIV/Koy4QuP6iLYbbz2ONDtZI8IYejaDJATxpp
SoIotqIhbZbb/iZgR8gGZixLloljEbi/DEWltLQL7pquCXlWir6339o0iL5vecG0PScyfUFKaIMG
y5SK3gJ1wKfNlhqv9x2mrUXVLRuPw5MQJ9xTnHDFeaLOddqstz4f7m54tu3B7UpktPGJREueM/RF
Ln0UxZgb81gSpYM32c49A+3wqFv5cnDVtxQORfazpA8PHk4Pvt2X7uG54riKMjozidDeVR6eGKKZ
m3yrI66G8d9A8LKuHs9ba54uBaRo2EytteFCPPCoqyb+sv4D6p8ITlOK19AOtzo49qNcpee9JGn8
HFgCuuvMWY+poNinmC1Ub0Hqh7V567kyUrKcnlVkw8GGdGuEbySIu1avjLXW0nxb4bLQtGJDi6w2
UU5Ul15REy2uqcNEJ4bKChjU4mQZBKLc/v5xlWhjSym0AWbmmdTwoEIZGG8c3b5Pp6hCUV0OZYYb
Q3FE4VgcPVQbs/P/LrdImM3e0+vVRcuLGzu15t1T5juUqcTd2DKIXAW1n5TBAdLlqXVW7kRZGUqt
oVBWRCjtgxQpiemtie5yh62MlX7k9cxD8IUD+K//vqSP0F5QZgxc2d/1ZcPG9IAbGUnG1UUI29ha
7d6eZNxcG5s0xm2Brp3Tsay0vAZFu2LRm627jo+i2GImGFmH2WXxdRI76DDQWjMBx+P9bngIPIIs
X5+giJCfLFn5p6Z18qy/9v8k0TU+pDo55B+RQwj86J4hepMKda5ecOm0Y92pIiUHX/jpy7F9GCUW
RMAhbeICqGOapwE15jZ4YboOD6iQjTtp3AEEZqkXL+9RxgzyrSfpB1qfNGWgSTSY1RX4HZl/LgmP
sGg3XlwBVJMHtPNkUj7q/423kK/7cZo2qdlY3x9ktU2MeotOw338OE+1qTP1pCjCFHG3/4Xf8l2s
VWzISwViX+oNfcxhq4dqusPr9RO1yGo+ghVhQuhex3Ok40m3Q14Mshj4BhwP/RI4SZKnMMo76Ef1
CRyRxzGOxL1bS4uwftnVzaPKl+L+t+yWx88DjP0WGW4he/J6JKRDTP/KR3XDuljLlPy43abiXkF0
e6uRxQ0wTmBPraQEuKrAVhjKecvQsSUUoPpjaqPaPkM3YJXNV3IfrMp1Rm34Y6W8PdcFrA3+qagL
YLIZ2WGfN4+mS8BZvIVqVSMWIUeHvjQ/5R02KxY0DPDT05ywlaYsag//lqmF+OR+lRS5U9NCth37
ohEdpiMoAJ0baDR3m1JXo3gPnmHdJVcxKrr+Rd7avoBv7kegpnKmjLMhXQ5wJbmZ+Hte6ciNfI18
XkHqZB0AyxlBSXtjEuGqlrox/K/6sxxs4pNF8lVT0VHHW2eaaoqn+EweLIXlBjIDjdSidudmRS/v
orrH9V3DizB7ZuVpZhzDz/J5Mul6LIVRuWscEjomui7TR3G9hs2tKSnjuohqCDG4J7Xi1JU7I2eg
CU+F44zYNTaBOyEy1mmBx8ahjBHSDyvCLtO5bDk7qE06XtBajXbEznnE8kIoiloxaRwRtbc5j3sr
J9NLiXvFyYuH9cyOXFxd5JsPQOmqadFNc/u7tuxOJkOPRdtcvZUmJO6aq0LULsLdpbi57Q2fPkqB
UMDAq/yCwEasxY3zN5pnM/H+Sf5j3T0hfAiODw8gY/3z/syhMYbzlO3dHCQrhDj+296bo/orBQ1+
PV71NYyPMBn4RI8lhGO9KYW5XAcxZLnb8tLq8ucNQbzvPkSkGcAuNk2b8ihLW/eYBBIlb8j6B7QI
UeGUn8Dv020LJFThLS6f49HQqH4VpV8EFRzF1KS7qxFJnaADSaoshbfsKzTEoLLNA9p2FQ1y4uzx
EExS8ZXJ+hxspE2A0EBGgG9E1LDcd1IYHKpzVKaHiwlHZgSInVuIcnqYsCU+AM+Ej5LPctUuL/L7
YjS8xSuuLtU2TzqKcuFcm5DB/+Qu/uXfC/BiEXEJGuajtKNBr7zSYuWqu6T7Fam0y+9JeT0CR24y
hgVkr8pBaL0SCs1rArSA90XBAxOjUKUPhe2pWg2ctzhOKXw6vKE/nZbdMBpJ4DC1TLiqG3+SKbnU
FwgR93W2ypmXJXGm6QtwQw3jp8LIe4kuPH+q7giqVOIcU4D0sa6XXuhcJRiVHD1f4upPnTktXq/h
dDcV6WFqdOszXJBBtv1vCRlZWYD62eOpHus+7AVxnRj57Ol8wrDiSJjqNw1w72qVRh2k1W7fvWnd
QPU4w4VosVUUvmePSKjOKWTdW2xb3p+117QUk99TRGjFXY2x4ilUN+bqQCq/RGDSs4xYqxmPBqYC
ZJwX5hvP5tFDUbRj33+kzTn9UpijRmsdtP/Kc24CIt5CDDknarA9nJyINzKElJlqyLz7/XydVs5A
pebwoXVbajbWWRMvAGS/jC31xawzUoLUU/1M+jRQoPDeodlVjJu16TtxmhFvgQzm1CVMsQUs5OdK
25C5Q2e1/JFYOWFpcfkYShtPcDnemZl6GFklJrmhBSzKkAq03NBQ+Wng/pKWph2HkhxjEc7zETYl
0ryrQ8WwNmLmKaWbzsGE7NyrA9xRVo/QTWqMPPEWUR66ueLW35LtbJKH17GjTk00fB7aQd3m3jwE
m1hAvaM0pOkiU2xWonWWs0sBz+BtykV6QgJKYE294nW6S7pom0WMD6NW2VYGXE/DAmtJ1/tELUrX
LupRqkFG8f1ER2yVEzC7Yp7qDGksXdt1gwm8FPWLnJMFo8CiJBAJgWTR7ehsqlRLCKe+eLeFLn7v
JL4PCmbAiejv2j5EcI/ehOdCUiP95XllegnZ8EdbiQuidn7v+U/lyVnIePFDdVLaDquQk2tsqxTw
EDy4BACtA6iWSrMCreTQM1mICz1LFbCO/0mmBzZqHI09vFtbkauIqzOZYM0e57jms3a9HSOh/qwe
zSW2AbBxSf1qnUpC0c29CM8gKFFm8EfBX645qnuIWCaYlT8TqnXteHMk4I6/Ofg/jIOKn+heUEjx
iARjIajry08VuYehePwssRiDv19dPbVaDlifuB4hsj0nYHfyr0Fr4p/1zXVJis0hAkQkl28NqzEE
5ViMP492tZm1Z5/5c5UAQewVu7fJQr7wxjEmLxUUOw0DMSRHixXrlYMXQXUIdwGwKgcQkaLNgNQv
+vyKezF4kTCc4ABQPjXyGVRBe/V9suwWtWmbPUI9F5zrfX+3ZxvYL3SmfO/uAHla30PimoFlWkqE
/oPUOQLdgWphZlD02Cx9lPH28jVYLHZTH8QG6LWSnvbia8gKOtJnsJI2BEEzgV1MStRTPMbIw01C
T+kwvOw5rucXAV1BzkdfXBNc4K1ZVcc7pLwMAqBasZEs+wxOJOt4CCGq0FaQwo5+HlMOcYQkZv8d
cVAmfKUmbgZBxSMch1GgGdnQ/fepl26S55NE/h6Xs5UpAzmLykjpUlWN5HONURBX73UsE3yMF88B
znOgbzVKMVWP/Fn5H7WteE6g0tgHqWO0MM9NIucE2b1kiDLsTPFpSmxmbgpdBXK8nuYdRqpHrddD
jdWUKxsJqYGCBRpHUhV6ezHWJ6ACZWEqqCGZMpohFFVIJm1haU+Vb+X/ZEo9wbt6mi01KmDG98C1
ekpaWSh4EdF/bii3L7ytsIjqdEFi3nSmWC6miet4EpNV7Ai3fXUBDBClPy9ALMKAW6EMk566o8xU
wzK9IZR2pWR7bLugDZKtCqYyZTLIgfIDKMwnRu+ANjH6zMtldoopnqr+Uit9vmz0xthOKbL/DUCm
UI94kvBK8qIQtq2XvI+eOl2EQkL2wWjC4F2i9p8LkqvE5ogqNpUFWh1zeWdhbwWzzzLGstgOG+aC
+3kRKlg4bV5XC+6zHPqAIaCFzw9DdLjdy0YqfTRu6e1a+qD8K71sGnhfNBk1vSB4URrSI/f2hlgd
3V73SJPB19/UDy44ZpaTyfsP8rEffp69wqxCGduAqQac2TgD4LrxGz+sH494DWgTPQkYLF5+BpSX
yCG3HKpX5JAgUPNr5Q48uHSNIpiL7j7W+VCWhl9xfZpTr6CqBt/zUoGkr3Cc0bpnUoPQbaJUmnOf
BdlChyZt1J7DumRnEMxW7gECTzF5ehjfgYYI5C2TO+6vkEy2qioPZhZIdEsEF72VgSQIzZ8Hpvfb
Z+2Cadsm6Yrv2bcqPtsEn5babTYkqnWDu67Lezny8MbJUy543x4Q9dIVhOy3gB6N7NvwZ/xl8rxS
E9Kvlz1cESRJ4nhORjTV4UXuDu7q5nbdA30CmCC22lDHYDT1T/wfmss16nkGKq/DxoSb9OTriZB6
tSCK/QdqXXCUfKWzD0jbJc6f/ogx6cJ5s+nqGqkidff4I2ot7vESqszhsYN1VIJJrfba8dbpF87Q
AvO1PflHwtFnEZj3RL8JaJe2T3e6FkM/NFz/Z2h7f6HLhrQ5zTu0xLE08T2AlHQwqFJWF4YYAGps
ci6UQqeniVcS0pLsIAxk1j/4nM/eC6nOYA0lJI0s5x81E0LDdEPRanAIKlGGo9potensTNqbipPT
TKW7Z+7QoZ3WB9d/xuu7UyOFVLu7xWUtRWvs/cGawtLuxcytSE7SH4wYkAd3EESUMLXb0jgUoXwz
OwPF10ctRWT2xmJCx0QGBYSQqN7Xc0pxo11zAAFYu4X8GSS+Ubmk50YCIhklf29jm9F47xsLjGeA
sAFJAPJW25TfXtdflXd4gq27NymL652ZSwM6gYwWTK4H/sgaLA49A9rbxjO2AAMIV2i8m73kwoel
g2KGG+OPSeX7ty7thMos8vWjTedeEIpXdzcyPen9XUoaGSkAxFP2L0xpdbYlJXmVauHircQRUMiA
BNa0mZpBiiSj7dsuTCHmVcFlRv5E/JK0EMZnGWTBntAKevy5ZWMvKXfotk8H6rW6byXKqZHf21iX
mENNAA1AQFmXwjB3/7JkWziF5upoOqDmQ7S7aZUTInXNWWVZ4DRT5ei58SCs+bdppaAf95PzYzwA
0jUpIxbtSg1wn4KtsLDxv8z1PVGhYzBzoBARavoH6k9qiPBveJs0zTEHy1uLTOrD6zwja62aMXKo
kvVL1lj1fttywtAGI/Y24vGbfZJKvb4Y7zS6uoMYyU9lFxENV1eumS0V9zFTvLivsyJXeUMaW2ZR
NAYEQ+o95PNreKlWupzWEoQKqWVTBilcOmPk1AO+VA8GcGgwRkEg2BdwWWY8y+qr26iHm6tPT5Ks
XOH5C3Gnm804VO7Z+Vgzr3IwVnPZxfsyEXxl3BzxMWWCpSeEbDxFrFsF2LmAbn6IVLqjIbvPKthG
esgr5EtnEsiKEjKqsLJOIQiefB9IRB90kKIelUMTz+WLp76a3gTHgdhRd7xMa6ENxzDXAocSWmeQ
TUnCYgW+O/s1V3hQsZtPaB/nmHpPhUimeFT5ld2a/Xvf2kl67ngtGrw5HGWJIZoJ1uSAaVCoZlU5
YrSj505uf39TwCyK4YuJfr1/qLaPFm3H6fNE8RTEkpv6KdsTPEV31wHwKhFsiWM7bcH/8+w7Nqmv
gff6VQT6QXbWX1S8SaDmXPFJfyVVwfdhF/FzEBnz9eyoahtn6i9oDwWhQxGwKM2ZGYIbY4cmHzmg
7OipttVxKy+YAuegiBY7xZO4BVhOrJ6Kb1DZBTcj8zzYdYs/3k9BuLyVq1xHvDJS61BlGqxZ+IIf
u8dx+2+a9J37WrCb9hcRI/oizq+L0Uflf97K+/SYepEqitGrDofGM44hz3EO2Ty8nxzOuSf2HEPf
ISjO1SRCNNKj9KVWQXO/1Vn1olYZVzS0fdDZBGdZwwT8ik8kKy1F0APPUyo9FY4B7eYM7EjXHwDv
R9lzf38TZia0YRdGjX+YWkwGYHbXRW6kvvuS55cp5YrhYxPac2ZyY1Z0NlmnwjrNS7UajtPY0fXB
OSwO/N9mhEYSA8KC2t90tsMqwkEb5gXZ/WjIPrkfp0NUC2VpLKakOgyz1zKCl0PeGV15+T1T6qDO
y3+pe7cHt1exdCvJ/84MJC/l1398K82YhNMD40RqxwiZzG+WHZk8A9chc5L8cEsQR4OpcVrfDG1U
0/6XPjm8MYNHM1FC0Ncsl19X7Ba5pYkLxjFHHLcsl7M33/VrFn424tzjXMLNpwIrsbeEZ1AUw9VL
qGgJkkG9MxcGDbZqeG6hRBNDLldZ69NVphzLgOCe/jy47m5tsVE/DKL5XueDlQXdoXypg4rowaR5
zjOBd1HfpOI2CGMlBHwagBz+KdBKLoI/UCpxUXLSVwYBhV05BI/We+kzkkf06fxxFiAYQIQ9bKmF
2KlS28vzGRBq78oJDtF3K9QkGPA3De06cJtzS5577vgCBnQtxX/hqtvO03dCYMeNEo0F88laWDQQ
rlMzdcPYr+M/3Z3gJbQoJTbEGLYwhzLmq1VKvWa7beHCTEwXw287emaV0TtfUXrZGXLrQANO7GVg
ucXysDYwXS5e0/wTHyNTQk547osnvmyN4yoWpoe2WqVkgvRgBSOxK9lqlrfKIohEPtNTDcUOzoBo
lWjCK5M0ypovY1xg8YdzRp3zwcRGuVdBrM1cE0G2WllgOICwknz2V15Vf0OCwRZhHGj28ejgEq31
qiJvO4kmJ3/D2Pa1GUfG1IGwDG0fGo8TVzPpz8L+OgmKcy3R13JN6of5s9qizQsOBM5spTbLFbXN
/fZo5jj+4dBgmHYSLXH1ryXEIQVhacJ1CccResceRoJbAV4pinhJ7OE9tL4rb8wShL7wyJd1+dAo
k8S03h6cJbZoVJsIpjpxJfLvyv7664smuS4eZHEI9KPi0sjTyayh6Lh87+rtrix4in5AmMlUeXkT
qw7OqrzfwYnMtH5pzzK5A6QNYenJaMUvJnEOyxQXEmurHaMCKF28dUc1DVamj/JAzlyb001yWs7z
J+K55e4Xs9RKqs2DmQP7hcSvbA1IW0qkydfMmvq7MavBe1MrTfN5PvckLdJVD6ie0U8+YR3uDD/G
TZjWBW2WxocVdFD1g2msO3VYRIhaf/0a+gucXSxwzgoiQT/CBXjTI5ANAF+FHP8fu3eo1VucY48A
XZZuaml4BSZbSkHSoI9XaShZQaVRJt+hxoOhW/Jumz/PdTQghMMcsR30dDKsw85mAGAnPQKLry5p
29qfvZJ+nbC+JX2Ags4/osLNXYnZ7j3wYmZhdhRU/Pt9qeOSkMRnjW7A2p6FNJdBH+TRMvaAxq/0
9dGb+mhZpmwEqFZmwC8xCMV30GPxcSQ7Y2f2i3Et0TZriR/AtJ0IYh9H1QVagivsJe6y0MLojZ49
1pAb6Au7yglDQM3IFftejA1tWOZI0LLcpRs1K5Olqv9EGIluTiXQycHkiABviNVR2nI0ulxZj7wd
KrYV/tyBNDoUueefT+sk3IaHDWgP320Xz+dQtTp9R4gm8c4GN1Ueqe5yt78CHPolsJSP2LVy5S+d
xIhcTqOPrch0shTheNoapukfOtiPzhlsUanjoAVf+SVWEeOecS6EXaqOLZqNiOm2tTCuKyzFJgRx
yOjlY5OWlKpmJWn+/NCjYUPbJKii6DVmV2CUdnMBeOZeuJ4HCNtWm4fl4YQCELekREokYBxv1UzH
LBbsOApgh2PeLBp/Xfxyq9ATt1Qb7NTbcN85fTpm8ohahXREM/11uL65b9zMi0okAwA9dJbyicsp
dfqyUk+eiC9CY7b7N00Y+7dhjxXDI0+60wusDqDi2XEJqRLV7vjktMChjZDv2efe620NxrQz/bqd
Z0/y55eu10W6b1se6Qk/aca50A2YZNS+J+igSSPlpMYSsbRRHgWLP1DkDDFcTMYhHd55lLV5Eeit
/EMPt4UlIW2k3yMkcxBU0onQcFFyy5A/01JbeRl7/6w0Dpm2PPLMquJ+sGs0S2l49StquufzUnWS
e5Y9kQpQi2tbHs6EcNzV3TDg6Hst+TWJsd5pJmQM+7s4pbEM1OZlOIhpJlEB0Jnn0WDK8m1lNxM1
hE2KY9GGJeMFc5u/x+Ex7VjOLRWfSUOM4xoxS0eJJrMt1CVhB/aATpI1yLw8YW4TOZjQ9pRMgBxA
/e7cq96tPqBQ/2jll0Im9QT3W4N6ceOlO9aK0T2Z7eaSVGL37Iwjr2WxRa8myCod2xTL8ViNiUZb
zYEZZywnWTjSoeDuUcCZHhd2FmbNzc0F3SPARh2WNHWR/NExgu6W1lVCl0GH3u+G+QEg66OVKee2
B9a6l9YefAY9dIgd4r9U702CpJbIjk8QJfvtf3K1kru/ia5YVxylbBmx9H5EdvTlA46/ejqPcCjQ
+MVYK5jGYvMd2UMeWJVZZAbfUeXBDZlov1jG+UPoq8v88++dJMdZlx0WxHpbnNcqDg72BL9koRyD
uGEvuuNURISfaSlVlQA96sWupObUD8f5YMsmZfa5n+sTzYSAoEKyO6wBLR36l/qdMOS2I64lRGqZ
3WktvnaF81U8jeDnHPK1J+/xP7jcw9pWKAA9xGm+MD35hYnh8AkwvwjZg7WaDs86NFbO3M2L3cV9
rneHZd/HcDYSuAbK6TUhIFk02TEAfFbtoHNEIHbI1h6X8nKF1ylm66EJKVZA/41+Y6g+0siYk5eH
yGyDaqDNV5z8slW4IWVT945cbAYsnbMoYvQz7DgAI5TyvukBoMklXNB620ZOi9wV8EjODsfV550T
hQ87Frcj5LZV2Cm3bIfnk9JjJpS6vjGQhJK9giatI2YnEQ7ImJhqKWRYAKo6x17N438wIkqAuEhV
pZBsI+XDUB0mlwVwOAWC+0EbJZmcBsHYY7Tj0jkGHi5XrspXETgzZpC2Z2Ma8Absw1UhZPCTFa+6
LvZA7DKYHdcMX5JLyyCnpT2BriTCzaFhwSdqKq7l/QMQiyRL0yysKbvhxHGZ0zJQ7/2/F8azfG2u
JKA+RAaUrZfG6wuyLoPGXcjIDFnx30VCYVAm8oculxHcnQT412JerTrABPvdkqaGu2dJWPub/Hq+
S1pSSiC3ctdREgMPHhjiLjHr94y4a0Rhj2J2J2T81gkhgsHfWZp2fzKdbVu6Dpj5Bk+j2C3BEvTl
IkIC0zqAtrXyOSPu8+eUwHelVsw4oHrF4Qa81xxAMph5LRbEuA5Z6k2KZOGEfQ8F4feI+BJj8NBT
SIpHInQ1lG/ivL8MKMkcCrdtXING7SVTLI8FOmgyymtIau7QU0lSttM2h4bYRjOcAw9TiUxJiwIF
TovFbM4ThZwzlyQFdlcutfW8hsr0IVIW6LQ8l7Yt2df5avBCIkwH3qC4mq26MP2Wywl9QL9JqJAx
7MupZNDF0kBuGVMEv9M4R/yMyx/wQh7e/1pt96gJHZ45NzBM7S/jLmpqCsH4MdDr1hr16vOazMoP
1L6d+WQADpJlaxaBeGyS92WPuR++aUCGFo7lkH1z3KUChbSPIJBiRyN4/Mp7rLK7B2O/R6QID8Vy
ZlYrzuQQ+9SN8AfG4LxXH5DNYsyxibeeikLccyJa/74pKFx2+b8iRgBSblYL1kAL9ysjwvUhtNN6
kDCQe96oRa1UP+esmIyhRIyQ01I7NbMewH/knNioBKB2dGinunMNEpLWEX3b8GL8W3X7GetRtza1
IQIEMUz0pk7g+/oef+WbnQaFAxgY3O8cxMW99vToxdP4182pbxECG61WJR53wtTBfB/Sk5QHRnkc
UJjtpSVtb+uDz3DvAjBZUVYkAA5ljuouDsHxkRkEJXbveyI/RkunEvVzDnoNrc+zb9u7TxfRk+RH
djBtRPvKSghK30vbwvOnntATmZWXWPiEDagx+2Fdzn64jbNcrj3CJIMT7qOZH85g3VEmbty9QGzD
nCaelAuJNqQvOjApKkVwaLPHEQPbk5AphqaPL6IFqRCA8z3FuWneyQ7ay1UdWvUMrET2KIXzWihD
bgxad/970FNPbuZtYuwvWx2xenyvTbWIzVQCDHI7tCt4RNIn4vE7otsV0NBHtvQO0TRM/lJw70S7
EgQFPC4rNCLiBzu3tlwpGDEVh+Dj8Fb9XGcqHU2FoCxZYMVYkRlT6ya9VmXK2RiNaVKyapTNgoGh
adL2w0Kb2ymw6daU31m6Pq6f4pQ5P6AmsyE9n1Ven4im+YstYNTA+HHfYYQsm9XaFpi1JHWj2TbD
zyE3CUrNgZzk8Nobht2XuikfmqpadyapxzgDPPlcjOKv35OUf4+2yv+0b4Daf0iz6ZVy2bPy+VKZ
83jbLrmRecODhgTn+gMWn5BQ5M8fSJ6IJ6aw0OHpGAZlyhxOEYPcXnwqZ0LgFEbljPF07xbuHn5I
BNekxXmWU5trOlWuvRFfkK7EgYDNMDshBChjAjPPPFI7OYwLxsl+IbxZJo0MmzE1F5f7CLKA5nPH
e+b3MW+ehjK8x3Z/0EwB3MtIaI3gIm2nNKpsSvCnL0zxmIb0AN0M61c7O1vYgdCQ1exqTPEZboAN
hT6MqyLDQ1/GYQmUtyRjCT8sxfC0b9NfKVrUNFScXmb8/v9K5OJ/ulXA85FmTMUDMgQJBvvzguTE
+GI5aS7lbrMRUUwGRL2QrDAUAcT5i0goCTNwaBTtIWkUSoIEp7f1GOGVXjAXO/mUkOLmFKo/ORTc
BBGjtED+W8D5GUfmVrKWCbA18PAFMGmajRlvyw/+lZend00yCnxi870fCdkoqapIk3ti0PW3CwH/
2gyNFpWvRCWtI1+s6BDrgbpHheeZbSaJtI1o5olh4PJrbm4yvM94LxEIDMOV/12JM6HMbGjTakNc
y+dlFUcMl+jt9dYFqMwWnN4B2aQhlOnUdP73EZS+/TZi1QgU42IHlmb1Qrca0EXp38BrKrXhHW/d
O8PfcbzF1CJCRHSXkfzOOVlZ0utZ7L4jymNMasw0RDDG4xOikG/4FYbqwo909Oo64USokFO4+y4t
BlYvhZc11SW7paQVnZVmaYvbDVNQKXn51fj3LvyS5WTZjlOkxuT2PggJAOw41x7Pba94ABPHTx2S
qkq0ZrknVloOClsW4aC9UD73fiKxsRjmPBryVBbYsBldhvkuVLe7rbX9qMGC89HdAt3SOnGEALnN
shOsTi9HOV+1JqhuunF6Yog2loeunYy94RD/cWpcXIIea00mgeY5WmEPRWARRaXdJcEfNMrxxPKv
sQNYofVqwDIBah8yMAhlhoU4D/nWmCNb/8wTCt6zKuPeSQ6GCuHGthWI3cDVrUBla4v8+6TxMkVJ
7flR7sb4d3hcHr6NkrXs5tjjo0cI/arUV3fXgcAaiv1zbFKJFsxC40aAWdXEnGXzqUbw+MI0RL0Z
CDAObFW2wPpnvOXP2JO6A+ZZMcZB+ccdJb7vc+jN1pvAXCDAA+d71dQa25JP+mqPtXC7PtYiKnKx
5rRCwZvEq5erS5zkly1zQ4scpxY3F6qgWewD4Jo4EHRPdclRn9Ia/Qy641qpCzfw6HKbDYto0hlZ
ZtGdezb9/KwATy3E6I+W1qGe3sJxcN91pB6ydqDIUabAdIuc2C2mFU32h75gAa7v2ifN03ej61pr
SAQ/vaS/LpxRYqIeeU/ertvYAwWc6p0xA67hrpFWMUPD7fRnlji8JSkmPTOFLIDJQ2PFyOXwXonF
29D5xzUCC1zIL3tPRX8KI+o6fOo0RaybS3e26GF/EdKm4MEeM6gc/ZSb8GuQlz10ZVQO9f4WQ4HE
GRnG3fKPSOZWscBpGnc04Ghcu8/8BOdais/GKKo8GJBmL7r28lMA0Bn21+JCZfKRrZs28+mcfqsW
yPAs32rgz7yq+AZG/QDwT4+EbnvdPVtn7hx5hZHcS26Oh729mtKVa9HXTkSh1pcAWfrjNCCR31Km
5/SxzSkQWARmKTrRnB1uh9GD3bq3N4rdexV/58S3keaFXgj9sB6x3uZ1c5BpnS8E2S3hl8z1matS
9K49QM0UOeaDg4nqAmWV7/IIosjRVICcW1yllG90mbmIrvsxUQ5KvkY0JzcQndC2r+Ls7NJnCbNg
RO1f7vNr8wKtVouQFgHICQrLpsYJLAWBIp9f+YHx8c33YMh6qpFPneApwkOZhTbsAate8iE5mmeQ
TZd2feCD83JK9fSXNvKNwAJKAOG5nRYyifkZTSAwxcfS56XT+7+5DXNgm+dBG4SFr4nmmBoJsjio
VuXIFOXgYR8+rrPWME0fBVAYfmsEc0UdeiaeAUOVnu6D0drzPzFEFUF3DkrWfVtD6undp0sP76ky
dpClw+UPu2ja8pY2xISBWs+gBYxqylkGXV5Cw7RGJ6FTC60EORf7cr3WAUadz/Hf3iu2V6Q4tXFS
cgMvNtT1ujJgVCCsaT7Ldbicwkuo3StoVKJkZcSzvNELrbHR1pDX6Y+euWLv72DXcnHlN6QgTNn3
/zsVy4lcrB1y/KwGdAtlETAqcncA577WRM9UolOUXRwUMYm7EUZl6Fz+7Gx0K9QpCM5WJEmSuA7O
j4Jlt9WqHRUgOkYLdk6MZYJIqpT3c7xFw2ISdmjKdqCMAFPSKTelEzdKBm1Dt/TNK3pNKHuq2tGi
kTLyoz3MwUZBeLaSKtKS0fvP0huGdfjABB8TBAFI7Q3KlYYKDN240justFmGxiMaj8vauYYY/6jm
KdoB/zbwnLDezXuJ8upfzbsLV1cSTjxZEgkRKv2xLlZu9hDkTCe4Eb22KtdCtJPXUpArCsac1cN0
Y51plKnb8sEV69bPErpY4nfrtLNURivIdC8VKFnGqypAg3XmEwfxm3Ti6sgTBGsQA9GEGlUFtSxr
q3nM+KQ1/ICWpplx3hW/GVguhERj7/bKJLW5pYEeAy+acyIhl4uN0EcVzVLoDwV2RPpPYayst074
EPiRBLTQWkyPBe6/xioQyVIlYTLlNybrayxUaDSI1LqbAU908ZpNWHeAc4g9RvUd1pp+mksWKL8h
7D+ZqiC5ZpXSvIKffJwYoe4ZvuGR/flXQFWN4OWK3WOF9qu+Xp1DlmHF6gjdxYQMQPHDWgnCxO38
+k5ENx/aJzHKh8YxRxhMhFx3Y1uv9xVQLdUZ4aJQuY6ZwaMap5r6HoZ3bAY56QeCZIFKnpyBNhoi
zih/+dqcT2hT1hfk+xtOTziF6+w5SAQyESvGYz47UmCZiU1yEzNCtjw4SCNmwHtiHjVIplSvwpPw
SOqIxAu7e42lOQIw/KWdVvVZ9Dk9diKa/VnnJ5CNYwmzgPD04pLP/OwS0bPwXy7x33It5aoU1tAw
OmCu8Nz3cgxe4N8ANc9Al5jBSnm4juqJxkBcuAB0KvQkw2jGHMOMZiqGOCUPm/tXfVW5PtjrB68i
OZ4W7nBuV1wrSdijkBWDiWSYlRhTvBsHzJbmiIEiQ0c/o2J9VlfenjGSo1ddDmdTt3Mk+BQv2Job
wuCAB83DdC4GII1ABEk9beUGXanXBZzTFr/+mdG8jS7Ovh97IDDWjh3yqeqPc2u2JSPg6rf4/VC2
+SWV/x/E1vCOGy+ZdCs205iq1e2C+uOpbilIt4AOxJ204dtM+RkVFEK+9gAR+iB7Ycl65tFC60bt
NLoifAMWfwvg0GD3DHoneDJBBRl4gSiAFuLgn0WT/dNbda8xm5jnzMwzfPe0b1G0GPzImYwuBTyh
mazDwht/9D5Z8PiTyG1AAwhRFbxlnSDP54Yd9/bDvVmkiX5ffxD1xzs0fsrBlhrDCnIJj4zjrUx4
TxK69xNQ0pJHSk249NuGrglggueLpT5MU1b+8fPUJVaHaoDCkgydXP3RsbxW1pQaUb3sctjhnGZy
nLFx02dN1P3UwgFA6f90/sIj6A0TtZ0efqGtqiHXdtEvE2ox1XdyzJRXeq6VmsHEqkoVeGK3IEIY
uE/vtJufeKkrH41qWKT3xddN8oAvGVuJvmlAK+aWGFy/zG3dgCUssC3FzVr74Q5EQeR5vO3TVnXH
+1VrA8TJcw61mJiVJDIBLP1WPKurdohD2d0oLuEnWdeP51kZyOg1BuJiEULn1/+CsGO5L8I/13CV
yaS8Hr5z1zsf56F8nyHsYpOZLRP6lKa8TtjPbJeEqY9wq4bk9u4ws4ivJXBhOvzJgKW11hIpEpOS
+Ghe+PQOX5e3O+HaRMJUAfz3jV7xGTxHeJFxFpIydZ8bqxR5kZ2TRVaNMGlvie/eVVQU+NPfMxvw
jJR/51fFrahbdq3ZJqqmy/GJRDcrNKH9YMaxGntgTd6/HG4i+bJJsrmpVOvvz+81Zso6B9AWjYbh
wXJfgAJzY1hqHQ5vzjkeYWq80wyAYh/6qz3CaTbjK5mRDUbhHKFhc9t76m+zGyPAlwZqdGtsErwH
MkKgWwtEHH6SkdcCV7t/LRqHyMXQpbbxuPVO31ybFhLEj6HtR4PXYTk7DFFa3iT9bDL/PViFRgwh
NfYcjRz3VtcVAykiOmRn2YXbcwlpogxFSriVI6VvLT0UJbfxSHelKc5uatP3KsKfq/Z2IYFJuAIX
BoOkpgDIOSxOjFrN8v2FHkzwDktbK7qipKhoMS1z9pUqUfFjWvp5R29rdDGNmewDDjNw9ufPej2l
3KbdKPoHyIFF+jf+4Rjq6sYIlSJpXUaRKfu8KRwO2BTXZjsjkme5ZNt3CYO74O+P61oZLZd7NLK/
Pwvuv1e8kZmcyRXHyP5gZ0sLwSbYENuSFV/z9aNpBXZi58yVLTWfIX+WOqJALA4niMf1tEym5yco
uvlpqCiH9gtdGYriisgMH8GfZZUgqma3R5Z84Y1fhaMMz4Bp8jCdFCm/YvTY3Wa2du/A71KY24UL
CCfWzMrM8OmgOyQlCukpsvmg8SOKXjINdr59iMAyac5KczHxv1jMQDcIxRAfNUQlKiVu5YC4VRgL
wsuP9vlrC2mdRAV+jJBqO2D9saBzQOCIvSu7VdUkVqytU7P5C7bsST7nCXuCoPBizHRbQlNfV+Ey
PZW8+CbwxXFHxwmC3ui5Rzw/mCuJJVtZJBIhxo2wIGFamx/8a2p0Lu4kuGeWeKZijDQXiYbK3kNK
5dyGA1cS+BRyS6qYAsyLcpIRfHQakQuwdAas7BJYFdPSSnAqhTYV/EgzCoQzyx/G4MtUYXMZhO5q
Utbj5zqSzoSo6I/MH81DANWrxdUrxe2wYGSTJ4ZDlZqvEGOY+gLFMX3yAO/Iv9IfLjqJhZUwE7AF
jcJf2kVSZnUj6+bJjEWEJzWK0fXInqvMI+cj2pp1W+mEAQxeUm/ygGDDoXHv2TeV8jl1KULWwrcb
VgfG3hWq2NFOjdusGKC0K/NTN1fcAHWWWx0CGmS14vPIq5Dp2lVkxGrnQhzErdk1VeqhJhWd1toy
5QvdhBO1Yua1tJ93aLvgv6baF5lym0p/MPHuvgY1OJdVF3iSJCS6gSjf/PjGq+ULvdql0nAdaWIp
TLNiT98R+iksWn4GBTYjEZKdR3V6J6g+p2k/OcMGczlo5J9hzK2VVuTGkZL8wzQPply5ljhVJAv5
i/kAZLUjdS6c8z1aOBugwKobsieZUPrzZsvfRADnJzDjFQApuIaREfZrUPxYqqJYGkJ2gzvUjAVn
9NSLbS6ZYdOSMUmzW2YLvy2T6Rm2ZOoKDDGafZal/LryOgMQ2TFkcnthB+EkJyZWVGr54SxfoEL6
4ZM3HclXyFFRu0/X6OtH5reCZsi0RSW1rrEg5djYNRxEYv/fd7MOP02wgELY71f4NCFmFF7M6MQ2
dmN3dwyp1/1s6ExbqjvN9orpHDiPY2RyFQx+wTkRVfgrkEbKUoYjiGS6Vp4RwlgScGA1mlBRK+73
YZnbXA7bHB9CYX5rGNEzqHiBm9BLB3rfevKwbBF6mMVxJsla7DZ/S0D98AS/Ap5hI6S8bqz/qiva
lttjNHZbwrhWLqoMNzL0OU+R5geuKG0P+0jGoogCxK8bbKz8g+wI+y7FYtRS+xwgxoN6NABfjF57
tIdQQeiQiVQCPdQwcJmE6kOHx2uVzhCFKlllDHIvbpSxicMT6jdtwaoy5K3Kffdh4ycltvs0SZkK
0Dl+Gu7H6OwpbEeE4GNGwdiIPo3RbeEdXkAtzUiOmdHf+aThhv+q85cPo1Gsu2wwaeotf4B+QH02
o5QHniTCYxtZGx2EMXXxHKPiBKoKJzONMWEzfXrMDPZAi///AlS550xU81MJONJ1wKbo3hOnu1UB
LyORJQyuPH3iw7i2n7C62cBRBEdqmDExiy1aIe5mOkjeWmcQA8mHYtrbLG4TTToqvMGnmedelXzT
nwtq7BI1wyV1EE8LEVaA2oB9vyMoLzpNOUDjJBZrZqIQAsrcG6H3WdLjfLu3lzBxYo9lfg0Q9qHW
0apR+6pUCe/qncuVpwNFqRu15I2LiTYQbwVdaInjFJqEVzskyWsM6NUoguBS90ne5uI9P5puXYQ+
Xyr2vgA6IJo34wwUAds+ved2fEdA3SMiIAmFcCnmPGW8Scpqqe63vMkWutCi97j/IDBUG7quxCqz
2JA+GyhQVoiIgP5k8GP5dEIcT0+Z6dhg/PcrfHWslx15chrl7LTFO30pi917s4XFpTatyDAN4bz+
vuNGimNSN35fxS/MF93XE9M6X4EM78d4hAfa+MvZcrWEOiwmbe7iyxcWds9HUNcDkz1FrQYXsw3D
bpK2JwQbumxWP9gvmWm6m3+JbQh+vNWtVV6GNRmgI+ID/SFARv35n0wC2wjY7rWiR0p0IKa/OmCE
Z11EEFuNOWoCcQUfkaybV6YbSMsOPyR9YgnkOFApuzTjSj5OcU45P8XR6Vmbe82BZ/cXacECg0wl
U42IjWFqUYd8WkWFPqkWvhcYuqjWQusKIYZWcZsoxLt5VlseYJ6lp309YWVrGeVpmlLCR32/ZgsR
3tDx9xZje094nWNX8YPSivYboTa3j6nIC5x763Q8yglCgQFAwn+bCYUy7b8H0adUpZcH+MGvwTk0
d47pSLzhXgRbe8Lv9LInVKhdxIfQdB2Y1YsimeAxJdc1BB46vCiY7OQBrAf5UsAdF8euvB1yLhSx
n1HD3LS3VFhPkzFv5eoutgV71oZO6XCIyh4slrd4sFoS4HaS7reHOJMc79uGr4ffyCyh2WEDwjmi
F2YVDmzCQTiqP2mKhDaezXQ7OCqRkKYWCUpmnJXFTo7Rt1NG0foZMQq4Gr8fs+I3VUEJgliZwndI
famHMJ3L3PFv2ThqXn+QQVHtqz5yKZvhCN4JwRIa4kBGEsA0hya3nxCNJcQGcsgnU/neMJ44/lGL
P++lXRSQnimepS96xYoHp4xe8BMQAyor/U8lPY9aILR7QDKmXHFhi/yjYDvfCCGQfJ8tI4cwyDHW
Cz0SqZ/3b6EcMHdMM5+pKl+wC8bdJFe/22+tgDxBkEBTzhfpNqgDmyiCqLFDWjfWKcpxa6/CAzn4
06tlJfXwl3bwaeZ3TE5FTMDSSlmeak4en0eY0qVCkfGmN9nAcwNrE/gyZ+hcV6lQCWox20j6DJp4
0PfnjMTZzMLCO3fVaHoYvG5Oq6SE5F8QHfBWf3NaGm0hqq97mqe1ZJFGfwz261pXSVJwF86BGTXg
Ue/kSV4OkwzRmxZf0JRJ7go6pXJzmTBuYf+8pz+nvEaWVenDLBJ2yxskw2fIPe1rBM4IW/p91Vji
8lHrWnZyUWT7+mMeKJClZ1CH/V5d9+SHLqKhF1htNJv2NdezGt8Rfs3iY9Hv6ogkUn0D+I87Qjd0
TSRbGcrOMwbvLHNS/1hFG2FUJpT1dPhBEq3iIOAqCA2mfeKw1XI1Br8u0WTAgqctCQIIqhtLkMUU
Z6mZtWy+z9tev2a+ZWDFWZC1kJOxKWe2TWas3FstxcpPw2CdzrKcnWLnE8ZoQzceN4Ivy/nTUjlW
T/cMvnHSeicjIUPztN6Ty1+70KfzJxsHSY4CtHipAusVttz8MmSHIvuWPQ6/+yqdRX4PqVeoF28L
L74CISnvI+dBuUjtYQH0+BzRqc9ZATq9lunMb3SIt6ea/dERld+CkUJJoPpw2eo8sQx+Ps0uYFqE
wacGYPdmqQYIsbukl7R/tR4STDeSrM/ykQupjbkpVZdWxpOuvin9Th2/tHIx3lc/n8KkGfDjydpY
tqtfG5jSmpwgtfLTm9aURC8NEAgs9+K2DU3V3dSvOzXX4cj9bYnTrp/H1/VbpnYYM3BUWLHdf//U
Kq1ReqA99IjAvnCO+wtChLcn5wmr2qMDMDIBlnrzcKVO4mKTE4UGgTsi3nLt+PLMKCvRzjSIQy5u
lO27FCQ1vaa9XfiHAwPhyP1A6HYC0GJmg5zb1X6PTiF3Qnf5/Pl9j0iap10e/fheFs3AsUx2W83B
O/mI66rgoDyEHjTNyaBIpaG71EniCmJdHdrvtFLQ832RUmeyN4XZ3+75j37yvzRtoSfcscsE0xES
0A6l9L1UXWbr/XIbh3Vh8RpV3mrNPircjeh7dbsnvWhw4xVrYbly/FJ3FH5V3mqa8pfFAkp9oqVJ
xe1JZ310tbpqOA2FoeFxoqupoF2gEZsJj9N5kgzzKc7TgRZ2g4LhhxfMYta4mHOnpbPZw3hS/XP2
LelVeC3AEz9FmHAlvIMT7cdgvJdeepRBeuGbo3eUhCraXunGD2YMDlvafgkDkkQReE7gEc3jfh7a
6IYNefaU8dnNghLQ6pMEV5NDQJjzAhCb+BJZRLgQS665gZ3pxT/X0/kMDkFaYXjjlqipVQEhJFf4
Gq5pH8yDpz9zmju7afumzBIdIq+F3ictdBiMIZoBN+lO8NH6VtuFPG79u+vNstitfO0YdxcPcFVz
f1hJdUQ+Qy1g6OMqlBwsUnDC2RjI2TIVRZgsWEsZlhi2DuUW4mZwWfitg3xPonqpoCdtVA4UvjPn
ozKsA69UiMNhFz1CrHd8pSpQMTtX5f7KyAJEddEZZ3orSeUqnPxjCT/RO8cm6de8a0zPOb8Ru1Dv
ix4dzagEAblR2YFM75lMWV3TJTW9nPA6A6lRVE485KcgHeyaIhm8ArFBoke+4d1IcDxcgLGVhnq+
Ay4Q+7h+xOg9DQd/afrmTaPmOCfesD/V9WVMicPckkCf+ezEDnc42FJAX6WQOPqg+rMHHF/UL6Ou
VTj55g8WWEYbRYCEAJpLbDdOZN3qbdxMe4mJZ0r/83L9/ITzU699Mv7PAWd0AsVYMPEbYyPfvtSg
4imjPXvezYnwUnafkZQESPefyqg/nYGVocogI8UsRvrDw9b8BpRqaaDew/OnUXnCHK330YcWv/og
Vr5X0VQoZvQ1eYvLQQkd010NeKW23x5Yw6oIWZycJGo+33vzjHNNgbVHSy9iL7WL9MGOTJKBymU8
IVuvF7sCuWHKJSPNkNWsrcgOVa1Xc+6MUwldxdtk0SjSvwnJFPTuWgzVRJFRcA69Jb7nNC9s5cwC
HpQFUk7I1otIob/WXOBH+lGjs1zASgMe+Rc7BqGnV/IKhxl3w1xkYIj2os8wchGWFzBmRG09dm2r
VVxH6Ow2yuO1Y2m4nd7Z2IbULyVRwWKV2JXd1VrMtcFvoetloTiKhCGnZ9nmfqINyZtkyzlwfVSy
BoP7SagDZQ6zlGHXBB4kHodVoAGUOnbhZ30iqdgdJ/RkT6DSbW24h42OcjVDOLHxAEphWweWWCqx
uL/tX7kN07zVmeEO7/1zV5X2tGf+1aB/EM8KpRm6fLTmLIpwuNChAsXQLSu5rfmCfBgGWHQLgmYn
GyQY7ofNXfCZf6+DAYRpjy7d1ISvsHSGdHM+tiGvAGPc3iBHqBQHgpjT12UUMm1wGndxA8EdcpSe
Ej3scZfoNVYAZ5grXJA+nqBcpcstovdgGqnIDufeeHJ+Pe1gzd3ki142tnO+2WdkBTslW8K6eupV
jisvVajKrb4/hW5xnY4WgLLsBlXCVbiGo29ffCj2ZCXSC7/7reeaSCug5qjfNjxGfycqUE+MbsF9
+oVDexipeC5NIqsz6sKkH5rFFVIahp3LGBylLXTiyCnt4zkHFxsyS/607KtOQSLKJag3ytQ47Gru
qI+Sd2fzvDjVO5osv7vDvjDd9jtBhKETuor2UzzbBqZAfXttUOaNoDiMA2Y+cIKYEphidp+wz09D
oQujam4fYL1SaVmcgP4K+l8nOI8Cz4MOug1NAYE9jRnt9ApypueWEn8iw6SVQdGgvJj85zjRE5UT
ZSn6jwsIx5oCJplLJ8x+H2H1CS3tfMhwWNvMWGLmVIaftLB+ueUjvJiBD7vspKMkIbYtgN/EK2YV
ibCMr4XdZb73dvicYIJwxEDSWOYr3eXWrQcjeCuZ6GrjNqUk7CwGhe2yPdFrJ49nviVt2j/M++u8
KUa2mM/EBb1KwjemSitoVCAw9cQrtVQHPyNPwXTp1waWAobqFWxid917irDI2d02qIB4SJLoHvaG
H+bPlvxOvNk7ogAnZnySz8w6rDvDSByEMclZVv+2bRAOKfC6xaV6o/a3xpgb8DKkI8SSJc64lLzY
ybRQXOAEohRJxBhK5/gtM+ya1uucv6Gy6lnBGBWHfd5YRfM+VCShXEyR0NUc6t6P2U561vnsKmHs
+w/2l+68xHO3aK/Aa4MJmxZh8bb/+N7VWoLdSyEO6d0gKGjpwRzulWM9dYTjDo9E3sqDe/i59BX8
BweLCKA2WiVgA6KoNLPA5mkWqyq+E+om/Rvd4qoME1WG6w3KgNb4quWf5FHninH8xElJu5FxN/ce
/w1BlycfFjD7LhhZWx1oVgF/iKjrEaszsPkTD/4fpsvBaSgEbmvtQ0+FSe6b+QcPS8B2la9LqO6d
+aecoijkMllIW/b4DZaX3eQsbx5+i0g6rQwtUJDT9h371trhtHCGoba5c78MmuM6jcHuPBQJLqXR
w/TIfsK/gv7hsN5ouJ2xvEJIOkhCaUuDK7M6QAcPgnWjKqlD3oEFW5cX9UXdNrtWgyvi+FPy/5UJ
uQzNLq2B5m6X1SwxiZnMiJrMHVNXPSYNS/eAUqUT7uCRraLriMZ1QTibT7eCoDcihujclv0L5ccD
YfqCO7sUcaDHpuwbj8+b5BCWjROSvSWMA2xIDj/hPgxkhSE3m852Ph5rEh/OaZY5MSaqMI5RhNFk
3WMlOHd9KJNWo3Y6FZ0r0vENqtsIsLEOYK0twyI3S+XwZ+IDG/dOHLSjVHo3f4Ho03xpKYzbz9jd
S0LMSbzGSIkWcI5PQ7AATA56tPPaIPiol6EzhlEOVpk5aYE6g+60dDPSHLoBVIwnlWAo8NeE/B6u
OooZvSYxjWuCC0XQrzkUFq3NaSlgaDOkUH7oj+r2Gz3i7nmpjsdwjM9jWEuOFr73rCqdXnWsoA6h
WLTLUL1sWPmKl6fysuDPynKVnthEL2ghaeCLM9IUAfq9NA0yMstjggzfRClOwcS0Wnd45Qd28W4u
F91F10lvVFKBouzVlfn663K9aA0t7lTNMemV0RujCLCCdXygLbvY+gJOZZCdlkgPl3Y9oyEpXEeH
rUqOpzJZQK9atfU7qEOTCOqPQou6yw3r923z9NcnTVel0F0M2joCCGNBE6qVR3znEOF6Vd5JY5Fb
no3H61OtqZbI61RNWeERrUt7GH7gr9Z0zDFEKO3ETxHjEfsZCF3OuDtBU0R/b8in73W9DasQB7YZ
z55kwEnpeGuAVLn5ouUT4AOlFfyksYIAcz4t8EU+p9eOd/SnOXKSUSLjZTD4VTV5Gr53C/cXsc5g
oOHlpxN3Bnvq1nO1IiSjtPwApiya1CErqBLYkuGKW6ue7LcSr9hfhZPwlicgU9oKA2vRIU6/uofv
jw4Oa/UQglV239Q5CTNK1m5y8HhjcelK6mXseHrHNego5NQDDR08eWcWP7438gAONIPXTh7Kcg0c
RQedflqeExvG8a/pCNmRR5K0Twj8G8YJmWxMnUphWZvOguyAGX7MSmKEeZ4RvpXeyNg6FiOJT1Ng
gFn1TtbE4DLZMR/MORqiNEPmc9zJuhzLYFoPdZFwu2+Ur6LPuUaljMlJmURrp62oh8Svrody7S4a
gN/M+s8Bw8Xm1hXefn4Wx1qnIkyIZsENxJC1lyyxKarFl3wUSFOlflPV9hgrVX0kj0QbHfhHhZEA
6olVkhkckGWyReul6l3ReTdwK4GGhu+RtuW/ChlYK2hbIO6THhtf6jlt074ywuzmtjgodETT8xrM
FX+cpvAQsTTC68CEQsXueKnyd1QCaNf4ghw00ceRF/6ad3/XtmoQijJSIAiMHUn4Bn4JR7erPHEa
4LWyYg3M+OiMVPBilSWTLPbjHaFlUI8qtz6/Xqt7R0hL5GX8hOYHf8qLvod4ZOKKvJQjIZIyWead
OJ1dNsxa52+cvmAT/QM5ml/Z6PuXYk59XidJ+yU4q8fkyIZVr51HbYnHul6d7NJMkvZYpyjXAG9X
1UJHPGz+n+9tRgjundyo3I3Nt/xIdBXXJy5pm1VnLb8n2GjU2f8Yrd7FX+7LoaXWPo7tO9my+ivz
ixtNyD018GztGHG5KzTgfb7CVqhzaeWMwaKZxY6dn+UIwgijOdd/eVqhELD281kRC4y8zD420m3N
8mJg74ZgHXjiTdSiLx+l5nxQl9MyHF49Dgl9UrmL/WC8OPgtVGBuYIsVpjChKX1+DtWy7lvnAjhT
13EDwCTjor+DgPd0r82brEdejzO1fJwpvv+FwoIoXlgDpTN5CAvPvZfBxyodmuAOlQEiDZ9qR94O
DP4iDka3tNE9ZbFJcGp0K0AnR2BWwj3iWmAFOatlmuZ1KaSuMjgHxEntXzUcT9NsxNeRJoPksz1I
2F/IgI2HGpbgeqvpWDADCSAB/QIlkMuYgcDskDCOvzIO0L6/gJvw+/YN7xyHLedUjuxUsIvjk0py
aGJ5yBEScNe82i5sHPxptZfqT/hzWV5hcneAc+wv+svXF5x5yKMonyriM+gDCpQFHYUoukD4oa9e
FxAJQ5gnoxeaVHoqADwPMhRA3Gh9TIu/qxCATNyjYx/uQr76VsHLtaxZvvIrLXLpHCUvwuMu+ppv
t7ZDtswcJfzxlAFFVnik6yzaTASGAQAdcid3HmCFDYdk9cSBN59dv6CZhIHyDcY9Tht6pvOc+Tn/
Qi40/powLnuaVhw9LAtIFEHW4/r2AysNdP0yVBgpnW8xTwptwfPeOxEuglPCRTI8hX48TDUT5/pJ
lIUYz/y0dM5lN9F1vW3eFPyWaPmAMn25O/VR34qHcd/IcGn/RfjwBlj7UPLxSuQEkm7iSJGmXLI6
RgRUXHCI2jxg3Scb+9orNcuId6JxN8VRk5XOhy5G/z7jXeguzEMrlyK7lGIctioq/GNjnbuUxt+B
bvmi3BGZC2bEpMsIWIDAQ2d6Lw97r8bBGmOughNaEWyFcJDj7R1zvfkCDB8tKHw5DeiKck3vRj+T
ED4UP6gWvu8Up/i0/GJ08yu8EQU2ql+WeXkuhujrz8ERrsqpSUDklsF408opTuvlYyVRfvULP2YB
aQEiPwVL3eHgxLkiQFwwa95YB+jcurwPusOh6go6NegnxjLl9/oeme/TzzsJx1RFTGEcYSIAN74j
bZMhr//uZy6MfoTajDRlWYteKiCdGFr5om4UBNQmazgUtjrYIeJZ+c3fehkAic7RxaeFkugm1KrJ
tuf37GQkl+fLbXzUULuozjrcuaYWJ1nJCOSuHYR+1loFcyqMzLTHtjulbPB9/pC1AdleblcmhmAp
SKpcUZLzSoxx1MWEsIN9Tbr1x5Pp9loJH0JHOC9Vfn4k/iSJlxtUrmj7+vNfbmRPD5bHmO4nlbvj
x0h7ISZXkx5FXJPA2QOFvpkGV2KxIMi8apWgHIwRoS6m35XwO3Pt3YDt9a99qxzSzq0qHPzrvOmc
WvCvzExYuxwuoz8V9TzWK3ajoNI4IMBDBsk5ks5Z9j3iHoJ2l9vWN/PJwd3ChqUl0D2C3VZ5qeHx
DGAgR9DQRjTna55xQ1man4/30tgHOAIrkt9Xz7fPkzgzUSSl8OrYOmxs1ncRLAArcDgDbF5sk0wQ
9oPKi7QHsyHjrTnFiBJFSfpsvEE49J+oMzGzstN/UuLDeyzPL1Nplw3XKak6FwqJxP7412LLC8bL
hYW3muxeJb8G4U77S6+Gv00dWJY5yLNZW1ERCLgLL+xWtXr2b9WNdgPlKptFxtHItmsBvqYePQ69
Kvi4tUBiEQ19rKjv1EhtAwniuMcuQ+u33RdeQF1FUswtSsQkPH9t/EIoOmQTJa+CyuH0dYXo/Opo
RGwa36tc8rKnoyD3wBom/+wGgPWOsXWwErYTN3DJN3JpoTfEp31AX5x9PaNOyjJ/1/44dQNXDlOR
oP7x8bwknoSvgbw85hPPesRUCFjp/J6E/Lk/WJe+O9+A2mxOXp9yYDtAeFNjN/9R56E0w83M/eC1
tAynoC2APp+3zlxtcIzJ1iflq1+iWRpGUA/b+gQ+T+8BVoj3/Stc71UzL6ywFzAnlmYlA+MJxEcK
CWVmoDlP39Z/ToiOQx7kVO7XP9IIq1DudTn8JJEz+A1p7f2XvlwMoocklIOoBhTezkW3fZg5jSJA
5CoiTbocFsCTCNy847db5r2i2eAzBkYqLwp5GYxgn2JSqYVBYcNY4gwCWKOlNKysJyfgmiU7iq99
VgSXmqz6qXigF+elik+FaP5S7KXvlWpKl1DT26OqhWtMVsUqWG/v9LDtgDY1g0WZbuRdqtfN2dfv
moxeCBmZ8TKq5+VMUEvuUlFGNyWY9HvxCayTRQNlOa9EHkuFOgb7zQvICfvnoxQXFUwBppjjXpv3
y6NLVu+VGzbbJ26poPa8KTUs6F39h4JDZ+0jDR3G20hZXZUosv30RKW+YWtL3JulTH9XSAsuvKxf
SjLFszLYIK+rNRYs3gzjX9mUGzdW83nmpDBpGsgATEJg889+DsfXm8RaGhWXTXP0OoG5S1tFsGXi
vBtuTdJ5ccaIVLizKNV4iCsZYF+5sQUAgaMc4qmIP4+QfbM8T9Ij+4+8rZfgKmKUdHugqz48BH5/
XpxEDoQhG1cSWna39ttK0RV8Mw5FbIWmUn+eexDiNKNPC/BkyE8WsPLPEusCo8495gGrfmKY+863
GPNyYsD8F9xy55frGfNxAopUBDMUfodBzCjVVMA2lSJReaihe2F7Fa8oyzBJj6nsUYArOQZD8zwS
kx2WP90fd8WpOl+vJrgyMLQfd5k9l0ily8JAcSI7fAPaVkF/FabgHd4nZGeRGSjaAPMKeHI3crXO
+znEAKeYpdyu1K8PC+pe9g9duBNpycHPszuLGIh5Y1J+89MxBgdltX8EVamEczdpPHTbjx+uWQ7M
hTUBeBLLRiPbej23NheE+1K693Sle5l6VPoW7seCoy8E8nFjHcuUihFY2D4qVToHCKDs/hLcwQMa
ohQSvsj/eTZaB8B98oXL2ZFKhIn5SmnNgPFUTFV+OWzH6uG78PeBRCw5vRZksSmrg1nK+cEmi2jF
FXqTgQelnhRlW8BxQMrsngfIIiMUap5Rk/uvmTvjBJCiZSA12G4WN4TfqEK/kmL+71fw4ygrm7Uf
ZCtQayAr4pvUDJbUZQ4qxBe2at0KSt37enZwMXzp9RWU6PzLBHppUAYAHPIEoJPS0AhwTa3lm2E6
0AJU3ch35ySBx9TC5luO+cAjFAwtcy4jwpzQ0+jstmW9QSxMVQBHN6cRDjjyrI5/tiI9o1mBvEJL
49NWsrEFNwCXy+OeCm6lwH/9TU8ReuAJMk7GJ73w9oQ1Bn3etzckKQ5Z5NtMT1i3HmS2AziE6Fma
dJyNZjcc55G/sT+mlijlEPbBqAklElOcRQQQv1Zesr24yfcc4kN0/NiOTvsRcNXgH3oItzfsuipT
bLLkY4JJodgvllfYcSjl2pLVD2LRCnInhJJsLA4fnnVvHQzj9Kx97SqnBPxYECvMmI8cxRvgU9Vq
jkQoUHHb0cyKKg3P8BO9r6g3/B1gYkW8ORawIlE4hr7IwbtHu3pXcePU3SI597kk3RdUT4U+2ACF
ucFqRJrCUGl/1SPMb0j+OsAWWI2ryYn8gNnOfEWEgOrXKYWu5aDL1u0qcjDxWEfZmgNGvybcAEta
pM3vt/WNosPOUmbwFoDn7vn9jz/rScFSxen2I7CWw0eUjpDTpRYVbSXFIFSXnDEtdRTJAeze0Wvq
gbXO920xoSOioQjHH19oHLXoeP1zHJFeN41XLYJci3upRs44TL7UW7rOZdex10YwMXKM+AfgeGme
MkVNu7DiU7Qd3Rnz1ZR9EW/ZXJJiqts2OJktMmDXqG2i7boPRAAsGG5ZuTAbhEwxmSr6eLw9Oh1t
gqVSNLZEr2GaZR2gCwYliPGBHLMmoWhq9JbgLs1TrEmDj+rb0DF5xDvAnWHCXb/poySoFoxS/CDT
L5IfevgEW1az6t++ZyD2APVM6klq8gaBY0lvHXP3oI5rLV4WiySzq6c+5SHYY4qOqDCLM65tRQoJ
O8U6D+7avjWbGNyf89MyEJF9RD0+mKocBOdTbcmx8gwZAxkxITdVkKqnN27CcWr5U2cN1qWJXywl
1lwilvisKyKcA/hcU3wPD7ayJUZ6psfsnpUPCWue7aH7/DDfTXA/UoE1E8hH0h5CdFgxW2tgaEMb
f1X/GCPCnTy9XlgUbr27CbMCS/lIQCHDYFDq9eBQJ4R5ED5azN0mLOHf2zwNtKpCaPQn76IGVc7V
j/1so/za1mwMmzFZSeT5yqOVJQVNZSlT/Q7Kea5h/xTugrrLyFt377eQdt4JIgGOuxf8XOtzZZsL
PJJR2g5KlvThE0iCZuDNTjBTNhTly+N88thYJK5bTjbA9SpE2h5bl/mqAS4TeaHIvwi5X12uDqvJ
wFjFUAsrzem0O0WpANoDwe7/EqXw8bhRyxI8CvqPwPBMKXl8Ys+VSBpI6ciHnRZLeeQ0GpSNL/nt
6R2+l31m5sE/c4iH7lTrwT1StgkcWEySpVCYRze+u67CKIJLXbep69z7ruORJ3Qv21Zped4TUuIS
2wjMFiBkNXTOZds5nI2SenC8diHlGa09UGKh5DXjGIsGFfvRL9RjDhbmpNGPsT3g6RM8M+rKXOn9
I4coq7seJdcGtvocwDqtSNe0xBFIKsIws0qoGp/a1FUfB43/WRMJo62iWmUEl/FQrSowWd8CwaK4
k9a/y7EQHcnZdJW4+z757kwQ16FM+xOLVYxug//gcIzO8zleP9sxuvj7z96TKqgZaDgKFeOCqGgg
g3J3wXH07HPH9HOVgQ8tXiAG0VOvYgZkMEIF7GC0kN8hK03jCNbYKkXKUNjn2RFzdAbNgcWi109/
yWiWJ7ytVXsI4STBRdHYkkrC6+653lhJJcy+Ow51Q6PVu+yH/ynsLLnUyaGTUj1T5d2g846yjWKi
csLCoRLJu3u+Yor3ExRYW2SyWxv2f/eKN0irreSAXTJ5cuEhDUQVFfuWUG0P2A8TdRU5SWBAWi4t
tZrKYVU61JkN24DfafKSoNwcbA7u8Ag20/l5AF04KNxe1Z/736J7PxkvMjVcNsYDNEP4MFzyIJPE
yNzU8N3aGiyJOozkiOFDDBmbFdQH/P6+xVi7j1X8UKoS9JWKJby70ygnuQesviZ/3ksHqc4Bke3/
Bkq7S6d1gWtmJLWe3OELtJzN8A06pKWKivOno5JaVGho6MF+ea9B3vmhj/w5g7HdhfqSumET+eRN
er97D7j2NyTvuSv3d76+EouK/78oLdLJ68Zh7QyR8KMnXU6mkqd0x9EQ2W4QxCixO1z5/tmSeNaq
8oyrQEDzWgtfKrBpyuQ21Gg/x9hpcCbLMvYKjSDrhvpgnE90lc0G1LgjF4b2ISJDIwWRNdfmvRnM
DaYe2B5Ddxnxef4/t5YROlzs/+e8NzM8jyH6ReQhjRwC2gMEHOzLIkAyBOrFrqXNcjvQd2sqd3Se
j1PxkBq+H/gvj8VMefvufmOQnOraStCvP5x7ny2ezBmndkNV9U003TwysgQhrMpYGMpWb/BBV89K
G6fYuF6CCIbdtcXns4w5t2hB9u//5hPoh7GMIPQTJd3RN+7dHUCmH8s6YFsZEAZXCAFJTYCdT5da
qxmCr7LnWj5sD2rq+nyHkJf4Y1ZoJtjggMh50IBEWrlQOzz7dCFP0TLGPBxNnzcDed6AS1BO8V0P
JaOJFZjqhjolgwBFhYvjWoz0iLTu4z57Cn4hqF4g7c3y9UqCDkmYF2+4i6XHXNXp5J9LtaaciUGw
7Imr9Re0i6gJihPSngjtdbRgXqz0L6AO+MFzYWWsOWUs4Ci0AxEja+iA1FlXMHYYj1T+u0vfJk1d
22LJErYEC0ig6CdgqvQlf3trqF1PlH1tsG+ne8JEc2knS7qk2k6IFZpS4sQva+ddL0H9Qlkg4Fbu
UevQtWpbxOkOlLF8Nd3LAijFGtyazMXHG9vGxmSPlE9sHcDNR1kfFOpehWfKL0U4W7TCmSkxF6pa
ZJZR+ZQAL0ZjT7yzxn1rJLmInSvJM0DwDSWTzVQ0JSeu7SCOL2f8sSuKj1vL0+Beb6sKQHWoHEc6
XScf39xN5O6/0aTdo5E98ApXEYPHg1NxArJjdSznKb5I/RAS7bdrWJbVrdeEI0o8alKS8Z/Z/nNs
vW0tI7C0MQUogeiwiUSwH1Wt1u3g77jr55kB8y1afg12L7zAIepEbJUVkgmD9zf3Dklx7UumQV+e
/TgbcJnEOiCHhNMItloWyrLCzZJ2KVb6mvWa284l7sTYFKkmqwcq5k6uOCAW9vRmC6L3MNvNhwQ+
gW+vKLVSXxaCQQSCMvpqw07opp/eazByYDkg0nhxge1ky4ZCXptxkBs7vwYK8X/nBDj0RYM8nqRp
76ZHpEPijuaBurfbd2eG9CIgRzuM5cB1e9OXcUD4KHKyEkpO5EeF8JBGajxBmYP7OY/OWSEY5bAv
LJYjCDRzFe/tnixReexhEGt4/R/RjFyQTpA7VPn/cPtoK3Hg3v95ah178VQ+ypE/aT1xU6116TTX
AXJFoqhboK33vZc8IdKAN0dXg91fC1jNJNp2kL2qm0tzwVrJrTniEMDDehw8FjL1Uo3GvIiBTD7c
HD5AeEujsCS8NnI1hLoPmiuT+n90PMPEGBWMJ6vy6LjDAIEebptIOv4QOxsnRZYfMFLsX2ZzSHS/
3wM7Gd91dhHvlQPdu3vA+Ahclqr11Cs1J6D3b43T5RVYQboU2Rartrvul51NYnXQOLgJWzsNU/o4
omvz32sMo89a5oXONSeQbH0mVnqL8ZnKoKfqPgkd9LRoecv/GSpBBysqs4xS9qwLOaWHTZyvv6a3
w6fwxR/T0ftmaJYdUrh7Dkxl3/j6R3OgsRWBwZS+LIVjlv2bmZAUubSBHWVw0oJyOTOlrr03L35W
2nOW7Hb+mNnOQT9Bz9iOJaSiSywZBalZ5ZO9c2Mw/uwuSwX2PBWhCFgybDiRQMX0IWQF9VGHnUh1
ujawcWrE9BRCIKjrGnYQPooA78XK3zvKhvpTbTnz1fie4eO6kjTwnwbqxigp6V5U+vpawAZcg/NE
fT+utv+TQYbURidxAf8T1TgRjlYCPz5diN56OxoymQB6JfPrtEo7Lpu+e7SSBkgKLxDEpcTRSXi/
rN1VUilhmYUbJi6PE7Q3oC+pHSE1OrGHGhwTAKyQcF0GWEkj0dARwW2QkKurZA/Rhlr16odYfj8Q
e/LXOg9aPWv0sB1enw/uMn2NZfw+w9XJjFyNb2qHpKNKeC4embe9GW5h3V6kuEBz1ZkNyWE1qJst
IgLlFY/uAMsKj1kJ0oedsM0k7qqBkz2GQtOy266jP1sXZeuqEy+XltZYOWqOqCDOSswqUVOq5E+D
w5ODw4Xdt7wlEXmGER3e0qsoZtjZ80WDoccIo7zRfKZ3zkquAoBx3XBlcK7LnSib72sm/y4CFKWm
31dGMH305b4tCCFt0Sx2wlV3xDwgUtHXCP0hfPmrmfv5luOqKFQbVnca/MSvOtsTiFXGnoI5L/pw
AsAomAf3WJiiVVQLECD3xr7L1PeaGnrounD1rPNdb1WTpVRKY+w5gnklF8laqf0jpuc2e/vU+2do
GRPN4QbPpOvHkqI7zseFSvokzxp71J4VmGj2XUU4J8IfNeQdO40PjxqVgG26oLOSoGqWZlIyA3mA
IupP5xxZrxU1hjD+bbU1zHTWObU7Ens4+tbDGm5qVhOyD/n+1Ceas+UJsCWe+7qC21xYiZW9B2MD
xcIH1i4YlxhNgTYhARoFM1U1TUYxWSCmLK5D8eCby6syAjBkjFsxlMR9GBfeF3+1EtCA0GQr4ani
PIGwW4p5pgUzX3GIVTQuwOpUZSVwUqtTBG2EMSUEddBIe9JX+wO9O02QYo5wj5Jyyq4lqdtjnWQj
odqNjxYyJDyZEeZd9EYN0nLhV16Xe4vk30+OekabNaucDoZ+W5AgsPiLNHkIf1JS/EcTZtdo/c8T
gENltBlvIO/eJE6FQlPwPs6EWUcKIdOj6/kMtBjKrQPRqeq3kVoX4q3FRrwHcWCpARLWov1zLrlB
oG+Gg5U8WGwSy/e+HxnrwV/SiZ86o7izqX/MlvpzdEKP+8HKzxpAIWr0STt+AqyG4Kr2IbD5XXJS
fWMu+K8ID9WjU+k/T4SIvx31k1OT1wGZVKiJlPK8nP4gMASo5ft6SqbzFaLMwEEBivyLMYkgDsQy
T6QFbwB9CpAfqW+5ojhd4QsdWK1zGxyNt2dT50rL0s4QjyOkM8PL+NMn1socQBeSuWBNO2/qSaZe
Tx/Thi8WvTK8ofHzzVOX1YlmUegoPA5PM1c9VLQHHK46Nfq/lHttj2Rg1fGJrZ+Uaqu6XezreJr4
BIpBEpJKN98wU9REllCkAufQUE9/+D1VWmCxhPUe5EIKQxzJ2/0Iw8BzraLNy29/GRWkMX1OY+fV
4UqfY/NAUddWooAb8FGLCmct7ogbkXq5zmatl6YJND5IYyiL5SODIR+BHOxGEr+CSL2FG1Tnr30j
hmWJoDuFR93WvIXKLI1ZhXHP4mm525HZaLvMfPYqVq6fzQ8PFXgsRfoSZ6VSeMyC73+Tsjde18IA
7fqQr20pYAywQ9ziqF/zeTSMWjYbI0pMvJkm7CBnFb+38JQoUM/vNLK3XDDkuMCTTfG3Hs3hDu4b
d+TcGnQNb3xsBkWDQv2kEPoLtJaHBET2M/rwgP2S9Aj8tQyC4wbuY+VcHDPE9kNyg5xpGKL0YkoP
OI82nVkvduMzXWLjH05FmeM870sS6auT53KOMyevz70VH5egE6cLR+xZbqE5FKKYE+kmL8nxB+YQ
Wp42GghA1KA2MehxmVeGerEizhzNZzt3FR9SG5T88LoXDdyEYrzVsuW8+tAXV5BAUV9eN5++dGFz
5adZUmH9OZt6DComvJwkpalfbjFoW9WxCRzHuo0ya9TXrHzfQIq0sYNy3duO2ABbMDWQOoZHabMU
UDh2LZinL2aTwRxh9waWrrjW3tyFgmsUajHPH2t4ldr5OaZe2txoE2b6J69Qg67yakrez0DmyPRT
ABvTY96OcaOqZlZXFcOPIROYysmqYgUgSRwlQDIvEAX1tGbd6hIfz87zTpi7TXZgWnQxHd+1ST3/
TC+9wUo94a2SNNPJZMOm1NtiXeevOyDY1ojyC4chHWkxbhQWorKTiRyp41zZLYvuKOVtl0QR0tVf
H66pKZX+ddluRyTcdd+pFAWXkS3EXSPokzv53JmDRnZ+DRLNYzwvycBA+9t+LMEX64lR5uVYWKyi
qPEOLr6xuKuqCQo/c2F+LX3cQBZy7+SCVrPkYNTULdc2E06dpb5MiYh7JMF6JkY/qIjtC1zIAHc7
W0k8zXW/jSdot9gQsHFNVnWrXqB51Gw+b8Km45swNAb9nHwgdcdqJlG3QzDNZJO7lf1Bf/a309U2
Ds2+41uWy5QJ4CHVkvqh9N/t/q3ybdhX+4yC7BL0EGQSj+fG+295gOMRbRnbivWyFD/3CxW8YrxG
Npf/ACrbZd+170zH614g+HjDsQocFSaKoX00Wkz2ay0d7tBXf0XGaxgJbjsIWhi7f5/zyxnkaim8
Iq8m7QHkafNHg6ewP/CPcygk2VmATf42X68oZYXQnpRh0teJakZWGmFK6YHxMKohrVrB9keMtuJ2
ix2fMr3iEc5S/WbPZyhiYfGChZ3ej/nyewYs+hEQj3vWe4vBo8UIyLyXqu5QtrLjB8jg9o/uRb+p
51cW4czeF3p78e+F+i2A5aLMbW6+YvmGQx/fykJH3kZ3q+InLnTuWqvEzsecU6+tLl/6p8o38/Rt
u5a/LFCgX1Qr//gv8/BjhNBT5WOj0mxknbg9AIhMTgsbpp3BLTk20sELoneZNs52QD6JZJxMcSyF
cAjBxNhZTIW4KeGCTFPrArAMSa1WorJEAExB3YR5q31iwZ0bfQ6V/M0kvrljiaFh0LAysErLkugl
V9LSwsT1cob9KRvmn2937mGRS7P/2LIltIf0mkNBYNC+1I+Cf4KEKx14mugp5xUBfTIvPcgap8aB
OyNJi/SZN9Wwa9G3dj2ZaTDwS350w1XjIPPz8UD3nsU607Vf5cFcLBee0jPCxIu+sj+sadcTto4v
pV1rNkEF3D3yexLipW+qj1yxjKmB9LYM7OVSpYv9+oDqh/cZi+YUVGkR5c0dtYvg8R7/lEajFgCy
Wklvvdl6lo9Kxzvmo7rs4tyuF/tZXzp/VYXJ3yQ6XHpx8Qm+v3SFynRy8xjaoMLp4tTA6flFXf5p
1o/jvmozTqERjYA/QGjojWMwZdNisglk/jMF8epGFcValwIKgtZWJCfWAVS1+pajepMAYTh0Fq4q
tLgDPPYNcNY+myFBa6FwSQa24/ES639OKLiYffPgKM/Jzpkwy3mmUXdqk0vHz/LK1e6oKj3zZ9eW
+1eZEbabrvVQ92ZJxkALrb/go0cuOZuFvvjniuQk2u4Q1gnZAy/4ZCVlomSMRtxrFfA6QGlkXK9u
tQh3M+MSWXMPtgRHdQbK2X1OTAJSSQG1lir2WwCrziI5xxb8PK2VsvAHZOK41KYY7+3AT0KYUGij
2nSgKC+QP9NJUGx0WzzmEZssCBWsrZVxpN7LYhNqAlPK+tg1zS1UfwcOZAO1n3zkfxV3BQyWyPn3
YkI16xl1mfCtjPmuSpnwljNsncCgezp1u8DT/0hntExbj09SSEtuIQAJJHy1YErOTYD07oSlAvkm
e5+PG944RH/lm/Us8rsvqAbqiWtD+VR6iZd8zJzuWQYl1mVO2tgFXPoydkwJ92bBr+/j8A3PkW7o
8GdbI0RsBhTqR0ltxEeRRf6Z/5y7+o/dPrI18CI7GTs9v/gZaZsjhW6VVL5+pWG6G1PZ7t39DWYB
mGV1I2ijVP5G2mDbKC4RHlCvkMEF1jdNZa96Srfe6vaa5Hlkjm6wL8jo3gICw6/IhxNLgCbFZlt8
FZqGu1up67Cryl6zCMibYV3rJa+LrbPw2uk5V2nZscdpWe7kAlWHq5U+IL7ICzE4Xv6VNrHM1BAe
xvoBck/7FGvQD3KX7/cxvgVcb026bNXDTuzYq9lU48fYaXQzqagO5LmzEfOk1pqtSVPW87UXFYJU
/Fq0X+mVbTMjPX8hWwKlv6ovqAkk7e9qnSUG3j948PVO64fjqYqlASmExH9TMDBCSglnWieRQn0I
tscPpZFDY5Swcnt2PG6R7WrLdVHErG3mbbgV7au68cQhVnPS8KyVPJXTG8YD0f4i9hnJUxAt4+Kd
RyVYzrXX1+KpQeTuuyAAAFtJt9CVp6G1l5WvQFarStAs3QfkdmKJCGww1tTpPaFbnAAEx1UMsKPG
LdFtPqCbKnrrZAd4HFEdXTp/pjvbxLKFo0EV1Wp7//CEjI8vsa0Bv1mLUBeK28/p5Vmd89SDoU0E
DhzPrInTqZtHm9JSisbOL0fc4SvvgmZ3pdgUWbaGjIChp1Zx6dzSfj4NjEF3EkcspeIl1dRwp1hG
a2Vss2eYpDxp+cD4ieA+IkuoE4e9N0c1fF9tnozerU561PNrAX4YMrolk0CQcwylsoTRDJkVNxwy
pEEKIzwGKW6ecXO2MqNzo9dBvo8NJKEMwTXnhJW1GeP9NZ3I7KSvp9avA8EVaKew1BpMsMSlHGEq
0HMvIp2l4IfUyZT1tB3JhEM+LAfkRAzpw4NjXxdMGLHbC9r5dvrLiD/WyX4VtfIjagdEIxxGcFDq
v3KsqoOskYZ4LWqnDU9A6sEDeWrTpaObuuJWlRg7AtN4hNxzvjzJsKglNvTe24ogDc85COQOqmAZ
STz8GyCP3nSATxTIo6DQQnYIeOPjbRiKUi3+aAKKEj5ayWCw93/exQ0cZ8AsTzHeGuFNBVml11I3
22P+aqxtlkoTkWJNrT2YzZv5qFrz5WlGNIWcBCIvjTSWe9EvyIumOReu4CzhrDKoQ7S9sM3ofibw
DDMnbiPsks6Uej6WLaUiIfuKarNrYEYRc7neqCYjz6f2U8WtSdISEpeXW9gBQ15vi+htOuE2ndOB
cgijeHcjnKI+nxQyR27qzWwjVNkVu+mSGFwTGCpZZXmI2ZJNqOjrWVNo1x+ugugkdo+PJR/D9s8M
7K9aWblbCQiSQTpTbUKJIVLVEcXYxmP5i61x/were9eNIepw6ER7cGQB84hV6tXJfwjjnPbAY+M6
C9oiZhIZeo0vYLFqDawLqseQ5hH9ygStukhdnUMG/CjkqBXcB2vBmDPDoSISCmjGGsLUiaImSawC
FThjCgFZS81Nj93mHRzo73SD8bEhNc3H0TtVuEkWHYOMieKmsCC8JJkXuqGQsnE2YjmKk2SZGrjg
pUzZ9qohimrayCs5iAkU2E0rZq7GnUDVo+1P2DuBIyV4aet8KSjcrQTAJX7PLi0pCLqQMDH3JfIJ
EMJPTsSENLE2Z17S/1jEcjAfewqIDLFrJJy9fFKs61Z1jeAiwDbkFD/VZsZ3ntak9v+r6CyKBvXE
x0AsfKUfXMfeGXS5+eCWct3DM+iKAoIcgvSKC/vAQxdOaK03YFj9qs4ey6ebIqcCJue7ULmxQsxA
edldmiwWWIgeJs8sb5kUQT9qbEdEt9j+fpeev+xZGjHIO6b0OefI28/d3c+ex70TktJtPVDyryeZ
bgl9fpgiumooI1drsqTh8GebXfgpDRssPGPVfGyuH3WRyfjNRvj4PhGI9CtULBDuJOZhb93+p+O6
DZFGW1gH+rHX9M+3mU9KXylPGEzrTVrklaOahaMNNXlY48l6GrOz07dj8x6R3Tyb/1QeAofjXHL8
Tvb6EQpC0GLwCCkx2Fpq5YrJ8FB4znoVpIUqYTIUwtkp7Jo6ynUBOBo2uJDba+XGmyitwPLdjJek
6NX0xYEi8tz3DmDTJj+Lx7bBFmtabLYt/NMBqQhZIf0LdqM1mDB3Th1dPPmuuGdJ93xnvL4+eI8M
9nhkoh6yHjXh33Efj1egmQPn79CC1wdaO1ZXeu0QVlzivLcFcOaASY0bmkcp162rDnO9RhSO4LY3
nNp/J1MMD0qmr0Y91aLxafpLtPmaIFZVDxrJamQ6zjW4fkbikJl3u2c2vpeud9cbza1gYVcgTfZ+
mRj8L6ZPmRcRjbDi+xYyaBb67L5yNeSwKNScpAoOTY+5umwxEBCH6qeETbBATjDTmYtCcDc7mBMw
30rJkU0vauwY+CuI679Yhz9tOwYcUOHgrWjFDaJ5UR6JYgmfTHHTjst4yPj4mR9j8g8EtG8wIew8
NtviAZ6V7vqdtwwr7+8Ty7Nmv7Et/pxo373Q+8BohjO68vWF92Z3D0xuhy474pvbHwYCaX8et4a8
SnTc1QW1tKfDlMORor+4VdKHVrps7YoUq6yorPT75AMdRYKr57pfgdX2K8H+XbMtJYf8NqSbQEsQ
66hG40jnqBADpyUn7t3YtM2FVduzC0wZX7YEunecJ/k06bkqi9Z589Xe3BvLQCn+oY89WZzzoLLp
+2p4nUQ8u57U8GYt3HYH29pgA92wDDdeogDMRQX+RBb3NGBQMlSTRtUB2prrA4n4wH6uNDQf3lII
Gr0lh5dYvp1+jL281KaKPUNIXFP0UZ1Dn1ebZ0NjE+ed1YAqFAgczDNQNdTHjmfLys1UUhG+N/Pk
+1QUELhBs7MKIEFvrETFJfzslpkQ5hTysnX/ryEPIuhx3TfSU9UJFbC3QiK2FTtjDXLUyXUx3rQL
yfxMoprlUxt2qvQQ5+wbxSnDKbM71G6ArKadxJCWbG3JPLjBNAeG13fKwgd66Z8Ov+d5LDvCSw/1
ATVoHxGABIDf6OEEXNb8zVLvePL6PKRE5W4+AEfgV/dVn7hyyYYJRgMnULAA5MC/bU56tPJR0WY8
fXrAoler6S2ysg8A+LYeAYAMjRB/IsslkvZdo2P1QYi2Q6nMHAOjDD4ksENGDG2Dh0dyPx24jHHE
13B2DUuu1mCMVN7RJGIyH+hRCRv161PUhQGhWfqNKBAAwxYdbOawbGTRiXi3lIZjS5KeHOiHOAc+
DZa6HKwPdRmzkc8wRin7ascx8eyq0sFUuurmzyTw/k/zTBncx9JvxnQWHsWfr16Ho8RWcGGqTFg0
R1kW+rLzmIZ+l/HeJaHJ0Or9l2Ic8/dOMl/gax/OmOqc9xisj4ziKLjFL67wiTodKxnJyqVhzGro
Kour54uB+8BQ02qRMk0H8Gk6QyfQ8ORtyM+PFH/2DKx+pIILHxA1pwpXaCJs3GohxrQgDhkOe8Bm
GyL7JVY8UIsaGxLgl6Q2yrIlVO6WQ6HsagFloDqwPVYHtNs06x8AKMq2r/PLwzsCKp9/dSjJ/BkN
EZeO/eMzyEV05fDF0hi+viLrfsQNpXAEEXZSs/qZaxLPe7RmyPlS9WbnXiYsCmWbClBsUQus0a8j
AuEsYDeUdDccXaOW2WToEzNaBlgIx6AOvom+Ih5cMcr6ukCqaeBFBMfAsXFPEjmQZC0Bp1tIU2uJ
/RPMXbNPl9qfKPuZe5NAwRUmpmbXA99IuiPL6cudi0moQ9kybJHFIa0Wzll1LLVe55PQCcnA507u
kCDy25go4jnW/gMlBh7ShOGTO2eXGpZc0e12NrIxeBQdO0JrC+zfIXo0WM12gVoz3+f3i1UJuur9
47gbewrHSxTvb47MBDkE/rYlkRo+FDuI/dBEWU7mvqDdXNrSiyTDZpmBsnM3Pc4WMPvbcGR5Lwe5
CxA/UVgw9BN1T98v9e9r0UyveGlTXkjtMfN+a+hhHqSKqRyaBoHnvoVa2MH1L+GwG3Loo5qutQ2q
XUHeVGKttAeOelWfRMC+BfN2ESSC3mHnQwP7Bya9TRLZhqtx0JwJvD4CtitdlQL5zwbMvLyefSM7
T9jfdmP+26bTFKJI9LZLflS2pmV22RxSUnauCl8msmHmpqmHsYiz3O2hoVwLMemDSI34wAq2xM8P
n6yykwJdxjV1EW90/HDfABIBhJ23oql4KlgWAr/ZyN9bGNVgG2oMkroFNI8NOnMgIjZTlkxI8FYw
nZYEqFEoaTVYZ3p6qV9gOZyYuVF6LPFeHGw/XTg0zT2nex25Vf4hZIdduob4T9NmPGy2G+rd01xh
BgvxqXAYV3A2N4s5LsfZX9cPuVykp0XyonaJaIcRCQ+f70ufdWblI30rjQeZyQir34yGZMICI/tj
5o1SRBefxzDofNNm15NKCs1hYln2WlGMlwqgz5kQpvHlRRepgwRgXx0g9BexI9daCA30DbeFG9wu
zIbRa8/cVecClGEiIOxtgZrQeqvMyJyMacCsFJZmGXh8u8vsfxaaRxGvLPt/4eH3n1kCth4BqpqK
CqW9li6WD2eM4TQl1f94zft4EW2HqQdyQTWPf+3SXZdzREaaSNeqQlweU+ub9KTpAXJ7VzweAaqS
mvdFjmvhNbybA96sYbJW4a7aorwALmzfShc4lsRHFcSGXmrgRh2OuHmJUhbpYRppgThDytdpPwAc
+6uGxuKub9u+SeFpLIP4/XScbWwZHXUN1LgwiA2H9ntboSn6pWWyFxM/r/jcApawJrl0II2wqnwV
dratUs17JTw1K6qk/1jHn0SfIoqqXFEBNIVWKf7MxR3QVwyEdkdLusmk3nlpp6VACXXZ9V4y6U6Y
Se93AVB+I0ok3OVlZWQtbayBuMB+Jm50sPqiKKm/seRWQPMeE9Np31mJhZORkOl8NVdqjgxpBeYT
AWKfoPJUb4zfyfzKu1WLLjtTqrIWFvrDpaXv9bQJhFN/NhkwCJka/BpzE4IMMdaRVY5JLxlIrp+3
YNtqDhQHyVEu5PO2vacB6k8TJPXytzSa8uT8c5m6th8Ehglw3AFa871sdTYK7vHNODRwDqqZBDWH
zbGM+5hDnrSMetvVRzTigBUsO921qm03xA5HLKx/Y3nFl5i/mFQgGxjWRUqFb8jFPjW1j+MX/89S
mUnhNGTgWYSqye9Iak+143GAmpA4cxfey0OlK5BWds/UyAFySmyY0xK+ApoJTVbdlu0RdF4BjAwq
DGMf5cNUeCA4K/TkFU1oSSjkMzMgQ52FawBi7vu4pCh5mt8ZkXGccoEfDb3CcWkD+eZTe7+itYzD
+qUXGDa4DWhKd1mi5zmVlTbNqm/ZF7qQCMZFj7KKaa6vKgJwJzhUAR4Rf7VI4IOoPxvZCn3xJ/Dc
nXXl7NZqq1XLa0afMU3y6kMwhT2C+ktVZD/vfVg6EOwI5oda40bh3dswRLy9qbQA7YnMZpv37KZd
7hJW6ZIGxCcIx8ofnaW8asdq1jV4tQcbXNopFIiodgQS+E6HYhHWK5Sv+OUJijpY99KRd7vVf86Q
5jgbWvO6GWhzUhacM4m4dfN66h6EczRN5uKEU6IC/Qgzaw9QU6OJgvIIiES0lEKVtXXZsIwXor7V
HVFluZUGJ5b7jl2KhfO5xU44dk3Pv3c5BbEYqSAUzTOhJKwyqzi3so5K7HUqjB5ncaKkTSIn1oWg
6t/p2DqW74STJTURSN6GAnIOQuthnmCjp0d0OYVUo1r3vWphTe/1RLqPGRHqanTdNed0+19KKDmA
nLJ/E4pjItfJ0brICVQ9ttEBCvNk++HDhFTn+wNJQnTfMurqrZypx9ki/6Lj6hHhSxC25oItpqPQ
Z8Wozg5ca70btvgdkRaKJlbDk5KboJinSgBQbRgkXSoqoDj19L2rPVTT8NrMj3Ul8Nr9JhrWzJpM
WmVA7DNfgdizihwUPU4PJPjyUk2GcpckUuG+ymSlixrK0DW5agJoPfPx/Mo0jf+dkyan6hwjtjlZ
ojMwOy0tVZn8sk4b+vo1nbuleqyff5AnkiNDCpgT5U4aq8brX0QuAbfqm9+KjwSMKxpSeOzoiaqG
/Zr9ApbChB85fEF/o19/GYm7ykMQzWTojk5Lgbg7HmapTkABKOzX3fylHEvrmmnhMC1+Fr7vEZQn
J8BtxOQQpPRUy6W1hiXcErnTFBu9REt+x5n+bBCaywUTWPcTo2VxIO4jul2vmts5ZDPY7PvKh9Pd
916yovFmP1NdcmQCXP7/z3v5SbhBMFKkftgT9oE/MfBEBou6wj8SIfJlT2+U1O1oZUaDffSybeha
UwKvig9jrvNDIYjekw0gR98JVJch9m0YwOoKpeWbFPUNMfHthqNXlRA1D7DRydJm0hHFWzQNUcoV
J5edF16hr9XRwTFmwpfQ9OSsy3wHk/o6GbS1J93FhKsT6ik6J/NASynUbSilB3d5Xmq2kOPz2dMd
Uoy3mkT0z8TQ9IOvLN5cVK7DyJsiFhjTi/adP8BoSU/nF2S7a6XTOjQ7wapRLhldRnGEJ7oCP1Ul
xLCxsjSzgJAMatpii+IMNJ4p/SfoGygN7d6fQ4jvoC6bQOZ7ZRPUtry9ixFhStuwSs7B/wIorueT
14jUW4GQkdx81IlbGAEjsPlt6GtgD9qaWIQ6yk0RLtmanR0HyRvc9lJzyJ2+Ma4Y/L+j4fbkZEHB
tHMORp7scRxlvfnRknPpPw221QQ8D1EelttS6GwoGaEKyRRT+fNlSP743ZW+P78Hh/QIHwLgOcK6
0x/FhGglh6Nz8QdPSkLUGzWsN2AcMm4c/OUx3acFEmDrBHeWw5SzrU+mTmya3OqZT3wfYuHvtJnQ
LOLdQZuo2+FHXW8AhE4OQyqfqx6YIx/1LoEL4vJOWdA2Cev9Chr5h/H+deBJY3uc3NUeIS5n3iYz
J7Zmbrec3nZdcbCIfPQXnUEZIibxU/gzWmwPybnYjBb250E1BR1SKyByRNq0VdWTbQziibuv5mVO
Y9jilXrr4GH2yirR1sNTHsNsdGhabxPVucLv+5xiY8H7yhQitxCN7HJ/UxXAs8umNxN/zuOyvtSP
JeXaTBFjJmFJ6DCJ3E+nJ6yYEjN9+B8nqzzfKkEu1WMf7ZwOhATPkGhr7+zOsXCDcrzMHnSL4Uo1
td/yfdpS4sC5aNbHS86cxmc8uV8KQ35xjLFoq07lB4T6MGiHguKZBKx39lmt59McYiIkIODyJBgC
b2QzIuyth1Cu07sYLPiNAsTKB6Z1Ucbmjs2KSDwiOxp340T0rYqYmDHUkcs/TV4VBYIGGR6qck0u
0dxOpsTrdHM9TlIkUZAjV6fwR1eOJP59QEz3hl7kGtJ5hk1rLNOMWM+PR79Ht1ny5T0Ka56m2x59
as6WpF/5uLD04DoL23vEEWd4NFB2zGfTa8R2h4rN89ghwirSEcPXt8y3FBBgrxM/KsIGcqHkggXS
1H3W92YDol2lFneFOPCv0FwcgRE6EidJtKnClrCte1jRrkC/rVBsug+n7SEsuMWQblzQewhfEhwf
8EtGqDiUZJzhm7/jOPPqac8D5oY6ybn0SzLMVELhTd5lUL0injUzudRScZ6uaCvWml4XmGT4EPbw
wm0J7sMGpSqr1Ia2MGRQyfVeNxUXFwX/Jd8CnCQHDMmvrWktb8Pro4kIZWPvrtf9bVKM1dF/RL/x
tw5FTf6C9oY2CuwMURORbHRrBKWgRe9SWHsDiqqDSmaxniPd9dcZUNdxyd+xBAtV3OZIG4iPFuGr
UqLRfmL6NZJje+1Y7cyTUnj7mp/5MxQP0BwAVeQNl6V18spNYWm0HsEmI01QizLRR7ShO5wIIrjp
y7cFdvKu7Lde527dzLjxCkc1DBWm0cY+9ImMizeKrwu5FCdkVSjffDZJyzqh0f6IRuz4YwtlE0it
rOvu+eQBGyLL2/saAmGKghpCQ2d8E4TAIvQHmmQaeigLbXbf3ES2U/4Bu2ecCDnKt+3AnVhq2/Ey
jAuK2XQgC0YTATYNTafJdvTx6fJ/YcevgPlJ3CEnBQ9HtE7q3xwNpcraB6407EjM+OjSwZ4x0SBT
BBqyb6n8Y2tQPuSiT17yLMYAjptFMPyP7b44dbcieOxtvFgtglIpQBFTNOupV4z3v0cR/EazdU02
Yaikx43ZmL3Caj0fBrMCaY3fjmub4Tp6zcn3O5CnuzDxkzoLmjSG7wHXn/QI3sbHcWiRv4a6pycf
TmwAOfuteiwU/dTtiie+8GN7cSQOdsLNNSP/RINuHR4AuCefsHIJsEqPTAURbqzH4Pzr7WIW9cC2
tJfWNEEbA/WJN6tiYyRq8WTtMXDCIiIL8gcPGToz3v0ztIYqdlJe/+w//bVoyGk8SlcW3bzB6oS4
sNxmSnk4CDBMojkpjzhCit2PkywRFLS5wXzX/CXEdZoE1IG75vub32CPIK0Qi3Gkms4EIsLeu57F
sy56ZxkuIpt8kgsOMLz5OdRJLqubdqizNsS6hRQfNsvvgwP83VBP5EE4K5/hKTW9ON7687K7iZuK
32ZUbo5IGDxsn/ysEQxiT9/oOOCADqI/oncCok81aM6ko0Bdkh1ZwtTUa0Kmtji+qkhirPIDiHDz
D2dwDaT36CDk0uSl/CNVyhTG/MftJAdi3c6YcKPO+bYZDxyGyFPmld9/q1xW3KasYEUbzOzx/t7r
I9mDKe6W+yctBkPwNvRQISDmBh4vGMQaio9Gg9LfiFMCgVjOjLNlucp9STRbpjf0aPKX7lOVcp0v
ZnO0BgW95n+2xPxjMuASBPAFEXwSPntVGrZRCK6D2MdnK5edmEJH5TACCXNR/DkApzv4/OaDnUb2
mSv5FxMbVGhyh5GuQCRAwyMaI9cwkJ+Z5WFkhu6ao9QHtNJVv2SbhKhi55jwSMVVOkfyU/mopL1G
gl6Lk5yL+S4/XWXvNx0y7jcLjf1Zpd3aqY6ewHH8L2fSlDTPJ5S3Mgyac+6B9FEbQu3TyZt6r6Z1
J/3ZzgGbvh6T0oknug+NsvRsX7URGSr9mzFMiH+pDZYsWtRouyJfhpL9KWCKy7fLgMW32LQufKUX
0d1DIfDu78wqkW2DaJQeVjQMUgl3jhyxOl9Mc3wMXvVd0WhcYCs/Gvxx41sySTsCIsQTuY2YTbd0
EPYoelfmz8wu/vFLFHlX3AJD0qvMuHSjicEvI8W/KNIS73D2pu7+vGm4nHLUwHoHorN8NJg2WQIF
E63gc4Qf3t8ivXNQGzJRDDDw/ZqicjoFa5qsfNOOIscuXv7fjF8XYirtjLERt3Og1e00zXBrEmzu
BogppUuQH8enFfgHv/PXLLlBpKX7/vq4CpdniovwQ5W3gwn14oGPQ56hWI3QdKFXaoBQ44fqtGRe
euWlJ5T7m3Az4x3ZpDt/Cl3do0mIy4d6x2pB/7ShZ6zt4RWchHmNCsEHyb6qFLreEbXwJ1GLIwYG
bujM8CMgiVtCErxg0IIiXXlVGCgKQ6U0uBXz2LZA9IYfM5Yco1S2jsAEw3rlJTX9a/RraAKpeH0A
FHNzZbnbDIMizhRHMZRte66y58wbZQK4R2E/zYgTL8CTWZAi0FwvrLaro0vVg4PBeyq9KRKn4OAv
L9Mnp8W30rFxBGOHe7YrVe1tHntZFsSfze2HNnjs4KPxfiMmvTvv9A2FUB80Zj8Bo/JetPd6Wzau
YyW3ydIr71+LSSpKFlF0DdPiZWz5tJrPCi2pIdZWSVQd1ZLiDA47N3/TAvbNR5AJCPAaR/qYc5Ty
qq7P4NMa2E8Lbi0JHj9Ye5zPQ4jzSuqtom3caHm+p6tn+dVUFwMT3UBRJpxmdlDx4YY++rGGC9kc
btn9jTYmC24RnJOgE+b7iWKZNdUrcNeBaC1CZvTpZ+zo02bKxzFdm5HRGawaExJ89AWgGlvzMFmt
ocxnfwHvgxqYnI8aHJBMhnaLMu1NQtm3q3hZ8EEmXXRsZMzSZnt9lav53jvytMaAYX6NlrPVQZdy
pB0GedZqzBbz5w3hvW0Cy0ZqYicFLEPxwsQzvm9y+2NSUaRCd8rMVRnyoG+D2I3uyDH3y3XmADb5
DNWxGI7MG4cbJU8wxJ9DkutQvJfRoQgoItjIQj/Hvdewrdw5IchWVLwwMxn3zERDRQa2OL+qSafE
GPvzTFX3VIIUQrtSiJoX+9lZjVAyi9+/DegVhRdvTNSjxT0r1z8VUqGfFJwePYwCBm6UCD/CqDLw
tmbDI6QoIyKflzAubC4fRNzGgFs9MBU9MaiKgWjdM5HBqtT8ZoYkWckCf3JtGkC016JpaXZm25Hm
2TJJRzv90GvG5W8eIj7q2oOL6YG6mqPWjro+ubQHDv0dPiE2SGJnAYDURXYA413te/PrZwM9w4e6
bi+F6ReXRRRPK+gNNbDwi/wF3WQg2r5ml93TDIVG84ayK6ZZiAsyva2pMVTsi25LbdnnF+L7aTda
W/Qa829vrLQ/Ec9jh7L5aJLp0SeCRYR6V8AjncalLAAJfqlA5BmiwFXCJB03sMY+B6mBvYVp7U7Z
uwMpU4n/e4dQKDGvEP9J7oWDwx8+PXmJGOrKs0+ta2KYuZ+H5OW9UgPQqBawqrEIHoproTkPqpn1
MUijpIrFhbEvk1thA9uP5m9wVRZ0zzDetrgi9ht9ln+p3h9M+tk/on0zDX8fSpAATBAHen73+lMS
VeO09WGEMA+GWk3Hh5o6iLDsBEGT7E845x68tXdp+OUN0mnUvWjtSzEgblGQg0fao/VK6AQZUdGB
D7HjP5u7MnksZPT5AlbkcsY3M3Ap8/MTqcVMGBIZRpzi49ktITf3DdU3YQ2HNAduWe/tj9ROxcZ2
T+l0kLklOohO3N1ttkURe+U49b9WxO7Uj8iBffgxa4TOv8UzkWC66c+vQMkWOzjfBCb+vT9Iuc1w
9szHOKy8UExtiP9dB4BcqjE3aoFVZ1ww2/iBD36iCWGVXpJLwdsJNd4niaIyNXh5bBO67bMDSsy9
dtdrhTwOgUvJgvPJsItGn5KJLho/FIYrCaOBUPMzS4ow+xpo8ULVGYZ34rXW03frrAal2RQENQDY
tKSjpXNo/QIKXbZotJs/EuIyQNOfS9p5zCo9kcfVsGQEiSdscmvhc1/Nv3PRO8QE3G3qAVZ93Lvd
StrFlgD6HbTg4ZZ5Ky3ZcFZI/oHTGGlvqRTfvPs1eqKiCgQyvTFcGlNr9JH3sty5JGATzppyq2a2
CWEayix3Bm/wMZhFOeJhN7YUUbhHjcXBdG8VwfSCtFbutC2MzOGajS5lXQdUpwW+hPFC4Z6hCrJb
bde0t7J+y+saylsIGpI6jCdRzEvB3Fm4SnKWalr6xlAXpLM0/ZXVR9Ew6ZEYSAppvRIK2TZCQoMR
4bWIYvHQ/2CmVXx/hfydScwkPM0ce7WAHyRSkHDxtDSS4oJx2G/n04GKbsu4/aAIE5SV+Nu6oc99
fixyo0huOoVgn1SHIJnFR+EunB2GbKzHp4ZzfZIhPSPlcp8WBwALepaVjSMl1MeinUoiokUOt7OZ
E8KrLJPtCUWJ7fq40YGpUsZ6UwaLU/rppycUuJWrfqDMOhnMwbItM1zi0JIqXtJj7fS4swBfSRL9
drvd3o/8Qvty3gm9VrkeiyFp/DAEi03+XxxucWPf7NyxuzNin8GTRrQ384L4mhpljUJKAg4xIDnS
fAsJRqUaEV/iVIK+i4h5JhLnu0g4ZgARCbhUToJIMqIoiF51YGhaGJ9p5/EJVVnIJvi1WeK2kuKS
GI0C1l1IkkRK/CzvG2FU7HgLCE8zuoqoA6kgAH29NzG/oRF/Hv/jeBnbR9uWStaNtwjQTNI20jLy
Xa3k8FcsXDcBj/IHKJNZvZOik3OEErD5CnoLsUScLJEGkZDk9fhZOBW0zJnCeZFL7Im+dwImynM/
f/i0ctDQ9v93D7QMgQx4bbnUHY22SRoqVvtyCOCg21uVIMwo5G0KuS9n84hHIzjvIqJX3PbScAHl
JokohK3JzyGeia1FiC8tOT3wG+7DPkcrTCPwWg9f1RJyqHPOm/ZA85v6xm+fZNfoBOjiaNCM4HUb
agYtdQ4dLU55w3khOLwXyX/8bmGMqnskYH/y/GjDGowI5WcjLD1Aupx6/hoxIvjJuCY1lDCTk8ya
QfU6NgA7leQ24w+BrwWsvhqDyLcUZi1jLuOWXBgrscjn/otgpKkEsWQ2tf8DbjgOJHSY6nuzcsZ+
WZ7xJ9iCTW9KvNMBr0kAVg8EC4Z/IlB+cg7KUK/gfF0BQnA0n9TJFjQFdVzlBvif0NT8ciQvTJYd
ErXBslDjt/9rvmQoYpb34815zBvIo3ttMb79FPHTVWC9L2fWk3XqQcoiWu0WJi0XJNSIv0qhEbZT
LB10ROaqpzC2XWAUpClC3M9mMNrD3V8waeAvBV0CJWZFA7dB9zr9X1Q18v12UvsLASC3s4G3mHVH
Py1rbh7zTvAIAI+431BDBn6Mx255wE0hpRPlb/dYIwgIuKxLgFAkQm5PHQQnZmoiFihZZiOI8DCp
TTXZ5HsPk+i8msp9U3ueszEcR4onoH8VDxPPh4Vje3r1i8D7KzZQROG8Pvrg09uUMLP8BUpu7PX5
NVfSoYrzvvQvBX3/Mj9oSnb8pIELsl8z7RnHj/x+kJ8KbJsZbCyWvc9fOzET2ckC68bmyLpmmpmE
YFUmS74yN6Mp90tble0h6oLphMsiVY7Suha5SwuVcJc+rQqM6os0s9LrAtiqGs3esZil/IlVSlsQ
MVrES+LVg0vJLMF+/VQezpQOvWebrHETusul99lCkaQ5HCDN0Y7uw1uB3DYX9Cw0oF7ccw0BISfm
LDRmVb+/Uq8hi+zFnPsKoM8i4g+kFAUrd5QBPRfU0sFCBAJ8MLBUiWQq25+/OQyFu74b7V5E2y6K
B2RiidCWlZ6P0kmBBwbOM7LcgSXA/WcyahJnMPkoGsFXwSAPuYfpYur9k34dn2SI5ZTQ1mW8FCiB
/L/yAreV7lLNMIH8i75QI+BfDf/J4qJh78smZAd7Dei5k1o4qftT0x4nLhGSqUWpLPIuNO2vLvgR
If36CsOpByufm9CFcHh8aXDJ3kLC9AnZbhkAcmqEEwEciAGwwqyyMWhYv+PYHOXbzjm7RAp8yxRW
U9qy0nKqPdABja+Lzq8afKuEAbFNV3csHEYpmdpZd7ev58OJbH/Y9MbUCghhs+B7vd91J6t2ue0g
1LZvx4qAUHjdniCZ3VupajYgr89rhgO8OvwFN6Hzu0GwRTUA10QUh6uoBhDx/8b/8c6P+dGbJ4Xa
kQm6Zge1XWzw4nVCtWN4ej/KHRtEn1e5B2uB6EecKjUdGXE58R/ZypOmYrssjGe5/Dwmgwsx5gPm
Z+Whv2WW0doUx1RsGPYDW7HTJZKTESRQqKNFrFivgWhrDFy/kAuz7EqPKwcYy5n/2FYG71UySAyT
LbQn5Za4LESLABJNIwqWlozJhuV5oGaqNm/IF96qZfDU9K6nYPVHW+JfneFXjM63FbSziYl5s4an
sDBNBdO6EvoueQY9hyC7NGK9iAUYWNsKuybXuYuiU6PBjeEI92Of7hQyVXMMCGJRNRnCb/VpqB/l
dMbfHfvV7H4qR/zxcc050o/yjCPfEslG8hY7DKZnSkZMGSWss6yk10uGiBKvKlXnl9TUimML9JoM
xLB2BuqIWSH0570IiISvfoUpopJBqB7cqTDOGlLqRllX0CRrAzYxrUwGsYZ9oe9NI1n36GVs68He
inc+MV9tpzXKho4Ft6cMXrKvtaFYVuXlQn/uI92Wj4LRTe3nRu2ySqaW9Zco764Whp9TKZ0SzuTv
ltIs4tkr/NF9VKFup187lCvlp0Kd3q+UvTS50yRCMEy1RBs4RH84OY6hrRYmvxnIzxJhnqC5o+bd
51beDidzIEy4rXb5z+/tnCeh6Me+/LtTulhpByw4jgQiTM4hu8MT5tSldgugjaYR4TUoSVXS/hli
lZVMIvSiJ1ktkBx+pzAVYMD6uVpIQcMW3MHFg8EMEFKaQah6sh0Z8vrQC7XfVXF8BDsleakLUBxp
ls3ReKPfEArS7hDdK/SqKnENk0FYc3Fvp3gbP676Cj/HC7uX5LR5djjRqMr2ZETrlUMFMfdSKXGi
71Ynp6JmaFcT27RGFcfpv/nmC/+wDLShPvDVivt+CyCKLFcaZbF69zJ09QZwEsh+BDglCfOhfK0d
4bp81tsQ01h1gYd2W7rjb3loY0MArpHCVfaf/zGjs3CU/1RQAyPupw+Qje2xm8mJfHMLwU3S8FPA
3jJkpK3MyLePiJvMRlIj+qyedvmqVSGWNmrML/AsAN5dC1cuDnHbh1Tc+EmIprG0MqhhnGEO3C6m
vrYNCapKwv77u50IMBRMh43IReNzBSH7tXUxCjyU2FPgMETYD7t96B33LOARcSAe72EdSz3egVUb
7RsM3ZwGgau1I0rTEgB5B89Eqa7SgLOOEuqMI/MVlrPV2gnqZMVw5U3CuL2g1wlIotLQxAD16RWW
dzsdquqH/R/iwpCplBJT6lnKCA5Uu8EKOHgs1bdocgMI9trFKrqIVFnBNAa/n3efqfgNlcnJA0Lr
8KvIUbvTuLIJiXWI/uip21TJ+u40Ii60znuVUekzrOmBMf5DHr+FLjARJ3TmfHDIW69Ni49Mo88g
yk7DIuoK9PlLWPh/NGNBQUyi77Up+QTyNilHrrNWYaFkq+j2Rzx6+oazKctWT5/6GobRRCU7D3st
YfIVR4ZmCLIKXq0CjzcC+jZ+22TBK2M42jvE6MHB7lcEsYNq1UPpA5i2CZZRNv/RJAx2Psnt3uqR
9m1wVt0KcaMKd8OumEPL9TqvqL0D8o6TmVNYMqq7l9RpEDkxghAl3OR8Q6m6jtlQcPOJ2driESNU
ZnfKbe/UMMJ4pBScP5VmHmn7CKqgBbpNNWft3dQD9KKaLCLG/8VPBjdgngwWa9EJSpsEuM4cPyge
QWyMs+JArelag0JF3mhebOhJOKDq6xlw0c1bxMt+OMAzsZLpmumQmKqNm23FEelWPCSx0UuxgplM
xC0QydrZE/yNxvzAKcWQubrvKO95Tf7endm1GIHFW9ja8ZkNoTk4BjyeG2ShTESX1WeM1UXrrxes
7pwFNkkal3lkE9iSP5uYujIdeyNzvktBkAlIT3VZ0DAI+Tp1FmTGaMs1Bknqmf8T4DW1icZQCaxx
0T+xziN0K+p+F+dT5yf0HgScW1S0gHvsJCs6RA9yqBN3PKuln9E29fkNgO4Jb7MEfgSeIQcmjHUI
A4cptTKXMYkoLoCWPACi46QNaJZd6AV9BmGQKWYpjndh7MOp8YyDiBS8EvFRIfLeVQ9YxQcBXUtM
i/P7UbUAEm8eD06sTGL0eM43T7l09i6uX+qNFL7u3ss05L0ch4nasb8IxivGnWNjxCirE7G9ISmE
ybR+r2zhSnFDLa5utRD4R53hLcS39nFHUwbvoErMrcAzASQ1DYPichQ5eFp9HpGTIoz3EPfetlJk
aqQQZyXKk8hRkbJGgiX6V2AmddxMGtEDIn8aEEbZ7+GhGOVcJMLSXxusztyXYwtYnHaBSYlE6ETE
JJ8HwPpR2f/4ygPCYBeEqZIukAa3RU/Htj85GQ9taApj1B/SXfH1oRZ6yEWLNwX16daP6Vn9CuAr
253jRSNyYsOTkLyQ2/VV6DXBv7cOXnvvE82159I3CQAZrKCFxVlegflvJJODp0hlcBg9sjyIJ5nK
fN7W9JyrZS4iFLiizotG+Lt1x//oh+Kv0+cHPHGCan2riWahyzDFVoGzRe/Lf1harmyY+3N/9o79
EU2/mRaYWCUXcHGUHJ37zYhIKGwY7HWA9C3OBPOnlWOE5yRlRcKp02RsYhEP1IjcY3RxhrOIu9FB
BSfTMKFxpl5HTM4SZfnjFY18HtsLUfQHSIU2tONOSwdkeUDlLUSXf4rAudZU2deSIDNU8aHWH1x4
A6FLUMC7/Ow8tjbh8z1JkT0dYtkHknS8JX342ySaVXGNIpORIAsAwtwbNBBi1svtLX9E2w+/MrVr
vWBxppm8i3241q/8725yAN9pFTHUIXhVsJSu4+8ykSindxM1bDRKk9U78TMD05pb+OBAtE1+Ap1e
oZKKLHluFU80gOVXpq6qkL+o1BrcXJyGaD+xrvmSertqlYRG4jn7zEEXF7n8Q8uJy0jGlJd1rwdp
S0xV1WnQbvhyGtP+qy5oouSNsOq7I9PFwx//D38GMZ3k2IrZTz3nY2dunbTPaE8gPFOa1RX64p+X
aNhIJ8lBToid9QlaYZN5Xz8HHBxEZdEj9mikMHgVlWLY/skiXEtH5Z5+FwEYEwohjtuq/x8n17Go
OJLQBVCtAdUCcyZXXRto3/k1E3GhqjncuB9Jo582ZRLJH1gERrtoisZZQgiFDy/r7mH5KYJol7Fn
RR3Wj/HK3LL8OL8L1oI8x5yobGhmF95fR0L12SvYK8wmA+wkRxEIGcAfOU4W1ijciCd3/QjPLvWG
VlD5JO69ET3F/hC217+whq+BpJ6f1h7jceWm/GpIqpYNgGKphaYtN8h16XtS8trMne4pdnRbp2Z0
FftxR2gc0+rAHze02WZgCCqieLBFEn6nSXHNk16v/uQWp/H4alB/zi06TGtST0yWOKSP9g9EQlHR
kZmf/gQxmXlqHKsSG3NOeo/wB3LkjpcaT/w7i/h9tHGEOaQ7aCpzSxm/KTJXcKxrfUT5G4dCQSwK
LKTlJECxKf3sIl1jXW4ljBpqGJY8JHUi6Bpow6TzCjqFu5OWPq9qhk7+1Z/9RGuby/FmS2oLqzY3
4nI0KP+yqCG9EYSCDQptYoaav2T/BFxbXNKunD+OSA7kU7NsT2c/kyRRF/m/FjzskxidXD3oostC
4CM8gOcBh90z8oc5QXinR2JBOFL7AIoK3I6OUwlO+zWY2XbRU/RUxm+Uqz2vOQdu75D671OLpFoL
ZfAF9eFqSb+qxilKU3HOG5SR6I1PCiDMzBVI/zZ0aLAdlIVU8uG91LgQp0JhBBtTBmmmiYn7stiU
lKsybYn18XEhSoB7F43BIGw7xXMMhN5/ljT0zzTg9v6QynSGvwEKA0vyxE4oMjlb5uoSYUjl9t3e
i20OK8c6vp8l9hE58emv8ghZjoR/oBtx4MssCowOVi9Ua6kk0MjiXPs2HfvDsAldML5lT0Nfuz/H
PQKhCUuT1J8fOYBJCp4AMjGamOz4lM7OUICM/tT3NRW6aMSaUKyrboaQbRYfG5uZpcCDkTudHNXC
xrSVIVIR96goZ/CfiSu2pSbjw7i5FHHbSHEBrWplVYUpFxZNni6dTOFhzGkTXMV2jfu4oska64XQ
NDES3w4C+2l/yVbY06wc/eCuLZ/QtmFQTQ2NAQJr5TcUHkGRWCgw1oibgNHP34u0eC/ZyoBe80mS
v5ii8dHc7u3e0xURG7a47FFgRFl/xgOfDCL4sFSShrEyKdqiMYryhvdS5mKtuVS/aESHm694rd4/
VRvZCT/XltM9YWapvzEghNurRF6YQOicXZ1Un+bpX3E/JyzHOEQ4a6gVEps/kQ63uVagKLH3RMl9
1O2zdgnee+xmTX1Q9ayMsQGp+2wK/8PbxH0kiRlmXkUHVBP2lCkCkl8kACAi5fUfiP4J6QzSXVpc
0ktEJ2FGY8O59XsuuDV4BmcIvQHufkI4fvbiAnAq2n1FRFx15BcthQDA03HOwQ7hmfLdrS215c0c
GopZFYbVhh3XRZgsrJhNjJD6vRresTy9WoqqTd0mneyDYIA98Z732Wf4WQKDME+WzrnzpXKqpAjW
D5QYOHALyBBVhcV/N/wWRwwYlW8QRolE2gpKzopFUwU9SndHnMu6/T3RHXgQTcO1ghVKgJbJAAwZ
mCKHjnKarTGbqg9uBT2JwMjGR2M/mlXhpZhVVHvbSVopxW+QBO4uwG+G2zzshYOBOIgitSFJ8lSo
5tDVMiBRTw0+/ZdG6Lpwu9Rhy/Y70DMtgEB3D/mD1R77iPkii3UCzNjxId4X+I3WQ/X+bOFqM0Go
BVwekVAFn8MupwOWspq6im7lrSHg4gu3M0B93PiknihLHAbi67Rt4I6n7bGEPytWc/istnpTfqbI
deIs0t5bSoroAsbikrmltD4kbM7GeAOBhhV1tcc1tXL24sUJyrqF9NE1lOZZoJ/8UVk4708fw3TU
PbNoLB+8H40YFe4EnbMK0ejnI3XaA69FcILn5SCDTlTKEDhwsklJeq2tmj009sIf0VXHJN12/I9x
pqx6f/I9q23SCYsiJ30LIXgYEF0sITpXkUgQs7exBYv7osFFy3qjyGslLDY6Ch9ij0GOUnouWZZG
t7QUWDOYS8+jbBiL+c4+r+Myw7BX7p84/zgrhYhcRDCzyeRELb2D4UQWASoEjd7dDKwhrGcIqm5e
F3aen4rhQZv0/aXBFFLwG9lkx0O9FehdmAAMi6kZBidoX9oYqZjsxwW0gNBsKeg3mHIo8hTkQIXq
JUG2uCtKEB6YMq/k3Pzar8JYFrtEAVk/5bPw7Q2BxGhfuxcNKRzlPze6/6OodatdyhuAFCNVwe/W
L9d4TyavvfFcwKmPOx5WO2yckNXp2z6vHL/Yj6Nv3h5yE0aIGt+4poG+6VPaJ+6F3Pzb54Vz0g2/
VtThQSJebEGDqvPLhSoiq2qkmjMxhlzyhLnQMVeOnDJeF5z9fo4bboF7IXhlg7smc25ZowOo6f7C
Ryi7bquKyhpuN5IO+rfAcUXAD0LlIyWgvcasO+bm06ZFldwWVg9uyYbVBDTSNxnKbLSk2Z4/7He3
Pd+MK1RuLZ2JEVy0iChDnB8gqGUtpeXMflDboyG5+IFzx7x9eRhMHXfthoeoZZO532FytDnoq61p
mLsH0uUemCuLoZDEzLcyWpfSk37JKwd2qnJ9RvsUZMEDcsksNZfXLcAIxvC6C3mNk2k7xds9qCTk
H1Wn7btxUyZ9ECV7z1ZoL4d3mlx4LzBA+3yd1mtCPgOX5wiMT/UEmPQu3G8Yu2gSQ974K8L6FqT6
43SOZRwnehTyqclTfeS5AVhIz6pTF34yJ3TeemfLggf6qmZrYYT59N1G1d/mjRccrOPa+PnzMnEE
VHB/4p6KIskmd92mY5wLiTSn8AU14QUfXE+mChhZaAoZbrmOFtp7UsDjaCejyYugi+fJJPJCXNFC
4L0KiaSk9IYnoQPxtRZqfUn47j5XHNoWReMD+SPyTyLoZpzQ+wwljWULylA3VpCom8xftzxM6HBM
NcLW5uz1K7wa/LOrux8CT8N0lvc4cA4b9ANFhoCBq0iCbut9pN7gumqHaG1eLWaMOQLdxHH9dXYY
Vb3T4AobTlauY70IWwas3/3NY69/ctvxrsSpAA05/aEgPf+A52IwDdPQbbWkEgw4NAmUsHGn3wEu
7+9p3AxRwBigzbgBHOdamVIC9U1+c4AlHwqQu+a0XMVG2654Vb/+/E82GPZVAeU3VAj54e8tILyw
6eTr9yiqZXhSNAJ7VYVvFgaOiSh7X6vG2U6Ecaqs/q7xva/biD+pJc1ECas6UhtZ1d71CSO69ah8
gSZBeHXusbg9s9+qj2x8lnELA6zXnsEBwKcxh3aVJbKPmSACgTFYDODGhnb5ROFiqfS+qVOGzKHx
IAQM+Mpk6Gs0bgYfhgWp8t4laU1s5Nc6BChV1Wr8q7dowxQNx9+pq+ZaHI7A0i7Hv/ielRW/8r9Q
407W4FFNglA9zHlrVv2dMCunELw/kY6QvSuk+8rrcM1b4yD8AEAMnfRYs2zRwOYB9msFY6qayYKG
cNDIXh92uSHzO1312SGpHSsz39xgMflrvBT4zr5b0QKzxyaHKRKHuOgsikHS8I1k3tP5rHano+MG
IROuY18HpYF1yqhLCDuzr7CPhJoZyjljgOtAJgRqzTnk51EYDipynziHSEJJYVWSpGU6oFLrRfu3
TfUfXKL9IPm1f9EasH/MeAbHifrjPbGfvNXMpX3C+4VdqtBkUxJ3pTKZJ/Qom0ZWZN8S9PWI2zYq
TRjcPyKUzuv7Yr5uL0P9NC5MMQUbLW64dqBvDLHRvV4xjn6V3X0ofUhxwepFMXYwBhiFX2lVtgLw
pg5sBtL660uznsuWIcZ2agLs02viBh5GpAavvGnNgvjK1GsMCaKZn2kM6HJOdL0vX1iEnl+0PmJr
tRUZWWkIOpI27fY3Pj+qMnHMDNOvjh3UAw3/j4W6zpanoCeWJsnBQwOQQoUoN0RWc/l0q2fdSdVz
jYGtXU+fskOi7bc9OzG245dq4Mu6fWNp00ABX+t2beRCECVfaBMlucuvKgzPZuDG4RIkHAxEkJ4L
MtzUr3kVMkK14UIT0VHoA1gd7bPf8lJqi1JOBfayWY1eyDKFNFpNjMT2M16S+y6IdY5kERShIWz6
HeDVorLzvhObMfY6RunQ8tF1PactLFsF9oDczmBJf3NuMMo8H4M7Qgur4BMx1d+dsn0s4253DLqK
O4Dubm/v/yQXGN0tPtNrMugH+bGWH8iMFg1QnPec961pAKBPgYM8Ilz+/KLjYZEMh/Kvh6r4jRAx
ipCIWjbEu96KvqeWTg7JyO5UhdRVAPedTq2VxJT7JLh5rBEX6ls5q4kktXjONm3NkxnHyVXfvvF8
6CyjQkiEAi8iRyt4dhqj1smKasK7KlYjxx/rcUn2w5t5YYgNy54WMYqEkIxEuFujXKQRetEGh58a
tgKhrOS/cKwwlx1fGjMiVKsOl3bzpbXIzYp+cuRvW94t9JquSGF3vtm0qzEYrcBRwqa4d7Jh5z5G
YTC2FuA2+JuMzslqlhFBdxTNO3+ohDqD606jDLTjei7bVTCCVB73LiZaSVWIUVTjABoE4cJdyCHJ
isOPB8c2B5OUUnc+F6XLrV2/vKA60jpLHTQ0st0neYPwEjQZIGTLX7jS1XVA+7fNQVSVS9qKNvvx
ioGO1XpS5oLrn44qPOKyylf+CAWh5IXtt+81y/o3mnu8DGDJbr1icVUYcztr/jXg9Jywl5H0OY7M
dSUjykG1MpKB5K3XOjjvmMwTbm16ZenwZkkHY1Oca9PgOLcG3Np/LiDxxGBIo7Px7UyuUdpjRKjd
UOi5BvDq9vEnigJFV6CMUHc80cklWdJ5wCvnohmtnskXPzTDIMPm/iIbVZROgwCY+2MwCVDkv+St
QorFVKIQMmbPyfwfrHovzKfI9ON4wjMlC3VH5vIjHydXSRS9Y2oOWwgORmFphH1cnf9KUq/cMvol
2HzNIWVSQngqlWQzRFYtSTHIRx/U7/ZGiJrjet8N6jDvhpdHLL+VTxmFIHl5Z1sHBxCnowSeq0XF
4L03pfOCwh6nej8F3NL2ysB8Nc6apdkAYt0osHEoZ63RDCGp5xTKHDP8ZTL3Cj4NoIhfZ/TqkwDy
71Rx9opTBcT93ixfafhxisxo037jTnsK7dGJk64RFQvzfVCawqwl8m4NBT0REZjf8EMCEheV3wdu
8VQcKFSkHH8oqAWn4DNaO8lPvYHNpR70KdjeP0+n3B8HOQ/bb95b+xpKQEOUQes+t8wwqQJD+nCS
Iv0QG6y8FlGxhBPcYjqPP126/jHOUJXzK3nEYLlcYNVOoeBY3GzTWI8H+wgMSQHDaM3wcoOnf/59
LxNTq/vnaNu0FJMVI9kP5+Hoo4D78IC1ez+fWu/3msarcek7vxu+rUezefk5R2Ytyc0RGwV1wACn
Vh6wgSisqDrWQQQmg01T0RDVDlxAwbT/6Cc9C4A6Gyc+IFdmgzWV4bvMIyB8Km9R29t2jBUJcoLe
5QEEM+bPJmeaEeMbkvtL9U78Ig8st1bor4jqmBlTmfZVH8UUaZ8CKiVczUBKmN6P0wjjxRwZVdIK
j6Z8wO0zIaDXKl49L+MBIL7cKZEuCkrrXfmfpmP1sqcRonADSs0BmPu83miCRt7pkEqYUZKngqCF
f49nIc6Qhw9tes4pDorgqivbdAbTOwiTAUlOcymrmq1d53EokiIKlQ/z4DdKZSp09hWIoVTtiA2d
pKdQaAMHPQSWDoUQB5VEzZrRGZoY/zc/jJz1AmqHoGNfYD2OPZLsurroRD5FNXm4Qi6VvYEbxKOf
B9LJjGnQRsVq8jgHjAiDmeEjR7Q9eHuhxmuMm9BDSZ6dvpHLwOTM3vAFykX8G4gnYk4UZ33ag0Ru
iXgEqg/R8NoQaODSgr21VQFpUb/zBynemB6qaDRHi02r99unbaoBIbv9KGb4t/JQtFZ+YX0VSCd8
objiBj1Ap8jJMozhxu4FHpUGn8kj1dEuTzH51E41bJfigA111HcO6DVzs3lrARW26v1ttHvoD2cc
6u9nfFVDiFhVw3KJAEXvvERHYoLaPdxgZUk9BpzWTwa2C1H4BRRjv33LnAxKzN3IZq6NicFjZeqZ
hMlsQ0zR4Sql+YMF7nK4gL4EqE/RjwJIDY9Z/JT3iLb6P4Eq79jtjZfp2aLks0dNq1rUkj+/VvRt
gbbcZGZ0tqrUs2CudXsqvnMCHB0Q/8luusNnmdNY+diHh1e9k4sjwnTnZFZiQ1jeX07O9n01mUjg
6sRZVd5p/rAxMreOcacsyj9EbnZJi5l+A/KMYAj01X66awD1GTjMRiPadJBZgLNlqESAmU3vGi/q
mzeM/4G7LvsOnaxXuyYKUtgWuNxW2Hj0mj2WNmehdZFtsAr4GgT6fPJ8cwbkE2l7soLdfVDtbHhg
ir1a5oJNUvyCAT8l0IiYfawRtBtonK24Rp8g2t3Jqmnk8nPGwbMF1MRn0r3SWYq52ERKyYS4fcU2
S7TIZbnk4ev9h5KzUNwHyugncVzLro8MzUBAAObUvjfL9/FgAscD9hzKG0T7xUC+9Zb0DFWtxUI3
AbvkVFl6RjfaEbEu+N+a4G/RtEpBfPs+5V5GJynGrTF/XqD3m9J12xcuenqqRTaept703Xlpp97L
J6IFrTHWVrFMG6avH0tdE8QR07lCOvZhpT2vIpAP+pkS4oF7KGsRywQUhVjWMoV7zSr2xRw+aEts
B3RihZK1u1LuoZngIcOrTl25Al9T9ihK803qtj69i3RJJD06Zfsce8X/iItjvcyrP25wDVa/XfIJ
rRTtq5MqBZjSytEGRtZwyKNVpWbAFq7R/a7dne6eYWDEQ1i5NEWGrPQHeeE1b8DDb3UqYHoV2yo7
P7GjADxYFwZzo6VcUtt9kVeW/2oK9Y4oe+me6y1MmKQqQZpwIoxWPUcKnAh+TJKgdujCBqsxSuwg
0cs+JYgBDnDBswfpMGU1/GMaIMc1hdjEeqdu7FIz1car7R5RnVPTVmPl7/ISgiMdWNdRTtDbjN8o
kxFn28EIKbpHPJ6JpuovQ9WugzX+AsGehYfGaxYXP+939c/v/MvnDHnZXKopUeUa5Xj18/I4Hc5+
I8HbMXw4Xz05rr57gfxL9nbCVMLA9DJqJXEV4bQFA1S9Gk5EH4qnlShSQy0PVimP/hz6kIOCkOFm
t+ZNtWP2YdVwfMEJ/vlUygHMGM9smmjf7mej2I7v6cgL+x+ZR7mXODk9IVIu78znJe1HMgosF2bo
9mJDaPk0wZA5Exsfv+pQ3G9Jf9+TCRjDUh0GtZk8n+Vd5y3DSmOhqstC55BIvGROpETiOF7ZxTH9
dVZTgmEP2Yb/0G/uq8QqMnxii9askMkF6Ch+m98fbimf4FZgItSjlQzf9gX4XiKrq40R7WiBOU8b
hqND5szBQb6DkG8gzy+YH6ZZjKsy5PP8wUbrPUlUyDqhoUcbentoAN+tU/SlVjXk5Z8xnq86fhec
6rO+ecQPm2/DfSegB6OJaaji9FfFA1iNs/SQGOy9Bnz4w5bH/TNxHBqBlqCTP+VNK0Lx4k5kkHyT
kM+eD0pFqQwW9wBl8DSvQ+BtmQj1jMm4wA3kKE40qGfxooNK9w6dCpY6CNuk2CvHlhDq5Mw8gYiq
kaNrHXwvJbMK2UfJY+4QWealq1eaevDS7orTCB79hTPE8kyhIPPSCHx2GDPFyq9U67d/7Zti5y0i
gS1+loelGkjDoXYFkjDIx4W6Q6okPpLw+vVy8sTvCseNK2hnHvwdakB5g3FS2NdAy2BQGb+xSlLm
OwKq44FlkMvNoopUK4k0oqENJYdtX9rwaNO2ZPGZgLxTs+jmAkkwLdXz8Depy9W1j3xEcsukj5OT
x+6n7Agi9b+gfiiLGZCme8twoWnuWOIiFrJylHm128Ywo1DLO29QmZ/UImZelC3Y5UH95ot36e68
nfu9VplGl3WhYQbMLjFsYtT8FKbj0HMl9H3SzarhxAcTTv90Rgphxr5lmb6XboRP0+X+u5ByMMUr
twghgGIgIenOHEUmLPNH7X+SqFW11xDB+Ri6zVXR2S9135KfG5enTLfFywqCKSPP+iktRsUlbfb0
UY8k7y4A+LHPP1DTbaDlSQtGukk38FHqHkshIY3r0oov/BrHFvzKft35xNfFLBoVhqonyIlLAnAs
wO4PhyyFRypGkqJYgZKcRC+B/3vF/8VgHn1+a0qmOE12Ky3FBIug4ON6Axvbq99Gm5kv2ZUVJTlq
KZYhbpFYnSda/Qv/NbZ5b9PSKwhXFXBego1Q2nG9J8mflurcwnBEvrchIIUjEm+/1U33tG+WDXXL
A7T4h3t6VCLY97eh37eLIBs1prm4qYs9wQmLsmVrzMeKvvLit2MwTwQ8qXjOrrQuCZcSsc1g3K3r
IgAOag9GygRcEUeaScp6ip7+2vkhhfx+kX31HpmwctXoIa7DXf7ukqEOgFYDhYFJ+098TzALpk8l
MfS8FO6CmvtHn4kJElLwGgEkpLYuXtGTkhVgau4Lf1/gMwWPvleAgJXsT+e2E2jFcuW9iCGF5OuS
1JFpWls27o2ibf63ovnLssu3x/JGrZJp58xhovp1/qig4YO7cX+LhPyhaa8s2GPhyrWsdWBaWhV3
yR317/B34DoOLm5nvX+fkQwSiJGu030p/PBYUtGeUgHinxQB8zV34UsIn2VE4CS8dxp5trXCX/e5
yn9JqjSRCDkkYd3hMu6VPJDt7C5YGpAJ1SYXYDXRKoYZSEYNVIfFvspE/u926XZqXPLIehzPff54
H4m9U36aQPSZvCBPC0WGP+DINaAl30PjyFPTpFLaNKKQ0DLlxxywTV80NPC6sIn+KbR26pr8GYRx
m88tQz92CI8xrSo0wTI7UtM13O1jhRHgBf0Z+I9NWHFulzxAnzAvNx+ZIq4E23PwBh1407qAMnYN
zK6xq1LyLjMvGgRsMBAZA7nFNMI0CWheQYutorY+cmSqCCvlMRAAMhOe6La/uYHjlrfjnhAUh/O9
C4aQ+Jd2a1vN8+lxWtBfO98gLKrTrrraXIOwn8w44/FQBpZNveO6VFSKNIsW3GL2sVLKr7uA9jE/
IMTniuWfDOkk/kH8SOeltNQLAEol5dinrgos7SDAGI4ApK7KPfoss06uuBIpAPK02dE75d57C4FV
xHIOlwgvm2jXuouUPSpGao7e9BjRPd3w8zm9eKKnmNcomLU5FQWrstN5Mizjv2TDMS4s8SdcAukp
kRPgLvU/cWwNidl8C45fKERjB1sr2fKWNOMtKQ8Aj3IWv1ZSG2xYHmvSV4dK7kh76/BiOk36VHsm
V8kVon+dw0DYGp2wqQcjw9//xNuqaiqaKQzzAldkLVYtHtXSSjZ49js3mtZU0qUAYVkwkX/uQtV3
DR201NwDk24/eyFmHIlL98cD+3jXgtychl3K8LxCAleDDFgpfBXqE1Y79fKbsQJiJd2RL9eKDFCs
EszyVMkFtBGnr5+rGy+7sBWBxFoFd55nuUb20TMh33RWx0Y9KqeOvX4Vl+2r6yy6DJ6Kj39z0IYp
pKVt6Sm6JmAcZnRHAN0EQ7Srt84YtjRv0rQy2SGvRMlVpSNxZzmTFoaeuTXBC35ua78w0ICwNqVR
T6+WuceXdauQJLjJb9TSx9Vmng+xzVL/fyADln3FrZ62++NXCcY79X3SnekWGUUxr2LRfZPOon/p
erimfJwPeuN488mWHsFohXDHtI6h/u9oQSL/oUFOLzCh5VYFr+K7Qb2BpjAi9LdTuurcEY4rCsXR
gBBjKNRkgawXM87uQ22nR9KO+zYbtYd2NY30fQ1ycGP9W6eI2+16kX1qUXDX0JeonP3rOXSWWgpQ
e/eIVfV71mdXsn2d9BR8kzClUahvLEvA+z+Yw7RaiFGy5aO7LpmYucVEgTVRze7i0PfZQCE9JM1Q
OsjzMONToebaJDjEwfVbiFthdUlpNtkFVpsKwJB5OyyBqtNR/Dz7u7TmIJwTFphfKKLkkDUe4k6+
Y+2YuUZtB1QgSyTF/o7nEKjE4MKhubLswx81pwIZ9a8gvbUBpUjV/hlCR54wkkMPN2k9wz0Hhag5
YHXirPNMcLA6MUg7mjeKdjj2NyH1HcdJC9oUTGaxLE06sKPpmAyKQHv3wnKzBxgryQ+HGb+0/lBw
7rytN+ZhAmn64vOL5JFg10j04tW4TcwGSr7zIvgFFcKs49YHpAYguvOufs9aVSDAiFr5VjodbirR
Vsu0in7Kt5VcQHNTcmcp/TZPTkfeMwO+G5OP8i1GX7Lpmwjy+05LlmZpaNa/5VU3pQvGmymLdJ/0
paCspQXTYE5D20GmxBYHCR75SQjb7OZR/WlNrTwzVrYkssPfKdwX8uETlQP0pTCoxA/7aMzYAdFG
98RzQWdeEHxeNJxUvIXIC0grRb1ehhbblXyOun89T9peICtdKxu46ts69Xw4xStWmWyjRmYmHt0M
zlzyW/0wHKRoXJLfGdFF5KfHrfp4omH+9m5WP6VXddbzbU4fvqeozP9QZuiyeQX7UoddAw8Vlx4k
RYdBI+tbr5tBCqGx95dNJan745Fc3SvLwjJIg9awYLYlFoydhwd4dPVEwRxiQ4h3fO4TWW8zwPpY
9mtsKqfDiDLpKNm9exo234TIcyUuQUWtgVYt2tWVKNzMrG8GdEkwyS+rN9txhDMe1eHn6LrA7ttl
4wEaO9mPYz6PVcpUd4dQ+0a35azDkbfs3nSl+MjTKOLMk2eJKADdTSI+3LRTBIKRUqEgts/bdx9a
ol9rRlbnw/cFAZoKqS/5eBTIDzGWOTxwiJFn2j5j9QquAplaf9FrYgklNBA44e4TfTWSJoikh5Ki
POGwgtxg0+jLQOKL1kHiqxbyB8/CMUqASFGkDeaq4CJfUIKTMYtZLTt+SChLmdjm9JlZ/yYO/GEk
pkvj3clrt3xGLehfZrs/xsboy7//QWKPwa9LJIaUPEosvB9HAA2KsXzj3UMkMby6LTEAqtNVvo2e
DCVKT+Y5sjw0VwCYXDcW13muA+a4bEQSD20lw6O2DHLONPWGZhNlApCGV52h0M2tBxk9Uje5jvFB
yqpsKUE5JXSF87aCDC/gnblbTJTbbPPfOW7MB+F5PBXkkw00Dx2UBKVfocdljfmthrnMCNNIaGKE
A6odZnUmTIq23c8+hVnEdWIJUjrSSbNVQipq820hfRgHeFkZfurMlcuMdGuIXtSv6Gf9L903V8C6
i3bh6bJ72GhcW+e4mnAJzxsQ4eKfzgnQNz1mG8kwcLxLcc9NQsmpHP2JjSIf6dnIoCsQxqp8gTtt
9pJrggDZdYhrqUDl35cvNoRhecrTC3bIQRE/cNWkhk9RgN++XlI8dqNsGliEKg0Am/WijGGfDFMh
V/T2oS7qyq6UnHyXUhnyy1anKypwuSV8LKY5JF7MaT2CgDCBiAfo8Mko2RSwzEMchn08r3n9yA5F
/035t1K5H0tHFT2Cn+vhGpqUsNSDIR2SKCi99nTJ6Nbx5/jPZfbf+eRUHuHqKu2YK0pPh6tcQDX8
9nq1yfKJAE7HEhsvNWHN8AGDBd++kbm8vPrZJ5iJaI/pHR/wSaPxa+6UTgZKYoxKqwVHw6hNBLXk
bK9GMBI16ol+qVryG9XihVMi280x083twhElS0l6BP8P5NHUciSnmJhO3Hk+BtT+bav4LM0xNl63
FK7AgQzaWj2geI5fuPGjRnUsFLu+1B6qyj2xvydPly0Bymh2+p8ZqzsEn7jc/Z1ZqFvsKe7lueE+
66YSfpXpya1KKyEv65y9YTujcJZkpOIokPsT1mAWZL7HwyBDuJfrZrJrL5m0qLioN7AIzrAQtgCR
B4Yb2aMyfcDkkF5szcpZOF/9Nr6XsL3z1If7eUGLNqGEW4/rpED+iBfG7o92azI3D+uPzYm7bBQV
HVwQTSsOWfX+4vqQPeWVyKuPW/HiDBbMImXTIY+RK0RT2M6zc2L3EL5Kez+v5i76cRtO4CcfT53Z
ZZCE/18Ldoqw2jszuCU8SQNrzuxPQjyzXOMK71fCpntrWOpwu7ex4AGg5qu2UQ8/LXG7QBCIz44z
RkH/+TUVrBs1QjMR4H6UN7cAQ4Bqp5NJLEDsAIeZRZzpQJBdpUITl5kmVpEWC5IVKDxmJ0iZoae3
f2MUbOEns1d4Jze0UWpbeyetC6JjNarLBBxSDn7ht4u6YOjmKNNKroV/qrU8t5zigymhttcevPdR
8Gi+asKkqI6dYat3Jue/eBEjmHzwVm5W7GuNrryr7/1OADQWLpfMKuf188kZoTYq+Pq4lrxk2SBZ
JrcELuFAhx5jzlwqe95r7B8vcqabrJN4DLmINUW5HI8M0r2YCkWSLrecqWb7ijZY9IJRHHumxjPJ
QA4He6zcyuZmwhPuj1GyIa05ugVB0WUFHW8AZsWW6Jv03VPEcMW8apwUJz/g2OfCFDixRO+yxxrH
HQQ9dlM+B3a0Gd/3GnOLwRN7m5rJe+vX/O+ydvWO4+HHiHRLSqkDzcWjvPv9i7xJGvb0naLikSuK
ScC9l0jED4AoL4Yw5qbJwfN5TMjr2PHIGEicroMtwowQmPWzOUl/V9usO5YkCWwknDS+k82wWw0x
JnbSw/JuG14Rw8DVcSj+zAkeyyjUeEJqW1K/eQ2u1hgjjBMjDzxe767OgTKE10pDuwFHpV+/yM8R
UKoOif1ZVhTrz79kdfADeUhC7bOMZYzy3WG2jnHtbJg441qdA4aS2DM8VbLk67KuzqY+ql/SUQ2f
gqbWFLI1ExIMlr4TopHNRRA1SLVnxdMDLBIEANbswcV+t1DzpKjwXDsC2sfAurrvMJFRs/gGZVuF
ekJkVoZ2uFcZRLxroAWKt/0P18VyGSdxgVcAxZY6qLw/z/LoDNm/QxbrKpD2FTx5BUAuuoNlEi4x
3vkopkUPB34LjDpPOY/yvq7jWsT7ghRvV6MWAQC6Y9XkUIUfC7McI2YOjK8a8oi8BXd462GwcPGG
qnqbQ/jS3wnuzxxa9drIV9zDK+7ng1nTze7h/rbbsiw7LDfhmgIXzqJufrqWN6Hz5fAzAY3oBIhO
8sGRnFM3Xft/2sh/84/JNIb1tZu0uaVRO90oNIVS8RAGZHss3QifqV8uBgtNCLbRh4N3XnNbjv4H
Fkd9rus7ICsFRitC77/5TxCkFQWypaPynZNyu+taNO0LgFq7WgCYV+6LPTGpww3/W/Fha0rLmie/
TneAi2UBism3ola1Q8yY0w+nvGlpl1jeVSycyXgLR8kTrESOuzL9Ll6L6Qa/rmQATvAGLs+XNdjA
YuVgGJJs2Ebpy7id+FxFx1iHcJzTmCRrrHXYeVsMZoAGbbqfAec1kwyDcI7IKUz07bfIpuHHPuUG
3LzYYLY/xY6WVL1tTF3fJDm7PKNGxo65NvZuERKj9aN6EOxKKhnVRJjyElrkR0mAjJcr50QTx1d3
b9Fj+3KgeoUBbMfabQ6pKiXJx3v0kzJXp/b0tpOl+mq7wnFg9MYcnoe/k5HT+mYEk6e/nrlYxAas
CmyfXAKXkYfEuBdXECTTv7T4/qROjivRdkO5HQhILhU6+YUYeUh6DHfsZSVdhA/BlbfttFnFmh5g
L3hHtyGnWyxnAmFPUgLcCCmtgH/YrfK/pETN6ves0LJmKa+ekzwqEaJ4MtrcAqghQOUs3NRau76W
+lxPpioAyXCJutRNyqGJQm/5G/yGFRZLi+VL9mJDUmze67PEbd2Xnc4R4v/nXhCmnnFVLD8z70FC
cdWve82x4Hp/azJejH2iP3gz922KHmGK1FMYdOp79tPVCM64RHKUjNmceOSf+ZKGIuQMGz9/fXEK
UZ4PgSvtzTgqJBwQ6d3nkUr62tS0lnkVJY7OuBQzIXS/MMQhDQzirnd+iT5L6SAfWJU3iJoP3wZW
SZ/AG4exAhpa38N7OJF98+lKoXx+DUYQ/1vqMizjRC4MOdHCYfC3wmiP11FcNhI6ppu0V2h8ErjJ
6C2RdhWJzd3CszYbF2m1Ic3ChcguHLs9uXHx7f6WOJrNro3XnnD8ULaxqNp8+WLyRtOCGuNMW4yl
SWaYjYZK27O88rOFdwenHYuJkQ2tWzsi/Yg9sCJzhzWGwwJGBLZ54g8w6K82v0qAZiLn/N6gllli
izz0qCa7DODFU13rL8BlJFOZdb6xqKxOc0Du/Nofck5r6nRQRf1mNW9QfK7Zu26mkVbLbUvjYlh3
P/uootig66GKIKE91n2HqvtiILlDL62nGiJet8HK+5ObskhNghNWD4jzn+UW9ZgHP+0lYexCC+nX
JyRCbY/qbRQN7qoDGI/LklmYYwGOlYvTe9fEVgah41iO78ZPq6G5L6i/OAhrMuwvvSU6OZUCLC2b
ui2bZJ6o8e9MgsRBv6M5tHWhe082Y45D2WdsivTslvs5ZDCc1cswGaFF80eZTp1nzp9HPkt2HU/w
bDfiowJ3QvpGiODZ9X3trxQzMXvcH2AZSbXJt1HkECOBt2XEUqm6AeB/td5ktbyP8U4CnaaZQ2Em
QpgZY7SbVSq5puc8NuoUoi37jSHNzWpr71OfeN1mZUdkPMRp1610v8c7/m/TjlOjZPEz5qXaz61m
ud9494depuKEHQxAdpu8VoYkF1hEdCEDl2cF2OBm1phx5EutHkOvPzdxwiOZoHXx9+Z4XpuqyljO
/poWtqpyEpP3XvhiDi4m6pINemMiHJkL0cGTjB/D0kK6pCiG0BGX9vZPXU7htI0hFFk6mJAQVBom
ez7AgwEh5s4adl6PscbJ4iuSmfqNXaBGqXMj2k1qyHHIRvkk6Bv63Ki1xJB+wMWJsunFVmlndbow
vlTZdobDDt79TlkUKnEU99funTao6cACv1V/kX2IsEi1kM/braYS8NrYMATRs5W/QFyNRAjtzFiJ
qYgJ5Y3gm7Cx5jZz8zQmN5/NnSd+31zuNlURBTH6cx5MH4HFQpNTTexbcZw2ShMMAxp0WEVYyfxS
NxE8n8OiUuwWyiiLubwlHHchzPSsIlkBNKRXMslx8TVE0yMCwv3eKW2Kc360nL04V6kvFObgAp4z
1rh4eUzUF3RzxzBfSzzg7K0Y/PP9F2Lx1IZCUyijInfK7Ropfjkztoto+aT3yGgnmv3JCGpkRzQK
xh9DG6GukiLZLgqFFVxJXJoXljUkIlI3/nWzpJ5gYGSxttPDPzOeSNfdAqPwtXqFLpcp0q+OS18z
R5QpBCzD/klqzdbt8VswYIHJo9krI19sBkEhg8OfcBM/YO+RLFEMUXaUKNdxO0lGvDzrmqNuNIrt
bR6tU2VCL1A0eKK2jDjRmCWr3Z1IC2OWtCMk7M4zPPMRpuZOU0MoQLfNJb/QAVf0XKiFpWXDzZWm
G5dgfnetPl0itlubwuXVzaLRpmrvQ42oQt6wYjdUnr2fPB7itfAJVBF+plc4WqPsOvK3mvKbA7+A
GGdOhWlwhdBN1Yo0jKtPhp6+WqIEULBrWlcGGCF4Z00Gva/j1+iGyj+zDZtp+FqbbvPNOCiDkhuN
5w13QZ74aEfy/MUw+aZnG3MYMgpEbqGOpNNLHzLkSyh+NJKZaGeYpqwIOxpi9sRTzBx/0EFyMlL4
7m1NtzzKheIbfzzLTBH/bHZkoOH3QFp/NZOTP5bGrG23NUGPdbu+7CiY8bmgutCjaI9ELfVQ1f0r
Lcpv+mhXvCSAebJwQFiA4EQJIWVxhSRWUD2uiyfrRLNoLAKPf3syRK/pB2k6FUyGIRbu47acluil
JlfomlyBVyWGQP2FPXQbkCNnLxVktIAzejixht53IpHGBrzR1uABJMCsxgRRi9ugkBKC3RXXU/BJ
eB/Zow7BDKIGyHpoqtiiy6gQF/TOawu9Fi7iymGqBiDU3wcudOXzIL4TM4HnuPu7n2BljWu4kLCQ
qEFGkSycXuU/2kF1hNXOst4iGrIm4eb8aEpAfrHTUz3PGbnP0NDXz+dr9HzVXxEqIIB1Tltp2PCD
ZhNQ6GYhdwsixEHW6h8Nmdt76pBHLthytcFWW2v1uq2+DZlCff01dGSy+uA77UvYR/UcmLlMvam3
WIWm0Ci9wk1m9iU4TXoOL1XwNAPzuqFN4J85SAdsZrbYx5nY03q4ob8ETgIfDZJY036Ze4saVFOW
+w/lZ0gROUdWb+d4tCRPabFPTgveZKF/FxJIjm5mvbjponol5EueS4F3p6YDrmsLV3v18V1k7Snn
TREc0rLdoFGzonypUk39QL+zuXKDRDtfQqRkZjxvAJrcyRVfo0Ws7MkMZx/dzOmlZBefBuYWuGRd
UC8OWvM06TVwL/YeSe5SB+dnNFwd34CC3puas+biofWf39vxbBFK7ciArJ9aK3lLoZgDCbUIYwZl
BYOluCT5x3A765W4CoEKgPR5rJBgjyAMAhdIgTxRFQt3lmku8ZJ28sl9iAFrCUQR+eUP/akfjOH+
X2q9PzazIzjyusGYienv/MJS+V1vBWCeBMris9pF89KXy2KLSy53tnhhQ+CoGmheaj+/L/l4rrV8
xaS4GbG+IcfJV6WzRZM5uubh+Vq6ZnrKCCmNlLWCzmAhv9E1iTga4xu5igBhR/HRxCIA5oLGhQzV
uFOs9LN8Emp9shx/S8LCsGwYtTNVJHVqGImawRD7Y0UbJ16Tmhla+s7nu8QETbWL5DjEyUlRquHo
PJwJFqj7YQ8B2a5ZK10XPoOUm/nCNPJrdyuIHfg3a4IcTAMU6EiEiZ1R5cYDFdlaKUIqndL3NxVl
0qVEcfTl9qY2qHbDoFXcIudULcIrYeJsY3lThSfJ8B9XRgp8dO/MqEN461w07j6X+Prdanjj/ATA
HLadRL9sdUFJJZgwqfOM23VwL7NagYmfyz9TpwazkijKfeVv5r3ZrF06EfLetA4cmwrGSod7o7rL
Gz6D4VgdFlIJcYDWmmpPqrWMAsHLOC3wJ0CYs36Vp+6erGHZGJYuuqxZwN4LsEsQ9t0PlhBL2Uvd
b8DkAHbyaT9Sd+3I2BcR7W8naz0T1lSW4WfzIgDffKyhB2WDWgR13PChbybOMAzlh2li6J9nq03d
k86N7VaSUs+aEZJVeGmrpgfEs59ulOOcbA1kCFyDk2umMfVJmAxpKzOc7BdJMugIikiaQor+dIxq
isVS8C1kan9MUZmx700HXPsSTzDOI3Z8NUhBahkODiFVjIDfov9EK62f17sJtBgG3RCY0O7MEPHm
OXapd7wRuE9U+ypgApmC4+eUhMRBph68PLkDR/7sLQb4VZp7uw3iAY6AATmxOYTn//IqiWCu1/tf
Db/69E9jrU2SiTdUUkAtP98Oiw+RTScVqpQBL9JDvKLIcurLukYZurxZkBfhBSQXN3LA8Bu/aJEN
JnqysoKy51yHQeYPmk560/dy82k0BiFd1eHam9nLSlQx7fBKkC3c8Fn2xY8A+ya0eElerNlPUbhY
Kkvspi2KuX2UcaEfcSQAyLvJbvqQYaP1ZG9Db6qvrA+qbY0viDurRGg9AhAgE9O9nPR/Pqw2rwLN
ffWxi4LdoPGo5Gfw36g0zPYBQlMx0HQxA7f/+VdWWvmvjFL/St7Ifckn8GkQFA4JoNfL3SevZCFV
lGyfPyi2wRIdkmQGU/iKueyAlu0yrWbiaOVSonVm+OC/osfiVnD7j0K+Q8Pr3U859SAQ6riHsdqa
XEZGj9RMDf7s8jmlGxkKsAWIf0z7swqLdwp9aU0/boex4U4RAW9XK1peL+4g7wYWXpyaBJtCv0QN
SZfFSy72n2sy8odZhTOEGzKwtbuA/mS+QtHIFPe+q0ACH0SP1ktLByHo5/5qva8WYB3V3lSNdDRQ
cYVuO/R5vZhTaxI9gg0pJRyA+uUa6pIa6d8aIojXDz6GnJN+DmKstXQTF1bUuUDQQCpz1Q1eXmUT
Q/UzFtFKye7JyrMO0itsQRpFI9r5k48pZojoYxlLKq1KKKF/+hKwzMyDHEMuU3qAbW93+Jvpxav2
bkVrZmabI+RUHiplzflwT6/xUZKd5VxBC+IkOvq0h9chdmxK0Vl6ts7RymT/7++bsd8w5od3ovIJ
NFn9WvH8u0vGjQD4t8YW1rMIGNrOQyLhCx+VvxwIWYr0tPq9y4/WbZtSofeVVfPWViEa2/S4SmPi
0TqQ3worsi8MHKajp6KEj0k2+4saxOwysstOrB6zRHgo04MIG4ooU9rHtQ37g+EEvbC/mAEkNc6E
fYN4Z7PbPog2rtMajs63PxQFj+BdIdswwprzdbqD3bX8PJ+WoB1oP0OEzdWMBaebrwQ4By89KuHk
js3/+BP+0M8ok8BpjgRi4Mko1D+iaEcHDAvelXc4xoD46ApvHhZrlYI1FULfG3aNLsMeCV+a8O0W
4duCAObaShFwIFYB+791V6gjGNf4k6XbzkrNt/EkptUA9eDu3yM8kyBJjfNcPeba7bhY1vCZueJx
R5HdgWJYYpbDnz3zcKFT3pBzKkejiViZBh8tSi2PDM8KQdqluN4mkUtP/BeQ8UIry3GWuWTuUNd0
ZvnJp/yRF0sVRAj4AbW0tE2xjMdoqRVvatovCxhhdx54VItpwSiCuitOioAViNm0EJ3JhLHh8iml
CoOpTCWmObuUS50b+Ml48hBW6TLvmjeK3laY/k44yTgYGx4HlOwaMqQZX+zwzQPtjQAEG/eLAHaV
S+zLD+f7owcRNEOJjTZcsZ3eAIm8oj4YH4Q40okEIAiMU1DPl5cQtt+hj82LFToj1L32ZbGuZnrk
Ua3mkFsAR2sxyO1Jzpny3sPtftdtD/G/ErZA1yHouUmEzsC55vL6TC/j1hZAbXb6PAu8BFNxcX0A
1vChO5mYtX0eW7k94SF2Nv5NBB6IMz+HRSe96LbB1mwxBCuF1I5pdpWwnbQVKZgkuB+hOOqJqxAB
ePDqQr0DvKMGv0Wbk+xeSn9tJD8VIlXoTj9xBTVgYMuYh1qMN9dWiWsjc7AFXEGA3qjOT4XGxF7k
7hc1cZ62lkZ13oSaH40fu0MM/GhViENi+enmXHlRvhgSRMqkdCehMat764BtKPbE8DVAWHEJKjFq
YB1yrMvpkRElNZaAgIx7reJrDo6O4JjOkt2B22C5LUYhKGDAE9fAPB53pEINFVL++yxpbWB/x3Tn
MGyv9oaDErZARm//I1vGdEuyh5KDU94evPGGB2r4+tKwHvBfL0wOgkdHF7cLJdzg3iFiz/JvIYpm
+IqoTYdtRYnt2hrLkE+36WhL2hY9Mqv7ZgOiohvQUtn1laU3AmEGXh8Fqo+NKRJZ67aNqgoVDBNp
x3bnzxy8QYq7AYRkmBMBvv9iT2Dzi1uOWARt0TQwu29is4GbFaCDagsBKyGPXg5C/OYJOpvSTPhW
Rbo6JDvcFL3ndRp0IRl6w5lpKlmKxa2TxlE5w9K1zVPts0UbXJLIxFL9dlCsLopEbGbDxE9aUH+V
WFPWTfWQmC6cmKRK55jHQPxF8pkJ4mHQuVywP7YK3EKPy9Qq5uS0ic+H5iae2Rwv8hlg0ZK9FGMk
JZYO36P+g2pC63N21HvlvnFPPJRe12EcbFLbd/5o3cnGUc2t0xLuS4x30r+F2qd11xrwhPIxOLN+
CIRw+X5KzIABOHxgzFFEFUgjYeIIt1VMjnN4h7kH43+4oSceDVpr5LlZFiHfw7hDmerLQ+ekp80X
rLMxkIuunKqLSAHWyN/4bgvfBy2RqXxh3uY8CytxtT8xk+fI1tPNmQ3MMqKhlgfO8DUW2gS44K/D
A9G/yv0d7RExMiqVgsi3zcAMtd8Weg6cANBaZpzR5PmbKnhgPDm80OWxl8dPa/j/Ctcb3FUB8RLW
XabbPLeVlDMzpR0jGS6Ke50o81lfXYOPL72ldvxS5dzrzy4K5E708bpqlvfunBvgVCgmqfZk6rlk
xfKBpcakhIU3tQU5A67tYcTYFGULPVHHlfXJTsChBqP+0+bvW89qVdsacpnyURu5l5RMOOHak4bV
RvUsRKD3B9bi72ED7L9KjtjhTKnrNBolxikN/Dd6JHl2L0BhAvto0/8pyfnQHc9EvLoVg2JHBlF0
rAxCsY9rH1mvkPVfzzsfRHo4Y5z7zuO9BQWPhYRXSx8gDRzeOxtnB/ViLR/d9zb6JmF55YWqyFS4
RTSXD80sGU4MFlzIyiIKDZZGTRSzC8WJeiuR12t+v6553eQXnKT7FSDiLtFkXxL0jE158lrqKuHp
6H+vsRnRX0Zp3b6peCnWJ6KJNdoCSY2lsmBqIWhdkG/WuMFvJVh5paQBsmSKnB0dJ54r6mWjFXha
WlkRGjISZmAEbfhREKWykvxFxjuhnSNRKiyF9ObRjTrQGlS7ACRwjbB9q1JbkmnIsw/URO471rns
K2z0zEaImxBNMC5NdwUTH66yjaarVv6W7/vi9caDoMgOF9J4Vo0afT7IvUaI24Y9AsJMPKNbAkkH
D6cqlIsr1dQoZCsVdvfNVmF6pe6VkBSEzcJVvLxIm02LiMyz2K2cvXwITW+kcJassZPkmYVSDJyn
ZcKOj0bvGf3/Vrp5ZkkXEWxF5Z5l2chbGWOG7+XyYhek5SJH4FWy1ubk4fO2+sRunx+jrPeeoE0b
QXM/FdEr/cFiAEuFW+WpDjDgItrwykmSS6+o9OBt4QLva4TitHHjIln54Fnvliy/79iJ6/gzv62U
3KNISo8bF1eSGGmEkjZq9WXSVq9AR8Ieb9XImXeLefXtyAt5sHFfgKzjPZFM20QHLcH7/gU1YvAN
z3NimxrziUDyKYq/od/605+3eGAMscMmrJs2GDXT6M2uxdXS3ClpxgyQKINC2e65NRpy6IfdMxG3
QsvafR8jjhG1DCKBW9XYdOxVsX18Byr3kyGeeMRIiq4dv0k5NHlMuL1hHuwQjQB2d7vtbDzQc5jW
jfNYhyx0Q7w65Ny6NfQbGhtTLP20op/PsSsP8ZJt9TmGLiDHT6tKT2OFtL60MRtIZaPE0rvyP3Pq
CDbXFg+vCPnfHFlxf8lzf+Io3uGN+8X0OPJZoAICaL21sl7KUFvgnSo2slk1MzRxBPrPiDoXwC3K
XipVxNvGQx0A/o3sBsSWNI0kaJvDWTxAu/99UB8EdEnKx02QE6tJOr7fw7eLctm1xrwbWN544VRk
qha1AxYpCJVmK3yidi5VFQ4J6KFC1VLlXz57KS2KnFJYD6+Tp7lSKF4CdnWQxhYGo+GACzbmQCcX
pjgJJ78+3WFCt7zYJoA5mYm7S2AJXxzbnlh0mDX09+xZUeoE+1IjsAR3kcMAa06slsSTA932szBH
lnMIJZThX5jAf2NZ22r2XYC3hR0oI1QyOjJKZ3AsXWygo86miWwQ1277p6KeJrOdt9lrl4VQ+qyW
1MJbSawWGaVfUBO1lIMD1O7Bg3PMhJkl9+JWZRz5xQZtlUFlA4TTgNxrGMwgWWqJz+BAjM2ltoHX
JK3ZPsuwErLh5+bWyJDBmJKBaCFc1nkAcTdfIl5dHvYn+v+Eq9xgElXGKm1JNVUfH9Nv6kroZ0s9
xI7VjaOj6+qgV3zKIRihY+Dkpvi8bpsmZG1ZnUZ6PR2jEu+AKsBQ24HYHx50vJgD/ubdQ/u6H6wC
dagpxNViSb7BGDEKH7bBlYRcncxirZninSxMtG3Z/uMIM8+/aT1KpMxUWs+/CQYg0O9Dp1UisEHm
OUgjNT5aVf3Js6gHVooMSnhffCkDazrPEcGofRvrGa7DyC/g+qrhoicR+4+f+IcEOtpiHCCMQKSw
bdgJURqAdDRZaYZIm4mecap18Pf+u5mhMlSNsk+NCqojPuc+xYqlfybrJfTvd7VXQpzOWMt6PHrg
hMgBF1VMxpu+qj4KiCjdsdtUeNHVZoVkP3bz3DNTJBXlvqcpfTAuPGc7Snrlj6JybUmqYurz/i/o
3hjDQaF0KahoyZ3TaViuzIaA5FhnxVEEwJy5gzW8Qui3GF1EkprkGgmvvjgoWYFon10qiUhO7GqU
CXp0UfsBoWzL149Jis9LgCeMG93XHamBSxhXBgvKkpGl289QJbsEb9DUc1GpGDSYtxoyTqHqAKo/
G3GPiZK4kKetGVvzGVTBzQP3vMdlscn4noZOtK8txs46S3nuAUOKi0MJ8MptPImr0im2EQyV6uKe
CWEw6wsWySoKv/8NXlKMs5ib4BBwVCa/7UUgvFb2IOoEDBNfb3F4PlUqF3VCM7rMIzmH2gRlFoVe
MOBbXZjT0mPN3n0L8l6q/yMhJ7es1Mvj5sLAvrWV4joKYJxLfWj5Wd98Xh5dJiJk+zr3GF458Sak
0mp2u3Q82zQcbe8J5EoAge293qLza7ZFaqdReGmU+FLKqSxPOkwkiq59FV6TCvSlZUbrdYn1d1Oh
1GMELgVmBaQmyHWkKXQXhk/2B+b+i600ywz6GiopNMJ2zJz8eZL5RGzXKQI5IsBv8+Wb3ec89E/9
lBAlOaYkIzZRfGARHZbLPOqM2NFRTn1n3Wm8JtNl8Yrxe32TAq+Bkwp+KKo8kMPmO6g8iYff6j8r
ZSAvr05fcIcMdifHrYgIrwswJTqatm7Uoqy5a5OUePbIC7y94/aL09xyvFSkwXlec+4/+KaTtnrH
5nsFFOgXgQ6HZy3ZuKX4T09U/Brx1vgeUOM2ym/6tzVZOVi4eO3BCKuerO+xLfxy4DhZFN69vDoJ
Ywkxuh9o9zWAXYHn9wfXG8PnQ/9dwmF8KI3X7vf1VU6vZ11zQYyu9916VHhcUmvqbp3y0enbfugi
0tCntV5D7fB32GMsLmiJo42qeJmepR0E8aTLPl3rQZMP+vnJ3cZD+gNp6SbtfzjCOA5u3sJdj34X
A8C2kGJ+iiI2aNAseDNYB8s8+MSooQOgARRPjoDX3vk3gwecFZ9KOP6fU0M3DRrObCanJSIUlXdN
QShVD7ID4M9u68Cxx+3qexeub8XGY/qD5K0Gx1MHvfZFrM9XusSNetgMdo6TteLnkrca0JaPy8Cr
4l/nfvt4e7FOnchmeiZ7OiLVE4ixG5+/4PRXyByyxwnqQhCdeZwbsCR6peY3DZGfwZZFAismltku
i5xx+IZVOt7hLgx+BwNe7pFg5CdDBl/TSN+dErwrkeB1pkWoqVq+69HnS6oWQ8rgNnv4+ORHgkeW
IPz4w6G0gmp46YLTJlhNAAkrfHuqUe/aADxbcVWKCIWkJlMA0k8qPRELHsrNDGrHHeV0Di8P3mEO
DXum2xEoskM4gh+gtAV8DahSR/ueiKct35aKwRA2a0+dB1CLzhl7NnHNlwOOzKm7gOh/LFV/aIyx
P62NkLoI331ML1i+aU3kjrKURrn/a61KFyFofypIE8LqkmhMuqY0JkbpYLY+aSwqxD63+hmu09ei
iFN9N4GNxTF6/PZIMJyL1I2bCyGVg57a4RWp6GXLvZdz5saF2+1pI4grfSb1UeLu6AYXd2gBDUUm
VG4ui557tEPwmLXQ8Gjb9fuiuePDROJyR2hRgXBbwIjzY2ym/5O2kPEQIcrcDtaFcttrl+y7CGI7
NsbuYCVNNM9BZeBu8Ala+Pk/COpBEtrXHZFHsjYAQiCVReLD2xpnWxn4CJaOvbFkrOCmwFSOJMLB
GEMRCicxpg8wgt6IaDxTSZm+APXrfSAl7sXLxrY9gK4+oWbI/VoZ2q/JREaxsgtVKcPoFwd02B3z
ytV2JIxaF8pwzK58g5Us24eQG6vLdigSbk6BItx9HxtkIqJFyTbeyzJa9Woyugt+cydZp9+YM25y
jLw/vK6hrdTYLmgeUzySEkJSAFmpwmXUgrVGrIIIZavNQEWC4UoR6bnbaAG3nrUTv6vCb6Znqq0S
Wl8xqVGLTUXkVnCaV4DdIZ04QA9MeYl3ZrQXQncOLUwP60TTo72YoMYNuJsL5vwqTFfV38hgLtk6
6s1jiMP6gys4pTxt7ueczwttjBpn6DH1Z2qUyUT3Wm2kT3dRE6bBUz7WD3e8Up4T4ZtuxqDbOphW
T2eEkI6g1+NfLztL7N1enGtg/ihP8nOtUgqk8iq9hA0Mxblpzn73RK5W2vymeneCgXzyeWH30vTJ
QfB+PDiMSDV8Z04abTegGA50vzrn3Be+5pBxCx+zvcT4q7SJTvuYCVQGbWcjdAFtHAOX+uuhNbvt
heGkKNK44eOtEpjZ7XH2yOIxywcyh/unkC+qT1ViVT0hCa3XmVNBilBDXmYCJx0teiTtHnRHQu15
rwGQHtNXmPWNGWj+hYm3Li8ubdZSssqO3RGiu3btvxw9Ut8qS1ogS1kfBhDahgbh5Ze++OI/ninh
hO7oeGRvVxWgGF8GOkm82ExlaWPHmalDDs8kk82QWRhpTTIU0XaHS8giR6RxZBDXqgvfKuapDprn
UkJYt3fxEJHJ5Je9NQGVS92fx6jQT+yonbwIg2FhZb1xb5+/4siQkpJ+drkSQQ/nShK1nsJnSTjw
JVydKqHG3yvmJxqfgLTJhpXQiFD957tuCgFHLnNCXJurlRB8+r7MKllU9RntibauAdIae86XvMkn
eIAiRG2IWvb011iURDM7figAQiu9wJqYCbaMgCa8YZt7681FHx8QpDVZOwsznVUqj+cYxmQtYAZf
EKqNLQzC8Kg+QsNTLuKPLFcdeNTGyCUNT9AVuVAEmCnFcmGDqoIXIiVOvYheOU0ma6NWh1BdgsZH
Xr8PDbVc8JJo2HnkWX0PyAOOz26XmZ2INR+VqDVcZ/o9gI/Ro36xkKV7jwEidSvsL0R8u5qByyTz
LP3eQgUxRwCEhn8fCfBGX6u+asYgbNwvjtbWtxdBRRlUdWW4PV+Q9O1T42TxvpmeLAzkpCGhHASi
o5VoNbyx+4VhCIL5LWBf2ugGI+ZJFtNmLrKtDLqDfSs+Eoz7zmT0NBoUwRNX8TmEQIRnRXmnvx+C
TGgf9yQniE5NVEe+grD6XdYG2XjbJ+8qZRMZhYqJBY7FkSlxv45ZxhrF/sV7PBiWNCIPBXRT6jzh
wzaTFdorR3ZoyK9uS2wjn2U0nq3N5eON2JqgD4/aLQEAmZ5yLuWXoZkj+0RZmrYw1ZbBAz+RVSJY
SMkp5AaSsjh5Ktvj3Lkpx/puyR9wvRZGIPyALY+A/yPYsOKhB7M664XMrVchrrldC/F5i3UywNPU
m2IQUUcyOrvQMfTMFz1F+JGlnngbxAF+oIhTTkrE9ZdLpIimpAkGyKKqJDjoEtVCpK0fWV1PGzxy
PjHLPMWJt2Tl61MN1dzzSlz4Z3ZmcPIkioBWmhzOwsrca/+Ofnz1K4ChTuw80GyANEV8fObPIbs7
hEN5XwjCsqvWgbGkVip0RmXycq0kh//F7EbgLaCwypgod5U5mJ0YisBvKq6Eiq7UAYqYiCUlykkS
mp6aZXbcuwe/bOQW2OOAW0UlP0PYwP1vObgKGFmqSD9jbhF21kgf1bt1Mmpg17MGuM3A3gE/znXn
tMttKhfxXoZzxFDgH0z3VQLFAO7vGx4IuVyudimfEVtqMy6jHPyE3fZ+XwUbSvD4Cn1YO2FlmVZX
00Ch+xjWPMNXDdoBKI6urGGlBzH/0FZWXUvRW1v4d/6On/ygDlKU883xcTRzqKsPnNU7Pj6x03JK
M09Eo0tyhR/nLtEKxpQAK8smRhNzYofSijn30LSG32bAmDU88CtIerd9Au95BaINH24KGA1L6O/J
b16NPIzcMkzrM5VrRL+Sx4zncYKAV+1nSiYHF2UoY4AtwUb4t4HNiLCzwuw947KRzoayBJSS4sWy
Y9KqzEBCmSDuOWi4yVCfJpd0a6LN1JKDFjwDpK6WrnFn9DXQMymnMjXqZnWHaexjdzLg8DD66aYe
o9g/qONxFAZDb/qdCV9/FZE5b5IW5vL8ebDIV9mPvAws+HCF/dD8RBSVNtIGCfS/Nlsv507fIpL/
u1wMcYt05kVg75PWqtQf8hXP/6bTsx4M38xWWowh+fCYB1q/E3IdEmblAfVGB5fkQVQLBKcgShsx
sfV+ola0U3tEhbEmZC1ibOYpWFTSJmIib0i91J7aeBJEt/pVUAa3gdDlTSD9R3duBhz2dzYhwy1T
bU2HzE6H27lBRG6rQriwEl0HIcvFepjaBpAUBUbEYTstJZP2HOTzAGtuJumYJe3xfq4QpMP8js9r
68/iIjQL2HUffxICYBv/AX5qeWUpkjLTgV5iJMi2i8xcXQnqBrHxjvHkf+TixSEiVwP4z9wtd1sf
qY3COBBBuXtAJG+k2zejEDzVkOfnECfqzs8sYmOn8Br7q5YOrVWHVwqFYG5QIALM0B3FfKwceqM6
WaqM+zDjrc60yMeRyH2+xoKNgBDJ20LvOLRyISMNzyfkAVwS1yTr0GKz5ezgDPE8JUtLbQ2zTXxp
xmSoSws08/fXzwAQHLFwN6T3cny4vWU0t6TjGpA6j3H6mY/drGlXD49qUV+c+/Sh6HoADDBWdhe3
L46TNwYUwwh8p6aNaPdEhSvQN5r1mCrcBmHYs7+fhgXboVGJ7Du2j0h0vKUdn0tU/Rf1lEDiBPI8
NLHUyB1gBIMAaaVEn1N6PVz831A8vDwzmMqmziU/ceEDaGoFXwkxIm70Od4QLb9L7c0wkQoskUQm
hF6KRAam8+O/7QU20UCi8SSgtq2lb7K0foUo+y1TNyZRjeBTRhYhVifW+bnirfUBrqiepAdZo3xb
yqAXmwI3den1iCoZrww6Gl0a6ovHD/SekCQ4bL3urR80MOxmkyzeo+TLRpe7G9I6OvUcd0hRISLR
jrTXoAWBCVAHWRFpwGrhkStylBId5upzMw4bMx1r6oVPeV6VqY5Gm3Vqpx8dRdyKFztcUijWQjsA
8n51qP8MqGaklR6BXutJ6Mnao+ARRg78NZwfp1t3VLSK4mkldtY81mKP5NyawdS6qU778cgzeMz0
Y5207E7HTv+ZaqSNp7yKWxEKmvTI3QsLK/TAptbxD9Kt4QlGAOTdgvknCP2RrNsaVM+siqdlssgl
2F5cpqBO7DPO1tdlScp1zisKX/+kqS3X4ID6xBxt25MMQm6aAQRZ6oRwp4XPh3guG55X0H9jEFJr
uELEdLkQ5yVNx7TdYJAQhX0hb0CT7mSJ/gECe64SuKroyKZQgBXMc5Z/zuPaZ05fAvvNEu8zm8MI
saEnoJiMuPcxU7Ebm7vZHoTp3Ov4TKogYV+TtFf99O8JPfv3rG/DfBvHiTjPysVMna+AnMk/2r6D
wxFVClR571lFXEaXyd5cqVm+rdunY2aWvvz3LtUTnpL6OJ+UjKvUeD23GyJFYk7HjlfGD7P/wnmO
2za4cNkGXv4NCE/eSweTSbG0VZwM3QzkXW6c4ep9wLOi39T1K/NAEQ5g0u2s2JFlk2W/ZqZT+KMe
cN3Taal7U9MH9lH/dwYyu2CwmxrAyqbYhDyhrGQHCMUEjKO+Xe8pUKeH9QAyvMRby8Zg0hO/kWr8
oLwdxLEvpa9jpiol5pYkQlvnT5islGrLl0iSfVqJcKkhaEGNXgKK4TKuiSY81utY0sAM6GGXh8pR
COMDRvMT0Q7RbFBWu9cGyQAAAzvMTbtCSKH0JhLA1ZHdd35NIpEimAge8kO1y77LJaiNr1+T4gw/
weGUPvV0jSK/KBi8vfATRHLB9cqcw7OK/r/g4pGQb+1Vnduvrf9RCtn0wjBx/kFbtRA9nccM5OWd
r52sTHjvnmzeq7tQHjck1j24BX40kF7W7AIbKJND5Y+SFErFfARbZtsYi2ir9+YU/NB5qbwke0AL
MGqldDJ5rc72onH7JkgkCKnN7SN+8/YHT7HV/6u+UPa22CHGjL8Vip44WgsklZmUGUwFWpI6BYVi
LyG6NCEeA4/1ZnGbgmQmXP6DKBnTPEkVZk6xkEBap98dviyik0wHZ/2kITNvvucAwrihwjPUy8uj
pFGz8iH3MNnRN2Wx+Ms27SSu2ibNL4ynNRPhLpXP9uctPlbRDL4dFVu1+s83xDq5rVajAcr9LLqQ
lmWY9m14kA7Zqqx0gCa/yfOwkpWwge2f8t9HAAs2rzJKngWVqFJl14KotZKLo/4T3oP6lWwBBERm
Y/bpEmwH/1DLEYg5xXETN099didJBp8yrrOSrD7zGn85odMolEOvz2696ihXf0oZivnHEBCfWdrb
ceklkaMZ17b/kS37qz03+lp0QQoyQt6Kwnk32sZrewseBn5CefvkSGjirnHUR8yuGot3X4myyqOb
s5VykTVKPAEop22YUSOkFlIUJMt7buACoJEZ0A870Z9SKlo15WI4Z8tpsVzHBMV+qe0mPXti4Lqq
53Cy/MF2PSNnw4coqtcgEaEdaKigFWavu+ryQAAKrPdnuIueqkLqOgYhChSOX8x6ElSfYOe78vgm
hubqkrGvl6Io/nwMdpylQqfwXzfI31ulWG/JpSuZ/yxYj8+gOCzx5+HLPBWPC1zn6GuF+O+HCqfN
JE82hasVF9RUyCM8xy2sMHBGFuVxY2+5OXrv1nQpRHGK+Uv8a6WZybv6Tithog1YTXsLAPupDuKI
QqxyMHCdPoGRuRVo2vL8QNNYR05hNtEPRMNiRIcVUi0WWBgzjL0bqTw+Rf7t8tcnQiA2UPdCMxoD
3I/0kxeYKI4CpODCDOP/d4g2uM6kPjikwQ+UsSK4DLskq4yQn58naqQfYktGaEdltUOJO+kLLo+f
hC1uY1zjAND5fdqd5CxQl8PIy4lYVRKA28Zhxfi4UX26mVy3lUN4vY8efofAMCsMJ2noQPCNzuVM
P7BmXzJT27872iiORaEeVt4mLM+PXSbh8+4a4/hM6Ueu84TIlH9io+c66wzZIGZPVY3Jwq0Nwgi3
ZFF0/ewSONgFTurDVWaJfMPAHyafQx9xqo4epTmAvuEpCUolrYXk+oGMf+kHR+WaZ3/B4ohkJ0AA
WwSwwZZuhVs7bu/qXx30D1uuqqJqJnAnNgiaw2oxyOWTtQ6MOIZVDAt9TOLlsiJkoJxHVKqbNkOR
LBW8G5dY+1jNATmJyEYDF/NK2t4fbRyvjH7+RC1juxd8FHjhg7PlbeJ9YplKn8+AR3D9DzJPgC3v
jGv3f5VwuszvfPw0ynk/J2aqatiYc0t8W7UYj12MfsyJnsYBzncEwjEVPKSXbWcrwq0Whn7JntMz
GcIGuR7mit4p9mGr+WTr+eJ9TqehiOBW2WqREh6HzUN92esES0m0hix9ysPTS+ZsEcr7ELKFL1Dc
zihMdOONlNXUr4csgxz2VUmtqiAr5xp87C9JVk9DqgRZekMj0z6liybrPTZnBxrycsLOAbbquFgm
Qx6r5OQTbChGGzSxkcFTk2uzB/9uCigM7lVxf5xZmy751HZW80fyjIL61UuWuQIJO0nqUVziJMxb
Ob9/u8tixEnN8zzGuJNdcmhFOaHxCtoLD9Ov74eQ/MHQSnhKNeul7E8EXNFaoml2YqI2K7f78GsG
Q6TOsXySKZ5iXgxyed78m2GiEmjAdH+QPKe1T4bSgBC64y+KqDmrkLE3IRTvCuyVPHzEn3ugIOKZ
3CGr0gTwuEPTJ88dCVkWKpgG+HlkwFRzkK/flpLzSrCYGyDYe0CNyq4yrypC+XXMiyCSbr3IPelz
AqV/D3YptqzCG+aOQ4Vu/i73gTcTvPHQZwvkhT8lkpYsFgRn9K27mL0Mb+h2ILZnHs+EbZgL/a3Q
UrRyzUvsY1Djz/R0VhevqrdL6lLoFc3niOqvIPPlNOqMBDYhSFHtUS3J26h478cy5f49AFCwcFlW
WM2+4a4pBthRp2zYk3cy5wzltUMEjWp81oZ84tzdDtgI7CxOJndIb3QgcW4W1HfvUTmyV9OoqyQj
KLzSuZCK7t21JtHmRDJVqMIesoa5im+R9MavkALasOoDeBsgneyhbQBCsnLxT4hMIEyZW005cinl
oogfIgx0xezfoueV7RVmpOIvGNR7xCi5Bm+rfJeGmUoNwP+J6sceqXRIp5DroR4vMkXl9cSXq6t/
87e1iaWBf5DfnKPre1Xf2YZDBGn9bGuUd0XrqKRbbXuw2OyedGPYoopz+ixnxczxOYr3ABlwSd1U
GdI6xuLwOx+sejAYNas5COAHxIE+Rf2AMDi4jETjciJGaG3sBV7QUwyVh1Fdyd9QO/WJjiNRrzMN
SCKHpIqurGVrGsnZWqK4emAHhkDfGvG6BlC6E4aKp9L2rwLrLuBH/6nb1S2EH8khTgHllB9h1Xcm
cRXzjJgXC1L0u15nggg3r/ahVf04vSoNegM+SeiqlXez03H5CKMYPIzXdPMT2EQA1q6niHsvunpB
eKomfKyEWlUkpI6gSOpIHLGRyO71La1MvjLfzfpQmSXJweJd+RSui+Czd2X9QfoWN6lVmlDKIK7y
pM0NV6S36uM4UnugwOjLj2nfNc1W7LUxyQT/nn4UA3tdvNkMKXvWy7zazq0QTMmc68lHOssUJWxk
V3hLGmVAoVkJATjunOGt3k8ODUBElsfF6H+2EoNrcNQm3zm7SzbPm7BEIHgi53sjhrK2dY/5Yb5b
17N2Gjil9kzGMDMZghazUGnFz61kNY+idfSmc7/XfN9pUYpAm96jQzYPGZrh4NTRabzmSMReTXcd
Np9x/elVwNOI0rccF5h+k/pKJszRxvLEJ8l+mer0qxduq7EsITyG25neYegfnor2dZOTm5q4YRMj
+jTyKM6Tqm41v5wgbi2f9o1PKYk0dAbCAr5HnZa+hik6iikbuwR7hPzFRGfTHXKMoOFV2XUDfb30
9IqnSjEaicBV1NQi+LTDC0QHde/lj4vKiyxRNk+vaDl6sS8amycHQgDCaIVIW1xUL/5AOOitTyJj
7G0NMI0tfqIYcTGcV/oZcC5SkMZ14Xz/GCqFIZ42u6Yg6w9m/zQiIjT7XIVVdodK51J/7ctHQK07
GCmz3DPt8SidsU35NN7CIpbpMSAZ28/AETK59wZHjjQB4EMQb2pLJGurjE+FMlVkhExLUZ2z/yV7
o6HrEiTmLaUey6pp/a7HWYtJL7k2Q2WCBlXMN9DUM2X0yp+IFxCg01kXdkeYkRMQ5VQIjfrvbrxC
WjvBPmcR/8noqF8zf3NipeHxzdOm+7M0mPwcyqHJVvL5u+hI4Y2PffiqlVjcPgRLbyWtzHF8aCvx
neT9d55UX2/Y5SqHSKF3cs2N0kLWmMI+eH8sec0Iga/uTxOJ1E0rNSUCuekd43OXgc00eAdRxuSD
LI2oxQTu3Aj0p6PpdyQZT47kehyTGPq9kSYuyh0+8/LWXxc0mtYMQYFHxRW7RK3qFkZuqdPcmG5L
tlcRoIXmVjGDZg5roqnPDJnrnf4axpu9sV8Lnb4ZVUrcozgmL7DJvSvHO34IWE87hECZardlHAMA
GqHN+VSJ8fjweFnexDwTTG880wdiyDijL7q9kdR8uyhHyySSkZuLorSlrswoRAJOPzdL/sCwUQ4C
MouVYqGnpl2wwV2fgAzsnu6K0GLhTiivBIH9ZCX5ZpaY9sEjiXYo5VPFbiT3I0YX2JUhieJ8Km7u
8tglGq2/WCW8seq0/di8cRKbttYAKHHe925f4RS3rnl39eT7FGdP93QZTbaan1Urfn/tngHGDhPt
2qrhriNS91QPk0amCrqrdGdrQNKgzBaYE9lxGgD1Z3InPLvqJsI0gGh3qA6SvhsIDg38/IDQ6gwH
YEszKmvrkE6g+AQTJmNM6AN0Yjf3V5Sw/+nI4UudhHDi6lIFtf2kpJ2arukWGbOdMh6iiIyF9XpP
Odb8L5G0olup3JLobqVxLeY6Lp9g/nNAi1VMJeITG1/QgRk0zT5cKYCs65gDoZTKclDuST+xvIX1
eWbgHIbcXXGTmerIPjoUW8N2MlgG1D/akQwrOWhQNWS/8O4w126MT5OB41tPwCQ8hNLeuOjfjNnN
4XPWufkbyv8OlTSZLAKJbJonyquOyTQqMo0H6aFJurEuKmStLU6vsmP7svHHXSmTycTwSzB8ERX/
a658NVqUBJdOrQjD98KKEau6Y0yuOxZl2AtHzYv0o0myxbqHFbCCsnrEWUhNKdavnT+cG2j3lLkz
82E8iqJEZHBm6onH1rPCEuYIXkQSTIuP5kiT/etbWtmLg/wsLgmu/uC7jNI+b9/nVbY8URZTNjjJ
i6f0IHm19emLIAQETSRqGnTOJMV9cxIwnMOqU6I9zhi3gGejw8RQZ9g8Hmz5+6k3WUIBTUZEbzp1
xYaQ1X8pA6icIrc6f+FxFk14ckctUNv8bPROpMwa4hcrbvCeDuOjFhaqZbWOjw3xF+lOWzqDCTpq
IU2rfh6ideOMQbCii1QiWHJTHq24FQ/TC9nUVXs9zMfSmmTEHriHrCp0QvjgDjLKuZOtfJ+vKdJR
XSZpmLGi8uj0Ed4tA97XW2ySZgRp7ksONObaQRsTx5yFXjbsBc6K232IjEsHar6KM0xNTkIuGqYr
SfSUF5bVmZcPXLxOJEEzzI27pSWpe7ikFsCiK3mRwpLqk7R6cg1ZA8I4xY+BdmL4c++XWZ/+Ujgh
DXHhMjI3+xxEWaVvCQJaybg/TNOHQ4WCU5wj7BjRqbON4GkrnLcE0PRticgIAOIlWECcmDhU9Nz5
bGaHug7gYxOz5M4mbujGTMu8SLwzWP4EDN3CxbqJpy16zMNNYriqOnUA0ZIs0eAHKGUt2yLj81VP
+DaDNc2u0s+pRrGC//pLzbb52yqPWaJYmV7X9sPRmpEHbf7l7xriAMD3cJMYxSrN1RzDzt6HVqVA
l5MltxuENKXf1wBr2Fz8ORDNBSPj4cad2LPlppGunLHtEAm4meJ8CgunwrJkbC+WcT+11Ax2pFjC
ncUWHsp4teFDb2kAVXvo3EGEkqA33uiICdx5fajjcZmCOU7E8mgGf9ApRTNEDkOaOUu1cBihqg+h
CnJvolRx7/Zw/Bkd63kpUWM/b9+QS5g7Gn80q3vvxRyBm213sDpkM1X9LwW8UYXlXNV6c1l1KgLX
R0D4No44vZu3G2whcn53943m21lkFjFjxPf6QPBsdE5LaB3ZjW9kkAdLsYP6VgWAIyyzq7VF4crS
syzBeC3fYGE9Ly8bd4GbVfyR/c8JD2MF4unLZCYlOeC8PgbNJ4TJl6y3C77t8Jwd11ikPzdrKfmr
NnOGYnlge7TLQpt+mocCDR4n490Hm51UVoL/bksWQ/OuYVWNvohnv7VshnU1xRLiq71dLRSVdTH3
Kg0Ta2xtltfQYfadGrum7zFS3kBky0rT2BZCFUAAWkZl5ymVKEYBygTsyc1lOsUv6cp/HXZyp9Y7
0tczNHZOHrqLMxBeadWThrHzb4C6H8d5drZyGKzax0cH0tyq9YHlTRiJI7FEev+BArGqgcNUO+9u
RR/LPWJ1VQyIB2bTQ3MurRJtqPxygsyJ2DbDDaZuhpvACLrIxYSWfaZoBXmg5jmB/uQZCev2A10U
a3Y0WcKiGS0dMoCbPDDBkpfLudvWjRbYdOv5JarWQx0ZwHooBDBSCDj8aneorqU1skoN70J/OsJ9
pvAMCLN8JzVYbtrj2qg2q8vhQRxjyaDUiF9IqlO5MZlB8gCK13XuEE5h/hwb9i1F4GE9VQsoI1a+
JjQe8u1C1UW9BEIS+WH8CXuD7HOPyxzJzIDariYtM9ccSx6nZ06Q2AM0ofvFU3032qrb3bisvv3h
9BjdjLQeKG8qBswyYszcr2MyTPCi+brfnibawYkPphdCQaRaeKpub+FU2IFTkZtsVmDLsrekZzgW
f+n+sWt89jsY3jICT/clylC07n8CIVWELuIVhnN3mLIVtEc4EJdfGomk92SYviIHpsFj/lcZkyZI
D5FvppSB10AAjRAD3xHHKBU4T3BtZZZI8TD1wZ/exSsVMoFBzD8oRd6Vkej5LijIhDxiBXmQcLt7
Wc0l89/HQi3Vuig9czNWvfLqdPUeJXpZOvyeVL5Ff8eATOFaAJ/FqfpP3PvdrXrM1XSgF9dBHHyw
i/aH+0FMBg2B7AXgU8GdwLSzcQ0SiNLeNa2FLnq6VUUnhUSUFKpPVm3FcceFUh+78se1+2XyZ8TE
3IxWAo+taHCjZFynkjsuJYhLootSqVQLiFqyMtw7K+OfUt74OgtwiAXrgcB+9HzkJDeKs94Mb4td
8mgH6pGsu8bqx6/S93rn5lIzbFD9ShxpXCNR3hzhB3TVc4U+T1X9Lw06eN6Go57QPrpZP62p/+xY
IiWTSsU/1nDeSVKz3Y/jjmwbIPESEkP/Ia6e9CnpSGFaO8ixKGf3ti8p329rkea4kfIIP4xrg/Vo
dlWlNJlXk0pug789dbNLZ5Pc05H/JIG8nX/Z5g0ckEfVIhKO84i7WnA+m/tIEXgqv35Y6Coq3+zo
ISqXkniPBhfNR9f49ny9I/ihFJbGfKKaT9Xb1E9rQOCh8cVTxLi6DiaCX9LMe6p4VglbGpMrDAJs
c+FFH4H5Z/kBqV+Gu36uBfi0u0rakiKgujNefRd99IWEfBcOUneuv9F4iSD1FLm2ZpKDCtDUpbE/
XkqSMS2O4Dcu7wOxgvUkTNCI2kW4LM7fD1qeMwgppdhk+HvB8/r7GBMnRKg1bAvm3ITMt/jR6iUl
gVspO3qbXOtT+PgsxCoo6x2T1bNOsJVlBc9trjf/CE4dhdNlsjWul04ZFQRAEi6u9PK0SDb8y06r
hWmzZkcAbt+2WWuPQ3gAR6qp0jZzlbtefaLGKLL1/SebD7EWFUDZW2LxVVxDWn20+hvXD7pHiBR9
LKjTY0VYblcm0ZLHHhxBK8Oo8Wrnf5ZIUmanWy8ezma2rWY9oXlHxuHFknEhX3xIz5zZITcQ0Erz
UlAV26fZKl+owwzCohR0NPpWnDfwb1yzRpoEY/YREQ7mPezP+Ar5c+kisvd/f6eKGv6HlT6fpIEo
77ZkS0fnwaUjBnxEZ/zEYkGBXDbFTYlX/wj5O/iqhCbdgpTpgE3bKyQ4M9ItMsMp17EJgDCyIiMY
CiPJr6tCX8NHckKDYEYEZw5cxMPcpSa+BOXgMP7tVGDJMEb+9rspgB7NavVIkGNbcZ0JmGB3KFVj
vUXKLTM9L5HU8f7UInTLQ+Bn4RgtIfnQY+OkqUzxEULwccejnyZ2nC7GvthiItw9FmIC9XBw1J3b
jxkL+lWl/LcmRdmjZE6xGfQoz0PJWV/SNWVqxMeCVHIfp+GUYZ0gqUmU+K3KmkIxMXT/dAXiZmyN
iNIERKksOQoFImRQyw7iaCoW2D0oFf7QxzvaoonkW/Xuxol8m72yj3+BHU3TlAf/1C4R0ikg6DLw
oW3ulUi+6KIaZ7h9Oa+I4rd92O0BpbJpuO/mD845Ce0BJi8+qKu6014Z45UZFHEO7Pb0IpxFyE5Z
aOx4PYNkjBwunijDBsh4x2tw1U2w6RXDSsYLaGoHOrHA5M5dzESqA4KHVpUArCbWlvYFIAJlRAUl
bnA/xk+J/D/kPwDTaryyWskNyGkHIN5Xq0CtX2KRVMLGrtXvbbjW3jZjgoQPm2zi/Gdaeq8au8ms
RH54qDEFMI+K0SZTd/xpv/1UZzMFHBfRkttTETM25ssupwXq7sa3YG+li0PtAwCsplkXkAq6ylIB
pm5mdnIDpNqmM9kRiUUuSg39xveBUlHwsHuD7qDBMWig02TM6QN8T9klDrtVNAlK3U7KWVMtiD+S
tflaglcWT+pxJ3PsWUiIM2xOINzm4Px+IXex1bLorK6Bucp5Kht9k4DzuFfGb2gthKHLi92S8uqc
5xdqjF+PrzqcEPUbFT2VI6REsRRznIzH2BRbakoMNeRpUow0xQ4RMXHv47VqeC7f4ygwFj6ppVAf
oelzN4sdIAi66TFsspzuNHe76xiv4blQiGJiJy1r1a6Nd8ePUddI2H2nSC+uXPUVzWmrKI0tjiYA
Zohgq1rHrqvcp86Nr47j6ggFL45mekvtQooLQ4Deojnhz2F0UWRcTE8oZiXNVZmItPN5ez+ivy+w
3RKwd1iWhj/VbxBj1Ck6QXTZ+AtR/xQpG0OX0DOl45kEPcQEkAo4CirhkhmiKkZIsWO0oU3hMyQv
h+Pq1/FqBkxGSClKIb6FrWPSgOjhC01xYa2OAwR+x9qqDOVOlJ+0uIAk4ZtYSnYhwQKxmI5w/SLD
pLJJooemYGv0IEICGV0JyKpmw/M6nfnccABRYcDCwchvMYfJBw+IEomXwLWUuWfpksHZBxUdkjO5
KLwwoBw7M4FD8cO5BMkChV6tw6THg8079rS8F43Do1GT1/FwiNav4s24b3PsgQx3TaFwywDuTf+o
EmmcQMh1aIIPMUZRNB2D8hHkauh314z+5MxuGqYK04rHFnyACDG4oEl9mhZ8kiF1l1o5A0ayIec5
6C6azTzsEaYRlLHsK0bo9eDmCejZFAlhB7QDJLD6Z95befFe3JgeRH/xWkp3Dru8VujS0SJ5VcQ9
SHEjsfgXuL0lNimyw/Fxk/TTQC2s+vHHrs/Y4tMU6TmEE/65jeUFC53Uivs0ga24LJFKUVnwa13i
d7EFl9dQC26Y+WS/j8HmohHmULNIyl9JdiY9pRo+kHWy8PVU9qqpkIjXaNToVbcM4ntkUk9f5Y70
44yJY+MtTaqtG/byURtg3PgtNJqMTTuZ6I2JTOVEHmM4FbNXkRi0L+Bi5wAge9tr2aA0+urBKjdv
a4KLQJMv5bnrZQSa6ibonGLz3dZIR7IVt2INvTWPem4wqSWN0HaOAk386IioI/gElxGQ/Ux+N9Eb
iFctD3z18gpdVTFzfRCDc1I6FLOtgoRnCw2crwSOZeXNQjJkF0XmbUJdTeL++xJWoEYSlQGiervT
phVOrO7I1Vp6PcVylUPS5Mf3QWZD4VOVu1wojW/rrKiOHVRpA17xmiwHiZJ+MGdMpAa3nPTVpMmJ
IsPK5Tzyntg2+aDyeJNgGz/S22D5cPnFb4R44U50fVTxr/lL3Ifk7i6YGS2GHZoM1upurwXayJYv
CwZZajkynA36zjR/qwXLpoSrWKHdFm2T6sPotkjlFtqSncpLAhXuUoZ66pjaXnkOkxNkGTxE6fZJ
Ezlg7oOJojrrCx1ueqy2Ggo3FPeaLp/Z81HRpmSOSxidxl9SAfcd7ltHOxZtLDj26S0M6DWlacqD
08onQ8ZwWJxYcfmjkxzJ8ZjD/cKfskRZNuccmg6Dkn0zcp02m1Z5RqsAjEY6EpKn5KLGcVHFHmXo
lQVNgPMx5q+R868u251W9gmfSlw6i3Z3Y5Snqva6MR69N347iKOTjppLGbNhubYn5WHdsSD/pUDM
PRvPUvayv5PND3oRVoHfLzp8YAlhWbvQNYO5AUO8IE3ngcT5gGFj9gIecw/XXQxxV7d5YyIq2mos
iNm+AleuU8EI9m6vwwB4NeS3ZA4TuLn9UXwcKJb6h4bko2CAy81woFAg/SCglFErzQTzy6bv1XLP
plw/NOt+gbnUPpDjUHORKzIvAxZMVzbgVWWv7AKgajJ+OiaEvJ4EWhu0duSV8Xpxz746ZIOyYJai
PeW7Hkr7NIsJQLkq4znvWXzAI1EcWgGjY1i3pafgLsdF99y4Wm4HeVSz5Syq5iTyUHbuB4Xov7mH
O3MIApPa1ZRCQwAcXaZOSDFm1pGGUC9867txEcqPYCfJQw2IW8LyNZQ0WVpULgD/W3CQj9hbjoa0
PgFZH9VgplU4UWuony6AirZ72vIJFo5ESaXDNZyXIHQgNvbTXSVrcVClcg5pShUnIfIXpZkCNeaM
f/3+H5sNIyVNCRktOehPlwCcMZ63FOw2/cKFCxRmT/c6DMeJBTMzCYYyVQr3C3np585R47yR907z
0Sg9u/gJjoiEbk82//myKPtHW6J/k1pktJxiXTiDWTg+aURg9mLB1cqObAeDs6pknxIHOwjhPloP
HfNnXJ9L0rqMUGgaXnqM8EQKz4v93us6vQZyFHPxiAogC/1Sxl5u+o0+pYD5unRbdfesiYP5d9qT
PCrjVPqArGes9cBIlEB/go+WEbfAAa7VZttU9nlLte2GzphJ6QLcCOgcqZvEEDySonVUSuRvnB5F
UbKgBpd5PqUakbYs9Cmf0ErECuBxOMN4AQLmyzZbXfJA1fUVqLtKysdFSU67zswSgyc8HMTmu9sd
UYF0HVYVvvO2jg9CP08Ch9u+UcY9sL5eNOIYu0yuwkxek7u4dSuxU1AFb1VQmQ/J4f2/EpKTzqrL
+Fu9NfiN14bvF8TERoY2NxXMVkaNKWgQ57ioIPJYVCovzau73rm0f9u8WV4InwV3GFhGo1RKhEUp
iQavmgaqyyuT4pEDw+30V4rGd21PdWWwULKzw+t4dyxZ7ntodiwK6KZwiYff6nu6awYIsTmj8+zu
EnGB5llb/H9Mb17MwbSN4I71gILEqd7cmhoL8qNfg3GJr9FHvhdUwHviFVqN5lz++yfoi4hYvrPf
AJMIFNhHdpTsXdadZUdOmPtf+FAM/IaIaSNTeGXK3EomuUcgd38usieKn772EEf+KHDEJA3jNxRu
AHbf3LMRm+4Bz02wzZy9ZYIPkGlzMXiG0CyKhEgmv/ekrzxLcHy3aMLAhNajnMUZIvDqQZwjslEO
Vc8fADSHTTBjTus6Yz1Msz25zWxVOuyhFYIJPK+i3SVsBj3WhHYjMa17KUNdqGTp9UysOewAE+N/
xEdGykWbX4sqvfa4gRbFHQj/bYxLsRw2z0sXvKykMiRas54VNkisrw9YfRkWlDtLyCwOGeDvGip7
daxA76Sy11GssjksEvadaz161Dcx6v8bGtLHwqP7wTRfFf1hbCI5hOKnZAhuqFZNy0PV5sQA0z85
SdS7/Yq5ugYJB9tQrM7YPPW4Edb6ubGRrjt5T97GMQ2ECH4KPxIBJ4VnZwkpCkB1cyEEJA65un2X
UJtxLiF+iqDpY/XpnjubvqbUGTJoQA2EGv4e6sJYZKor0IZVcUtRyXP0TGgSbzr63ZEoQJXqy5UQ
DnJ+3LXMQSSWmSsEq0vd2cAFNn+0xXKz1uJcIyDWB+EduQlsFhij0ddy8V+raJITD66/dRt0Ssed
kkroyCHLRBbOlnWMyp6A/dXUcn4/++URFy7k7As5oKzXE7Q4XdIoEmPt1jxUslqE+BsTwE7Zslbs
vdvikQGpWJslMhdBUr8hLO2TDyCJX6NbwsyB44SknJaRZNpytSFyqHVCiqq9LMw/U39DYsuZYFWw
OQjzozc9hs9l5bCJYPqaphSc0aEYIFJaO9nTUdfqfI1N7BDLYpkCCcJa1IXPyobzpen/Fho+up1l
grgreda2gwn0OKACDJVDujga8EhVeKRsB+AzWNDbqNx/r3kk7Wfrh1M7vMJNMQcopdy7FlauCkgk
DOXosGQL3FrcnjPN9Z6UoHBZKeZo+If9nEPw/rKVZAJv1YlcEKtnwAPTPK789X71D9i/tyOeVwaW
mz3BhYa6MKEprt8HMJufVVJ0irj6vyls3JGiV1KGtvVxGl4jhVC9J1TzBqaKP6eh/KT+dghCiqBR
F3XXwfs7ceTcUP5wIlaLukiPfIgYe3tgvIK4+pKg+odbXk05My/aRwim7VM1A+FYvUODXOCr/SSq
04h2e7bk7LaqpPC+ER/6T/ZE5zT8WZr/JTQnfVh+S0vStxbH2cbliOdvBpKooKZzyRfoB1W6ftHn
iW+VcN9+TAjxS89d95OZDJYAkCfJSEGVTHnN62wdwhny2crtP0LNW/f1dr4iG+3QQlXZcq6yJDnp
ep14WSSiMHRcCPo9pBzqKLpIEmnKreqVfub9qMnqX0cgs4RgkRWqelAkQqgBRKXJouRVsLNS5I7i
D6eZZhQ7qdmkzK+M26aSyUHxWM4gQnwIhFsLh0fKjD5F3BYzJnpGXfl09aI5Azv2wybmTBJqBVm4
R3NN4FZL1gWY11F2YJ1gPYRaEj7xuXg7eT3fEnd1RGXu3vxCAmt3/6xmZDxR7qRTSMopI6N17x9R
87J/MOef2/6yYQ+DOVyzXtBdWbWrWWu3R5XLNzFJCdz5a3ZuT7QqvHST2Hv2NAVJjfQQCqebfFVm
XO+TUTE4jAPwiDgRGXQRZQa5y/fxrJJVZvvn78MRUuxqi1SPR2zK7VvppHoj6QM0RS1wzq1fNDy+
65gojiD/qu3w5FIgjSRxG1r0pI1La1VbJVs7DOiPKu7ZsnKbCDfUxyNRb7e13HcuKWS13P4iLpPq
wwidLrcrYZHOMi3FhpcodY8oNhXRGMowHIqCbueAOx+KPRGmDzPDkrwOotSHSWVYr9GBme8QA3MU
7bsZ832mXt7KKRF+wSw5MnCUkM9FVW2OidLRQnta56+2epr9hyVHvebC1GQ/q0uV2lWlCCs/2IJQ
zMNkCtIz0L/tbrfMV33T8CfRTX+2Le8liDjSFGW6bEsscanU/HXqKAimozCzZYxHNbh9BreIo9w3
EaM6HUTy91ChS72MKRFy7/WkKZY6fvUXE+5GIH3gDxJeimAik5XO6F7R4aP4odtTRtUrCRlTcXTq
qeEGM+UevbcveGDyb0LzI23l7BmCYBjIIdVf/PktZsnlha4CUfKVB031QCKlURB6iXYr+zGPg7uH
WVH+Mu6aCUQ4clHzh1/kWvHwm7RdyDuuwgGsDjRPME2Op6ssm12HB9XmuUWCRbZwH25d+HJxSzhq
Hq9Tdy8H2EjaNrmgvpj+ezbd3uYMv9xEwx8tXmg7RmqzWvXoVP5D66bnEsHbwUxeCjmJwvKKe/QE
7vCMMPwHI/HdXrhmcQIrv/pV2bvbpPycYD54AuuDug7pIsIwB96SjknK52UxPOJ6YAo8gk3kgjaw
pyYM3LY6ajtX6Du1JnRi6BTvCSRH7d2GS6IDNKscHmKk/w8HOSjY/mnx9viQFx7CEv0XUUOtEBTi
mtCWkDkT78LxJi1JNt2S0Phm3GBKrujCFqusqwCzSxmYDl7lcbdLUcNFKlYfM2IwdzIBBj/5cWvb
5CVK+o7g3B3uN6YGQJraaqo+tgsgimCoASPBn+7g8qhj6oquSKM2fTRtdPR1d7RkmHGbieteZc3x
LBZlZAUms1+YoQfkPGNp5v/Qa7vxmdgsf6GV73abR2PrVOEyf1diTJwo6656YOmMTTGjVRleqawW
RsXPwI835dysQ2YJSrd7FSvWLGBFrWQIOA47ybhGI9OJIT+Yfv25UgGlETRBEF0zpVSOYM0PlJDN
BeAPPkzdNSoUm+iaOPelFvia2JMTcQe57ma73ypj8S4EEd/GTQ3XkgVWr8f3zs3L9UVwAt6NcnZq
VSkXKBNiaiZvyb7EpYMDZKFcVOZqgdKf/CkvZuHEWxMUn4jHLZdNZyo0cFOKEBJ7JsoDn75KxW2U
p3XnTA4pFGjrIoLbQkVMHizxCsi5aV6aAb2eWhYFsHM0q9KgmSxdCnJshASSJ91B32FsljfkDUrw
AnNSdyt6j6bnar8kKenssE9EY85uQmS9NxRNKC5vy0iPTy2CVnzHO7Vqx7FQb3CH8aSEPSxqcEy8
M0pD/ETK3I23VLt5zJOf5zsoNqBg5zAp1bAffaHpzufgTjJLDKDoqE7c/9+xJesUJXcmwIPhNqih
/iPlsSJCoChkmhixTlEiGNaerIF/tpotJdgOrL40k5rInHpU9yXTSE9lkuBQ0L1bm3IDGdFFaPQv
muYsQQg1Oh7wxKtI8BMp5wXvuaFD0iApIT6ts6n+60UDxgT/TEbpY2z6wV7S9azXj4vplswC1FBE
UVbnE7hUe5K3C0CFIjEwUHwON+5/qwoX46xPeX+pnkC3Z+bkO7VFlVzBJvXynDyrD5r/vGgJqSJX
WWcCE3OK5c2Ly5ZD0DQPu5IIuYIr/bfG/Dd1C7/WrAUyJ8kNaJC1A6edzOHEqOoHWNUSZ/fcKdTB
S5ivNYc7yzG9By4rU4vX7Z9tT6ME5Y3J69jS/g2BAyNGT4kQd/mz70eElnMGJZB401Xh+w+v+PI4
cMag/sKDRREoDgtyeYj8b7qn9HR2JMxkj0hcGnk7YmZV49uqZqe4Sh45NaXkWgxpyH+0xg07qZS8
99vl1tvYjfDmg9JrivfOfr9V0FeJRNIDKKw7hObY89HTR3hMzPzlrmr4ybn32hdpLxlklSZAIiU8
jFOMkgQlYwZcTGgb5dgjfEplpB0DYtnEJm1gw2yYV398cyZf4NGHb/2LQ4oJNDQenCacXFrtUTeP
SWo/CpByUm4p/kcYJocenpcMl9fddAldTl4UdQI5TL+Ha2L6GXv9ze1N3oJW60CL3waKkUMZ1z1M
yv24E6h2y1DkQ2y20ZyS6W38n+mXJRepfWsXB8h9WqEPzbqtLY0OGmW6dMiLklT3rH3mfuCJvUhE
pavWATg3nP9zauExW0YdWSWbua8liyQnhomRUtZ9lJM4PuH9TFwOPZm6+zYZvIX6RIddVM1R8P9H
Mh1ambGmdMcSmG5OA95hzzEuPsEGn5oXKjAZwKLj51asLMzA2bQ5bUINQKHJnE4e6y17nek6qDOA
pCojo3y9oArZfpcBKFAFU0gIm2R6OvGRaZkxjfbf5+ASuL+kh0suBz4zis4euwAtJiUEEGKLsiEz
Td59vnIKAhPClDTZ4B/1kfiLekiFvRCjKoPMEMaMaDCNMohK3NwndG57TDZj9UW9XaGp9HgbCEvq
ArYB+pP1oJJResGNteokxXsvbXRORi3ougZ7FvCwKfjzSKXgvNTJyiKhScwPGAEoVR+LY8AzmFU1
bVwZYs7LDwoOjBIuuHLXxkto39NmkEatnmSzr+z7ud0SZQex1MhnHma/N+9jO8KMuTF8zowuPtzz
03JzN6RAxUSJPbkM1hLOFijoOUMfyPa7V3Y+pF+n3Bc6gFqJIPggET6Wqd6JGksYZEGQS1fTQO8H
SVAolkWceU1UfRvWCnuUB61J4vo+QFCVeo9SsN9eUjZZWruSD0iphku2HHQc5Z5eYZWZXtBvqXcw
sfMcRL746v+yIpRik8j2DkMmY6RghuyzySUcAspsfbPvmdVbGCrIcz3Mog7KyQRc/X+29i0gJmOG
9c5HFRG2vd96yfTC6mQUZD/64eFEw6U7G69Cxp6xXscuGD+KlvYZtdEamifgkaZXQkXHUz++QZmf
DMBRTpY8HIsZwkU7Hy1EiPnS7ZrMjwA6FHDNUhCd30OSfn52j+twZdzEvL9GsxaIgqMFofRowAeM
xfkziIHxZh7Gq97XTEqUgHdO0nzpkX4GJkNifdsE+l7sBbLFjLd6Cufw2SZ9gZePMfe0Br0fS0cL
VkVnXUPGHOFoOvork5aBBqhzelf7Cne+KbFo/jFEHQW85yHpTVyRmKr1Hb+4JSlk/B3foX+gRNdZ
pYyl5OIuthXAZq9GwK2z1qnsavOes+O8hQigYGo9ZDZuHeCvi2x1CRR2CTBwB2Ze3br9BbopLaLc
CtA69wWCHycggrFs66DmWB9PB1cbVjpy4RcUbv+2bAPNFKh+Aw0ooUXa0pSaUEfNGaHfJlyiVyuS
T7JUCQVWWZBDUU+PlEoDeGa8jJMmflrOYuEeHlpG0rfTzYvU/Q8Y0XpN/lYqklZhCMnZI9LlEtg+
62VwOP7MNlhMU2ho5yKjvS/MlP/8y9NtauQK+amJgqbkfRrCjuyzHRdoOphPWRgeAjIeC8eYOJ4e
Qp+Ny1aCMyIggbuv4n0nib1mAdQlSWe77w0vIIneNBPg1x4XM/BnZDAUG4PEZYLXVdik5eq6kTEr
v+qKIrxArxSR7Xid+7T1tAMAqsa720wYoMQsVmlmQOGXMef3C31aqyRYwcsBDKxpO94yEnv2oTvx
hRg8aKQRDpOpgXtdOLerO4dGQPo6bbBedeCePCuOQ7ch+EqfoAjfqHFEeor7H0TfaBK/1G0PuwDl
rHHg3lkxWYCEK2ur0l3L35GWPtkzOS6OaRETifg5/ZIbp+8hypCYDErGAWCj9+6MmmHmovfP7W3W
kxBMohyRiVtdQw1siYKZt1EiSTDv38YXmPtCClHRetgKSEkpslMXwoWwS02G08GUQITAPZxLx7Ri
4csrPRMBhWpzdyOeFovHfzifO5HmSUlK/mFabLrLZyrXpr9N51I0SyBFzbtBNdpxQtesfSu6Ma3i
F4OXtRl1dIfKthol5dXcBOoHHmvvo9fsDZFyPl0hn6nKa4Z1cmJctdCEWo83P4tBgeO2hSRefDS+
ZF/phMmM61YWpYyjnolSBVGClwn6E1kiFiodK0NaMFeAlrcgxyUpuSsKhh6vHYxb3FofL5as/moD
QFsXzD/VQXhQ9+hCkRX1BGC3LmKVm6/QG/ydWgMEWKK6S+w4wmExFtrhaHnrKIKSBkuo0VK1aYVS
2gw4vT4YaB9xB5BrWwAuIDqkFx2D7uGYaIg6th20pTQ5b00A6ux9uLF7dUyeW/kA0kR1ePSgWCgf
FNcRgjjw0Rgj/ndCP7ZrdZAKa6BWyQ1ghBWI4xePaxrOUhUPj8kJbf6m43fFXO0brG/gsev08hvM
3oDVr+0te/BcAN09CXg6dZPKNK+DZQSu2Gi9PGCfYSoABy/tp1383o8GzAYgMRPKw/q2Ge7V07ZJ
9ciYz+GLy4tUbeBmNGz8tntbGN5kNsdHGIIYFEGDEje+rvaUVgXCh1cf2kJ218cVJyRYrPhML9ef
pSMfW/dsvNGC2Tm8ULWPJkQyMQgJF8e4KYMlx2x6QATeoPLeIVmPKzgs7jYQdE7vGgVnTaVkLgls
CR8Y0cchpqLPnmOnkmy2+oCJq2IwSVBbArFutQy0TUxL/MXzakQnHF5yMBF/4SQDa+MUL0C/PB+Y
VhT3K7Pa90AkI2VwzWhS9w/vr5PSYCPyq2JgcnNrkqy2lPnv9Bv8F9mntHMQUKBhR/0Ub94/HsVv
nbMEQB/GiyxaIpsHgDy5lbETUFYcg6hyFsKGWs9fw75U/U0siyXCgCd0sCH1ElfGH+Y1l2IifVBu
t7ZO7ThLGSpaHmE6ZgMJd7j4OHTcMdLxDKkjT/Gy0fARyarhSukyn0/4R9HV9Vn1LKyT2FNdfLUM
n0LcnLiTToDO68FNtqP+Ve9AiV9ibcyXt7eCQfaGCzPDy2DE+uaFs6bTFNtKtKvUU9qPt3fPe+yj
1E6OP5mgHTfNEP3pgOCw95rcsiyjgOUDx3rBpqjBppF5ZWOfgv0sEJKNsIKoDkFowSivtdw8aDLy
T5wTUtsIUV77xKwkRsp1XG4Q98babhMQsw5s0G8ZubdCUL6rHLDPDpfJxUBI7sU+fc/P1l5mfaDk
mIZQ7xNxTNSJ2W8Fek6CQFZnxDYJvuBETz9/gvKN42JkkXmnBo+C3y5pI2etOLHoLDVLZiitbDwY
qcHYH1mAlR/Ypq3nUtB3DdFm1tlLg1p8/iqTFrApq3rlrY8WAIjrjCYBEEopCM1a8ZBI3Cii7LsE
SI8vMRxGblC+VmOSGiBsQpjGlYb+qlUltA68t2qHYh/KphK6uLCV0OzLZSA5CNTnHpeHXj+RlLJc
mG5tDC/zZqV2utM52OWcr+Eyp6+S3HQxIFkigfk+6GHNRdNGEXz7VqA6i7xyyGZ6JY+wrenUn9W8
mlXP7VWjYKlsTsDrJUd1mKVJujPT6Es8db+Si1fVGTLuEVvf3y3KGtTVrDphriABnt5VamNf46G+
uKDgf49w0RxxYP2j6A7q+fS9rrg8FhLAD/RamGL9X2SbZM0YXYxCmPyOUGaFnUTKTLu8GIjmIIg/
pvtsRz1MYNafwCl4eKCbc4MmqaYJihOUSKgr3Cop07UdMZ5LTgl6xmsDqCmhnqMZimqXhJXnAhU5
q3owzd8iOHC9qITsDAYRwAqtLDPqKvMAWeYOMGd0qkUYzqc0vRDE6IAZzUFCCP6MdKOqmDmE2SCn
owsW6CcLTqgGonzrX6Ct1pl8LLlCn+PeyENypTMP4PR2DCCSTXkAUhYidzNu1vbD/d7ES06Bd+gj
9RpzmO+690x9AnT78sNWGVZ8MiTWYla+PeXganpq5En3lSuaWytA2bxAr4Fe4YMTXY6YDAEgUqZS
X69EkBux0DyvYIZeEMQACoT6detKRIhiBovkNm0ifZ475EZqP1cn6/sQvin/JBIKWcWbh37CG4hW
BNSLBUnIF4bsy+77BTwhVWJvauQFn6U9TlyMrdAlbqCtMCbkRCTL20fUlhHAjTff6rGeEfqTbuVt
oK5WrVnWvj0xxIN8CvEqYLpTzx1yFZdJXBWjEd1AsUV+XEBPFqQmZtwWnT3cgLcCwTDbOQRtDOI4
spBIz2cIB1O0+pfZ7RVC+iTEr6U73nI7VOib0laB3eIPzWuDa7o68bGZGdjTqe3+gqgy+7urB8rn
2qeEW8Nr0U7zDM+SDkOc1NxppoHlO8dQKuZE0DGegjbSe+klSmXV3+nJQkqPonCIKvNRkBoeYWua
aqk2ljXWU1Kvq0kCYKR7Fq2rhLDdFoaJ5fx8PjsCs4HomIDL6fTXn0EelD56fCpIMPZfUbFCm2Ai
xyiKd4JnupcvlQ3Mf2ZDxwDSaj6Q2IUdZPYlmVUAfqd+GtlchNSSApjGQGRRicrTxG+qlNwtZJuF
1hnzzRYLhydrsVOrn55Z/yAbbdy+7anvRvwBn28nVhot158/jCxlws5wbABG5qkwqEC9N4Cm2osD
jJNYTxomIDBK1W4dbdDHYrLBxJBpRd1wrPaYXDa3C1sObPXwWpP5ATUR3BLRx/u9OGrBFIVWKJwg
NQx5M/PLM6NMxNj4732OFMVQ3ZgFPr67Fhir3vWtTrF92ePzZJrgfRJ1Ycz4N1hmJPdJ/OdKtNni
owajFGcFQUBFWE7plheY3RPeErWiaj2TsBbRUHfaqdBRx6BHPHmE2EZdeLh2OeB4T5L1dRs8zKq3
cmaZaSTOHe8pczaUUS76Zc1oQ3yXGMaqlgPWpwO/tk1VvOuZ+6Cb3ixovCihzOMcMhUTBQYuhLdg
C9KLgwrKyrhuvMwOXw5rRvygd8ftd2lj9+CgmaQsOPzBr5s9QJUClCXN36Y/1bnmEapMKj1YdMC7
B2/BpBVUKeT0zuFzJXxKv8wN5dsPQFbt1DEnVAbpsSZ4LRVmGN7E9zJ11w0KUyzv5dv7x9vk2hIB
ap1aK2frNCKQ5Q+FD3pZzekGLAFQSfvcu2lxn1kK//caYBMLlutXotVpwUoRfD2Nck2kARXpmEqf
VxEI8IdShZsRqxtnecHwTG9m1pgDZqZQI/t4uBQSrmdrdfXbtH/whXa+kobx1GINNc1B7SnrxO2D
EM38U9SZ+ZeM0ugVDUcIwLWZugHovaKCvmx3hSd2fVLEyQOJ/Ku2yUFZLZKqfwX4ncHtapAYVOMx
29siEw8oaTl0I/ZJ9YFNB8ysP4h5mAu7v5t9RDumOF3bkUeb3951aBSZIDOo310QiX4fI93hS5pc
Uh2rH9xWHOwCo3A8J/TQwlZNkQouNBZYroL+Bo7l98vX+lIedOwNQLIwMU1iJeO7ndJ9X/6NGnQW
fgxBaV9jX9LI2EWB3Y7e8fYxCebhBZ0bQMDMaGvMm9skMgAdsXpmmxv3u+x8ElYNJSDhGfALoTZN
31DCVeUlGXTa4wB/mCZfst5A6HHQO65vGuAlbyVJFSM3JfevaI663lBDc+88XvGVfZtsDYKPU2yl
v0Vy2gA9MjxXoIGBiisPizToZZsE5QD+2rLXmj2J+jYFiImzz9PztAyc3znaXMui+ayK6h9s2snp
CE5nwyzDNB2eXT1g2Hy7QRrF+o4OfTmK7MPNKw4F5WKlpgoldRLct2K6rE8TsLVHMaSKatDTq1eo
7eO2IW9zZ9bKUeomspWJPLgTaRyzUBAaSoLPX/HiRNToVd+1nZctozyK/nGKL8IBbeCz82qZnXGy
mCXbrvu/jtJYRzeJfWWq4YdhDf8tTLrueFZKj6IyNxWPS86XAsshQNfAEB91/ximvOEqMtnUjidj
VJuPymvyBGkmOs0luFdL2wElMgjrcWHxMrom4cPFMxJe8u3Iop5Lr2HAoPGBRyXcqcHF7Anvy9cI
I/BkCMNkZQdgGGeub5incKOlU+XNNKoPTMfCMkEjbHtS+ohyR8CC0UopSoxni5uBmablj82W66jX
fTzgDLQ4aD4KXqxzzO7nlRBuARF+IPgk2e+214tkAFPHFYbOvzcyxj9M92lfNM8sS/xjHNt2cAa5
HM1RnvvMKzgzHrtG7bop1hXeP+LMEfX0kRz+gFUiFMiKzqLppPMy9YDNM9AzduvwM1qf3MOUWX2u
ZJC16TA1H+vv6REVBPjPCaNBssiyyWaHXzyfyTpAo4WgkF+6B01nw6mXKGeGi5PAP2esRU9lB/Ir
SEj5LjpJ6pMdBoEfsDnLFL3CXHhClvtlz8W+mcMzu4AVUwTl3R5SgYz2Rn54GO2VEEvrhkq0yvH/
D0u7TUaTy3i6DOxqry7Mn4c8mYvUnvnTQJ9zQ9SmzPLYxOpQashkw8yilgDXRlo60vdL6s114DrK
a+V4tko6uR6MX4rft1Afmv0hQ+/kYaZVJkjYNJSOHRlmrF+ruCXIViQidmFWb6fB77LOLjQFal0G
eIea+usgxr5SZiq5QmS6BMyssOoESTcQ3YpnLpgrxH1pNvzkGXgYpYkIihKxVxKOGoRVb+gN6wNz
BL6JV9FHT/lu1HCoj5bhCggkw8wEeuD/Faj/UJ+khKkgZSHxVR6ONON0yrWQ2uFQUBdsLznMGs0b
/NU02CWxnizygeASJCbv9DpuEfw1lsmYXCGDCUqVDgn9NExNyLkIIkMml5RPu5w//uThJXyAUQ5i
osFlikdz/VrRU2WaltQbJEAvsZlt7R+sDiYnwyRO6lW65EKPUARasmFTHDhk11QME7yzoDN5IV/V
27M0QNrHwBYqqvULKuNJAxuqrRNd3EaWwP0EakxQQICes+4dze4SaehdOLfyA814oeHSydVMcRpp
dmcy1xnGht//cu5lFH9Yzb89Jx1/ySkxF4v0zOKR1R8upmeM3ygHZKreyyhrKSKAPW1fVzzMT3CU
DXUeBwM27PNLTLH8j20b5xGXYollsBpj9+e4yIJ3bKWyKhYgljhDL2b5u7KtMOqK0/+jmG0Z5rHQ
s1OwVSX75MSXJ+h2v173R2yyCj2Es5vPuBgeXcoYc5np+784BIBlegpyIspSBdGPtqSyRWVtOheV
KPtetpfjVuasmxQYyUrrHD0TqzEm8opFC3DqDbI9ExTLFK6PpqNod+OoZEiB7qj2zLQrRP/19VMe
n6NbP4emNECPsI9vuoNA/vyJ1mh3P/8Ka4xooBNtBoPG9Fa0guUHW5PHglHwH7kF7SheSMDZZzWv
BSUxpYZpIIwR6CbRa3fgMjdRsIPi8mZP5ORB93ShxPmjsDG5/60IXdUVW0l/5Vd0F6BOD5Tx8oad
tBRUHeyFVCQ/L2e9rLpcZr+8lK+jKp0kvXe8Tmo3CRCsicpgxqUNSNU4Li1vTrSHxBfJMO2kjzTT
Cg6+Unr/7bbiATHcgOrNFR2Iu93bkPgZI0DNOthC5IJoBbrvI6GkSEZ9e1rKS2ORIRKD5kjmzr6D
CGkwYaHHRrjiIqF9bdrGmoyfXs6cvezzLKScM9Tb6dCXoLbR8MCUx+noszX9VZhoLy5bOa2nsR3x
+7+cdw7wzNiBgP0t2eeyNiVA6BNL5rZzoBd5l6XfC5pfu9RHgqNkIK3qZ5SzzWax2HvuLIOoDtRT
V9mYLQYrfJe3XhDOozb8bkdEfLonhbB65opdEiANGQbdD7/XWMab28u4fIHmpf6U1J2X8AyDBK3l
A4B4QPCbXfB74i5tN75dIFrrxbU7ieh3Gq/ZykBdAu8lJQqQ/Mf09YbJDWdnHHNPvz8UNxCxhVjg
NmJW5PtxsDP/6Nwblxp96OQYGk4sakPD/xfSh9Cw7mbulXIPPa83l2jAXQvMI7Bv8uTxjfAIofzU
uXcdgLj3nQOKOGdRDjBTjW2gf3nZkWtvX6MFVqKXQ0XgcPD1vEpJIX61bcyOD+XTXUIfyhZKqzWl
jiQeoN+QBCPHQ9zg4FzsbQursCcWvuPE43KinsqP5MyTEy38+V7vIaj+4LmjnAzd6k8B2a5RTq/T
Ojvpy+FJOkvvYYVBe0xf9vw9QW6NUKj3ZPq7xzGww7kHdiwP5xrW9Ljm3YDgIcWWYfmlMbW81Url
JyRGza7HwEDn3AOfksKQHuHoLp+pTgS659G3DItMW5bU7bvEdLf4ijRGMz5/7JuG93DaigISkFlD
EJ2euBwPkgvCUQmX+LxFSjhSneyLRnZnGu8y89gkh6C+ZuPBn9hF+rBzKXk7gASx4f33Ybaub7xZ
bQmDKtnzcTsyCnICKvNj15aQghxpEF3IfH0fkds1/ad4H9q3c5x4GsUyO+kUWU5QxBcKUmaswPkW
21+3pzFIN+aTSjEonwQLB2IADAmj64wc6idzZaigawtuw32hw32JC2ScGBiThP45s8fcl3dHIG3D
in8eL9matBxKXtgD45Dg+Sz+RALiVxU9GUbnSlPs4AdS0oASP7W9oiK9BwYbXZNQx2sB50zkm+0G
oyXR4+AotLqksH5Pux6KyMZioF9CuG8DzjK8uovDH9MGtUwN9/Y6Xc/15aVbyfxHChcGx3PrmC4W
U2buNts64HL1PpX9Tv64XFwNs8ydXNRooFsPJ/3KGh8XsvAFWyu0S2okSNWdd/gEqKgs8H9SF9vR
YnuRgzpSXQt93J2OF/6a3ZrOWqtFtkdByAxhnI+2p1Qs7KB1WmThu22nmFahXAYqzO+rNzLkGHI7
vCLdGh70o0rYhWqcR11bszsz2nRFU9uQPzgAPyU5kMRij4AW3nv0OlVYLnF3sYF+hA0GK2WcB83Y
iWCKc+o5jWIMrE/4kPR16ag8URjCUvSey7cnY0W+MGP46MemhwHves5rDfiVClrNucxb63Bn62Jk
ubFQbUBG3ASVQFKw462l/HI4R5sXvPmlk+g4zwYh2o292vPxhO1mlIx2dMWSzfEJRwlagcvsrLfU
A6gcqZif8i6iEQqzogCb9W+OGZmF4bRzRlTctDks2nkw5eDlJzx2kc978ak9GtwDlCiIjz6Toayb
R6l31f5pl3gEzGlqjPxQIS6GZ3ywbbYVXdWlP+oYuP4L8llKoodHq7k9Thff8McjysCVBUaTZUK9
5KVsTv0Ul6wX2qlN0LDpp4NW2TbTGjt/ajFTGININ2AXhrUYQGD4S46sTSDxd7jgSnGm9udCarVN
9DsbFf8zjlmjKC41OF4T4Uo5R/vZ2YP1Zw/23q1ZtNyevMZJESrjpO/3CWWIDypv6q1YxtDmQXNJ
g0oRUXpnTg+7hwzVXb91kPyLIxtN/qJdk+BAzLh2vHKIwnJEghCCKZoLorSaftFyjb23mfhyVcAC
jIyVzCRhrEDTeBCLIx27gGJZP6OKMGWBwihVnonNSEPkPP5QljhU1mA2ICmWsuSIwZ+moOTT6h37
ye820209i/9eOqoEOtzyIu+jczFc7p0bBEBYn5kUwL+1qjvJ8RUsLcJPZnhjx/U/uxPbYwdP1LbL
Njx769QbOwI10xS/isc4M1PIjdxUTXHrmtuNU1LuEC7/OGNyVimqo1CRGKDQ5QLA3zkOxPMx/yn2
VY/lUbJSCJqS+N9stojgQM3aO4aYVhNR9G9cTs2fhBBTkgC9b+53RkvLMpKmF+aijynovlkc+B3r
UxfHkaUrAMvatAr+21ZVCVCsJa894kPjOF9DFoNXAXLBV61KBqK31hx9887RPYHdwNQAi6prCJoq
c568JQDiNloDUF46Cmt2mlveA0MkjwfOOUvhWA1B0Ou+fRWxEBX1YXPcSFRayxZtAsbXjp7e0zSg
+dTlV6Gd/C2VKrLHBbvRxcMpDU2qhZejZRI+NefRgBfQ7IbVBMcrnrjqk68hQVaO+5/Qhs9gLDKK
Y+nlez8mQ1SxB77c/XpanpNG4a8ohEuRAu10Ubn8abK3JEfeBt2XmqP98yWYF33NjfbDYDkezXAO
rWhhpeC4yAWir+kaETINjGIRJTmS+O85W2M0JF94FwT16IuY6/G+WPxsNHlyu1LVAnfF71/6pYt4
j5UPJgSqKHXLdQZxNQ7Ayq+g7o+1Cl3rygne74wMX7FZoYzpDL22KLImxao8y0iElehP0h45kqma
puH0jKPWk3akZ1Aa+qAHtXJaCcp84jBa/vliA+OWS3xSJEL/SM3l70SDixwOTAX+OpOuYq38ISIo
0cTzuRfuF8PR3H1i7UgV6T+eYjNtepHdaYOlSywYJjxuyyOMha0IanhoL65SRn17R35HjkMNa7ZR
jM/FVHH6hmA35mavspHwp80Cdpz3nR7fdcP2jr+FWnHH+SHm2Rqg5z+LBaqEVvRxRqu4dYg8YJcq
msUBmPvqcs6F5Srt5/rcCY59T36qqxozxLzxEdjeehpwR2VTlbM076Y1sy4Vd/TeRZNq1TCBbnxz
YJ32BqmVAxC/8K3nALIAfs92CqUy/uW1YtqM0GoxC9HRnqinmQQnSy6+423KxONfiezFqMAkkG0A
EVG0p/fAmB/gO9ZC79lzZ3I0UlarJhSbNChr9kTfrPjPA0eG3pfJVMBWFykxE8acv6uAXJulRcjt
LC2mFWf0toBZbDobxXuYwF0m/BAuXegyNRSgei6LE3Z84rqBiVbAeCrg80Tw4a1S5nzK9qd3/FPU
ugLutnfpRA+fH0hPa6bhFtpjDCWsNMLG3eGzaCHgsksmVXzPbrKdVFQ+ur7w6p2fB8R1EIQ5Aoew
MitGDiffPSlE6JKh7brI1RaQOaWYXuk+kGazONOrjR+nskvZOEM61qDfEOdHJptxcTF7zSMyziiH
kJv81o49zvSqKsbK3VjWLS7E7/LfcyftV6ix4VL67807OzAofUG26gd9It3zmojB7IcKcfzMocXm
bpZkoAP02ZpR2UUejqVfg/vDrajvoy1N1kg4MpnhqRiPC1FFV9cbK9QNOBRZYDseLsHBH2bvzRWD
8SPkFpWk3CISctwkzSdjykzYyFA2vKkYgLlzm3Bpz09YcS1qlSgBasdY/NZs8EbXvVrAhrk14l0+
3P17/ZeZrCTW1vXGWuCxE/3VNwD5zoJs403NwULVBD2QUFbPUtt30W3y1AnpP1H8wGff7ufyaTq4
Ls/ybbu0G1nnpc0PMIzHbK12A38tKw8jSX5gpIhNw4sd370PbbYXX51kAlQDEvHaB1uoGtnk4BOx
o1PBUjfpCt0cW3kEeaKNdXiMshEx6CoWxgNvpKcKJdXbEt02uDlwgmGbnJXe9st7a3DXjzJwyCKL
nq8vbzOPuey+g3s0VPAuyKz3ei3k2fp31KNXYOwHMT8i8s25PoTk1Y980eSHiulrKj4Vc5j5jLvi
M8IdenlFRjvoXGDwYDd0na0TvgWRsxlgjydxcL7jjy7GnRKPdJ/4HEJvyXm3NF0CQSzJNZD6cV95
dhoWb7iMwBL9nTDwIZ+GKGiqdo228EY8UrVk5rxFoV8rRVYX3ysG/93LIFnQuuemds4T/s/2CxX/
YsOu96UCa9gx15KJlPDrGxlpjxq+pm0lZf/7UZ+WEj+Mz94uqM4Vq40n3SYLRvxVlFVHb6Z3MrAm
gq5ie0muc4GojGDjXamcdlLvudq17T9Dv4A3SSoJVl9WdXWJVecD1V6Uz7N5hQSzH9gxltk8KtUN
qp2Mxr19Ooew5Eq1eKWbCb1JZKTttRsfVyosAdldCcGjOcZfFtToZC5ax5RYX24+Tg2mWTU40ozO
A7WTcgGEBeB0V7MxU8N5zO+bx4cMRp2sdWAkITczOdAX8GtPpkyHdsrNSOcZr34r3+gdyuvFG2l3
Utkg9VclFMPayKAnZWavTlVH8ZCMsoGO248U7ILAOjEFvNnEep0oQTYifYn5DLFDltBBoOvyNmSA
44h/SD2wyjCTjAWellnsniOFNAi4Bis4mLu6XWJfumkFx7vtjOI9RSn5earzTAVaLAs+aTbFVMPV
xna/42PJE3a5/Jl4XrHHJTjIhDNwVu1guda9Hhyxn5TEkM5MAruxlrBdKNU0eETJHbF5K5LkMKTD
2fhumIvPACSl0eD+1DO92Qdi3+5T93frJP6koX6814acONKd5S8zuypKp3ls4QFvJby/FkNzE6pz
FKPGcprzFBZ2OCMfa9vCRFezka25w5UF9hAtu/mvhIVjauGpxMKmyJ4+90JPgO6CPwTrwW2eGRMi
7icJJjdJk0i5g13Iz9msGWSU0IHh+bmO5rWFk8DUCqtsdzmkfU3QpENMfZjRHO05m8bciK+0T4wG
LfAJMdLfug+EovfuzNI8eahumeq+MBRU1NNP+fCh0yVSCmBpMdPJ3Z3C4pflUU9gBb/5pwMWksbj
aPEbU0mbeT7I92jTkxhX/9qqsYQMqSDlLIf7XnSnL8LRYEcyLpAHb/TGmqHQ/ewZa8DGE9gkk5tu
I8M08dpkC/DKRrGsQJGuOLTBKFfbDneC6Hzv0rOb/bZhJabGGxDCTkZXo2FyIuNdD/uNXco8LzJI
HL3dVBiewfg3+bawc6xo3P5F8Tb7EzVWrPk5jCMicAF6dPf39mRq3XpgQdL1gFXOKRLG7plazjmi
Gjr4d2/obIdVBQ5ZO7IjBicRxrkaSMF+oYR3TyUE0NWq9qElJcMuSf3JD6e7tfzQMREcVTrqsfMP
8mQ/vU3A0d36burYGqe/jr1YLpFTZsosDwGyH1/OzUXljHXz/ERdkkP7uOxoHle5Yvspce/lCOWi
22sReG74lVe/C3mV720FqQoRbE0W3wFNxGxFIBkpj4CUbt35M1ikuKZED0y2/1/wLe/1fppYi2oN
6aOIed8Cmo6eM3UteAP0bJZUSCEQydSGrBmftUoCivgOExAnrZW+/apdhnW31kfpYxHyb08msDLe
kKLf6y7OHXI3sB8jF51yXxPWUqkk4gUCRJj2ptRgNAasJlOP6OTTm7WyirZP4y3nKUPANlE3bFMr
7oCAwlAWRBWE90/YSbZcY/LbrXKs9CP18RQ2orOUjbLge9F4rPcdTJG1Lf3AZbMqtpJLXB7xRZJY
lc5DLvRxJsEv3FDOn5lexQAsFRJHS08hHtsSNgn+0Ja0YlDRTt92zSuXhQ7LB8+/Dmafuhv1wusF
VhswA1FGToh0ThQ12g5FKMuNu4NQn+PNCUyzyfh7T6+tlkRQMJi1TrpMpDEv3YmxWO4m7gnu2jOU
0wmS3cipQURRmDojYaX0C6QlvTSprxje+Xj5FHwFSiG8f2LlKrzqDt5sLO4bxagbdSjrC7P0C6vp
WZoMJlLMSwIjPjEZ9AKDNG3D8L8m1tv/3ctvjPAv7TelyAhePKmWf7Er5WiUr4Fgcyk5inoHcHgc
2bkfTPMNm3UvzOyzJphz9OkFYe0kyTv7GntvcbhFkEg54m5PTW6mBNkfmMZ0MGuivUeTIHj+nbrw
F82JlylZrM6Rrx0gju5HZ8Ftjgs65/4rmEYYY6cGfTV0JWw8KyV2gusMG+3O4Dm2dJR3CvlmXmjx
jQhp/Yg5ITUZyGtncIKKJXVG0872FkCXOHdr4v+wtM+EHv14CFtWWh0Ye/ysG4tjBWg/Hsbuz4u0
KI4RoRFfazRyKGAa0foX29ryOf/N6hDzkX+kTm5VIaRBRWvCD+mRJl4a6E+3HO84ysdqVELjphKx
6SckATbAYNPo/ySCJlV5m6xtV9+E3jA0t6s6/2v+05+Ru3SoRkzhsCJ7Z5cMlEtMsmRdaDL8DpBr
IgbjuGUUJ05+wQuUnpu+bivQ1nrosubru1Zx/gln6UUe0ENYQSuW+nxQmPc1U110Q86wnINcgBhs
f3H6MNiTaTG3maTSsfT74N9yh4RTZ5rv33R9PhLASDFG5TZQ5/9RO+VXGtt+XEsRZ/amaNjakAt8
EO3PMChmVR6idB8I8RRKvMFEwlDeeRRMZ5g5Pgn0htyBAXPofCuWHwbzuzs/DwzuYcXd30SMbM3H
vXpac10lUOm9MG1hIQ5j60Hq5yakNbVyO6hECTUQHfRsKIsxSQ1DTt80CDJfYCpG21FhrW9GAYct
FuqVGGRQJPCGSdrxjkccmJDa5gjfSunQJikr6dEOoznlNgcM5xVTWeWtzyKDakh7Bvp93YeRc6bI
0VkA7u3akYYJfyB+YuDQ9gIvtcBZ1svGJ/YN21kYQ6s0GPRKLzuxq5n50Wrk/YeLrZqcuR66gNkG
u3A52a6dmA9JLTRLzUD8Cob6ea7+rQu8zQzwk0QTDbbl8DCcAg0RkL9SSWojo3R28x8+Zce/5O9K
ub09hkLIPJvQDjMFrJnjHnhxjhvVmYSoBBULHg0M23YVmxnt0JL0u98NyAsql4jeGCaFuh6qhp84
mw9wOO8BMQNj/nYJgF+7sgGIqWz7EHOVV33GPqZxlEEE8KfvXPCpspaUiOxok/Jy0gEtU5y2UzP+
SphuWdlo9RArDTwe09RsPauzEfqR2b/ahl4DD+nOTWuFlYujN9UIJb47QyO5C7NHwUEuU0JWqI0O
ReziGw0z/xZobaJJFEZNJkB9y6omsVCbDdvzD0YWdgNLSW2Zybnkm7Uh3Pdk3io7YFZOypLBDZiQ
xyKaktSGXGJVM7xVUYGg+obm93h55V78vgtu9wihSQdvqvre2alqkRu7Ms52OVSPUiKeTV0+TZ4K
P7pyoOG+ejJDhMSjmdNb9w70cYxIJFa+E/ZNd9mWbl+DqaK8Tx8PB86gCgN51qsOYqpHBzy6u6+6
9N1RVNu+L4441oxbobG8axZhWDFdaIU34nKf4yxHmGkh+Nleg35QDKq5sN+pz0BqHfXql/+FXTXd
M05tqjfwwyaC2SoZ54scnTvzqbilexrYMq92hSSARp+WAGLfhvY/dNGMnq/ihAE+9O//upasceh5
N/bBYN1a6c4YdeT0sM8f46iIsIgaJIOD4YRma7kqZuyFy2m0RKq3qw/FOcXycSNEFLs2phRmZr5C
+cOO1z3QRnoua7B9kZLmjL10RuctHYbtqNmEk110v9WoOH3GKuYScK2TmVQoJjl4SawEYLkOYYW/
PLi+pl6okxH9B9Qscd5MYvVcQv8mFZS6AGbQbWc/kJrzuIS+A0Qu0v0nWYxlu4ZVqd0r821cidR8
Mu6YYuNbXvVggY47ZkqWCMf2odkoy4cziOCfMRFtubMxNkzFbsboXUU3jfvwnozWyFnAfZbbFomy
jxvC9yc9NXM7rNd0ZbsHqlK/G2eO7N05wZ76eSPx4F6fpdusARNPxSGIN50kFy4np5g2Yf6fMgAS
IfpwA8HyaTP5tzdNi9XVe2rz/bxspTy0OJyyIV9Q5soU0O+J57ew34hsIEZWN8QdYX66tNX2HXfF
Bhb2DjGSK6wdjc2fncPTU115WuFqRM2Y9TubZ9OkR5it3qX78fhHVos1EI5Uza+Xq6bhVKmvGuaL
DbwDSUgKk8SfBr9asGJjSR78Ekszj0NCzNhXp7juw6JOPAzbo7yBmCDrPCVh2xk3W3V1lC4B0azm
ntpuWpsRu5+t5dlHTCWpC5xlhl7a56xv9ZTeKOxLfYNcrDHEXeHX414+QoISus0DK2Hwh5TV3w+6
LYhhow0E9KcN2c+/S/fZIW9ydRIV7/VzZ7Wx+VM7arJv+iBNMEnm2G2jMJxUnUVB/+ipreXJH7dn
KCd/qepK9iwioDmhQPdKJwgiZbcB9NWexWraVU8LIzzs+xeTz9jKabGnKR7ZjlTTbVBw1ByZa1m1
nzdwR6VooPm9suCzqXzYF6sMhFqFQSkAGrK/RKZ5ZNxDX43Wubf6kcrRnhflpnENFedFVzE7Y8Yx
MGyNmknVdUMFRv532osJrTIP4DtWvWowMpoHxSEffGqYUic1CVE+rxt7JW6brMX1iBUYMjZ4fYiJ
Pcp9zOVSof1GfYCAWQXi91QWczmH45Y3Ng7GsiuCqOr+Ig8xsKT8p41/Z0tKqFILM1hjNHmZL94l
Phiev8Pe20pZ4/Pxi10nK9bYnie+esjF4xTTJcqI60hnYmamGFtdyokdMhDxo7OKfxjswMJosl7G
D+6fhhTJHqxrGr0n9lI9q+mDlG2D/VKta5MMbjic1eeoqO+5OjHd0p0Zx4VLy/4ocoznY4jQ4cmY
OwU3hmqfCtMHzx/tZfXC2FiSgY/o1ZFpABdyCggAsp23/dN1/jYFYvlWbISUF7e2yPUwABWDniU2
7JqJyiMXXvbrDCwv0rNgqWfrKA397NdJWYCnCh8/vfqeen8yC/hZuwYnevP1QlexL7pdre6M9tfY
gIo/TzsdaBcc/O5ElfXkjAVaRAribLJrhb5lEx2qujGhtFWKCs3ZzdnJu7kSfjH8lpF+esrdcYqV
Pn5e8GnoiQWhW5zh+AZ4BWVDj4ZXZr68Ume1x903I3hOUtshPyA8Gpjg7tyMAfDbtj+I+5z02KSD
XlgSOlnVc8j50Do4CsKrHWlnyilIr5Jynej7N8KOOQkMCx2WVnyk71w/9ou8FMrc+f+LdVMTGxIK
8vRSaFD16OS+qUsrb/AOSGXALMcre2+jjVMycEKoDpCMlYcqru4y4E5Vh9IMWDshdEzLF1iUwlRC
rYCliM2WOvMwZuFUydPjgxOw2Lt5VDYM3cx5ZaLXtx8trN+vKMcb3rbeHvVrA/tvImFFNfcnH5gc
NF+EFa46Nnyl3EPYwd72hmg9SEv5P8CPVcaF8ZIGl/n3Ayo864Qem3hLIzVpZaiz5/StAJ8MV30+
cB2RAfEUUZv9pZUnGiCEpsU3qO5ou86xd3Y1yFJMHvIq0RP2q1IyhQDEyryi8mpuZYV0AjhUhPnW
mYuJcbTOVI+2Yjl7S1V3lhdZOno+XuSZEDeElWci0N6jNLyMo5VEMwmXZR9QlFdm/xtcPRHGTusQ
rG4RbOIpRwrijl3TqOobImUslsZFc9xuwea7Fgt6C1AicUvS7SPEuU/OUj5wQ8YdqyZ5eGwS3TwT
r0BHxg3Gv8aT1Tns+xwRcguFRbW9kRQTZVVJz7ymygwcfnT9KmtTwlIBLXM34T0GRyGkiZT77qwp
JYiX91RTLLlVx+r5d+Xcg47zXOwDOozUzb/5Mm/Fgb49LJwELXJJxb202bCQ+/Eqsh/DS+bjj/oC
cj6uAcuMr1YcmBalbcOgA6p4uw/V4Ftew5Np+UyOT+EUiZD9ANZ4RhudJuGqfBesWjnYtklY4Ggd
R+V0TXxBKgJ4l/4DP97Um62sW/6cIHTFcGMxk71iviL2gThyir3m+TK3qj3GkZSuoYVf7MDRdtl1
hbtCDOg/Y6jZfQzs9hHmOBVDE7jJlP+hmX02nXOToVN0Dv8g/6JGil3e0uRJa3Lf5jkG9w4jHGVn
pCka+vleVuQrNGoySZEFHE9PFyJxQVBpkVO2YuQUCSvU6FHo5HKrMQNkyg6ki1aZ+4QYTRN4oja5
r6qvzI8eLxBgcd9F1fsWK+tGE3Gt+6OYtjtF10Ody6fyIRdLmTRam7SHh+F8CWUQKQ3NyYMhTlca
Yw/YPq1jwOvn7QGFS2024viT6//q3cVl8Sd2ZdODtfifpYQkuVnjcTTHYCd+raF2mo1pYZKrPDEh
lKqUUeXKB4RDOpyNFpYwobYuuE4Kh7JN7znrCjaS8br9xDHuTuJ1eeLRNTOl8ifk5dxG9Ylqhzf5
sO7mpqYyfGqvUEiNy+rY+7OZsI6UjP0wygFl4i5JG1f9nXS6KFzlh7kqEsNHjR0GqeWd/6M3424D
iOXj5S/E43KFRIQ5n+LsHmGe9wlaB0WDetNVW2/cGxfLc5PXcg3UXM30OgTVsLVFXrbmBWihbyeI
lGJ43zYWZsJgNbLfusX+jkr+x83z7uwgUMGqeQtJwSTlMbaJlHx2mtHQ1qOVEI6Gyt1rIYRkab84
GtYp5FsaIjxulMwQl1tVT+6UXQMuo/h9uLJiPPrUr06zTc3PjtxOtDUIe3P+zTHigXDoIBN/Qz1D
jouflCCHAe3XacJsh7O11nQQT0bCmjsBm/6kad26VAUbmzjyEE83moUQo2Z/C0XyxBjn9U9fu9ut
5EmD88MRx1FvHxmxIOw+mrXtSe/UbM9YLybVKoteB7AYiVON0GUZdvjcABwYweMY57DHPv8O7fNk
wr4EMUcKwD7nZWN9ZuvLnGdKORpda1j6eY/ZLS0CdAHK0Li+F2vz38GHSlVatpnEsYa5m64XvpDF
qUzK8kju2W4S1XKhuyUszoXAQT4Kn8d7oaDAJLXMYFpMP20KMv0wmRFdJdrUnY5ttVn6Sa8qYCeb
DajY8BiXN9qP/E3maY5h0c5e1G9o92STK90Ce7JZfWo47SesizIQpCQli6VyLJeiYvIZrlL/Q6Oy
gXhwyDrm8NJmgQBM2/+yRsqi2M+f52iFrR9c2OFSSuMPnJoDJ21ALYJHMZAvixKdmry8+VMy+E18
qJIZeLafoDDFQX6qcWUT6pdeMLfFvp2tK01D4SCrc0UHBLOEnM4oHCWSMWnPI3JoE0oBGgi5Xonn
VoG+tbv8/zJYVxHUTYvgJRGt0V+1+PXr4uFJMFOz6J5Qe3sZV86XxM2oFmgXC3GVwSP68HrG5Ws2
Vl04dfhEmw/5WvkdqYhLR9nFkmWUvx9yhVDX8Sav+idpJdzmTI/Co8mcObcS/IYN3rq9VKiT9hhb
tsasZw8aVaMCrhVRzMJEPOzcrknOvqtJPCOFNw1fO2pRCdIUGdu1KhkE7TaigXRLpwMzCfRe/4kh
MFUjn+d26EHnPOpt/oAJHP1drrLm0LHnU2Ai7EUWpSfiboTvQ9/9CSCsJScxLGE7Km1zeUkMjFvs
BfXI/JKSzzV2/RjfReEf7keIW4CzPO4DM9NLnFaXwV7cMxst6AI45X6fkgSNml3DKOimzM7GI7Zi
gaCCiPw258W4YPNfSh+3BjHIRxHHnboda2s4AjgvoaZRryCmfMLZafHrgnlDBQY7hdfytztL5Og/
GiLgVx4pBFy33C48MikZnceyzFSjZXXlqj80mdjdEoBSvlCr7L/rn2/JA8qMSP2Q9UurVKdwPvLo
W5fD6LQTjsPlq4+8vWeKKGpO0+rteIfwVya1K72daVX4SxiKWTPmUsulHzoKiqHRZSD9iT5SEH1u
ZOT8HWWqB40f1B7vYnA3lEzlVNpzCzA1ZOUKXEZdQ9vwOBAlThJsrioiaY/fyHOKj781U0wKVZmZ
bzIapqAMJXxF7YJ+Mw+z1a5OxmFNnBSAW6sgjm9Bgp+e3Kzq7bnh82JCFFuOiM/E3IVhyFM5Pes6
K8i/y00MV84YYj9cy6HanuohJyGmIeF8b2hnB8GRwkn6wrI3yNBJyNNG4m/E8yMTCwvrm1LxSPSl
c+stf+WpbNS+FhnyuSw3WlOoJfahXvuHsm0e2Yyjycm2TOwYvneLBBvrB2P76BKoHomqiYGk+d02
4fle9kOJrX3iMb+WJtujRUatjK5mjeTcmdQIZ8FZWYsIZD5kJxPB3Z4mVGzJmOG1HrQ4/6F16t9l
UEt8+ErvyHNzYqqbKGixPZ413HTX6+qbBS1MHQwZzeWTGY8C8hHyVOxPyycZtnavX4JZUNlwlIsh
AQrb69BNbzw3pk5JC5fogpAtzYfI28miRMCR/0FJPml6B7qSSsLn+Kt7S8kyg7cGhJiJlzwyLNdY
EcgDMcA7/orl+8syCd2xv1Vnf8QbrTat5UBGc02KMq+O5i3/9mk5S51g86dx9jAdpyDdlnHOAwwN
ha+CF6o0TuLwe2BBWBQXH14hVd3NwqOkcvySlRe1R1bafhrDOt6+B9L+0LqqhRwe4ytx9L3puUKv
OH4pBgsKbYmg9htn65ObhyxR+b4+K53YBWCN82o+eKwZi7pPSi+rWdq50OPiUDq9CckfcPOFpZw/
GnIj9d4YvEALOENujMncXTMNuYwmjhdSba0qKhVbDeYY2Q098su2n9Ertxqf43YIHxuUQlgiOg2e
4z9fjnO0T2cBGV403pFUXCxu7tKCM35+KFC97cHtGYJqhkXl6vkPvCAIRIw/0HcovaOIMnANOJDK
UYMcWjXJlM+iE3jjyr3v4DZrlHA5cy/oV93kXxBUSaM4MHqPqdx1UyQdzrH6KbmUskZIJWyIE7wU
PLu5/xF3w7qosTjXMxqsWLHmnD3mzyTfIW2qnEIPeAArR8cUU//H7ujRx7z8ch0hS4a3YG0G9tOP
PJ3vk4ZT329pdMNtipCikQOMMf1z3oURswMPLWwpxh5NrIqrHTTenTj66pcO6hIJGgtp1X+YeJNu
pDTVhLciNfoIanEeCaNy0CUcnqeWO2IpY2A3XUg2U1nJBYvRhi/b/RulAhahZhoaxUD8BWcsSt+r
fpBl7HCEquR1JdDyn11RJPILSn+OwZlhqrQlzkkbmjz6F8K6AWq8wNpsFgt8cp3WLcQy1/56APII
epgekWdgJwEB750XxyLtTTOqqLLjJe5JH/GmUtEAYPpSny/trDwErYCxICoEasFKICJ4lyIb9U7G
1WkfpKB6wDVD67q2qfyx394XuwkR1mpSvFX6P7Qy8IJdqgqvYnDEnriPTkhsXKqKptozmWGbeZHi
uSG3IoIZoNA2pW+q4CZ6nWpNF+rBQ275LR5Z1P0Eo7oM0+yO1ABnzm1aiFTDHk6ZuOmLhWE3vnyP
iIFo0XlzeV+j5MVsmtbA9YSnTbwqZ4vWAtNuiIcH3W27G1VGQdg0Dw0oPmQjgaElkUSbBeaiBVrW
3CvsXen9P+zNmELI7Ut5AmJ1raoWQt8N8ArLi/YWufBOfKAsOVHyDRf9FzLn54oQoYE5hP9Pj0Lw
x9FBdtvYdNdmjKigIMftFFEE0UL0z7jkHOtjNSJC6nHcZ0Y7YsNVae2kRxKNPk//+3M4sRVnMH+n
5MesuoPUV+UkqssMX3vHrriGiD2s+MN5cjWINT8vi/+0N3WXmXM/V6JTbkOmw8laj2WGFgz0SbB1
0f9Fac0MY60cS7nNMN2NzQsCkNpFNQkoc4lny05/shc7sZ5PO6dTppk8RmixgNZcxOPf7wNs2lt5
WkSIYZcmWYWHB4f4oM8P63wAptlsLnZKTBwS5ReMBKU3edLsGwBzHN+gLb7EKeJtWjrYTNXRcBKl
0PWqV2hkuPN36WRceDTFu8bOCqpQipsIXhPzWcK2+oIpumVoT7pGt32M1KnUDXzFxJBIV30UH4Hr
0QqUxV1iw5KsoWn/FhvEUIpSycJq/1RNiXI4TJX61O/i+HuHtSZzveETgiV3kzYsT8jDZO0tZ7Ok
1hKF67dwtLo9IqJZcjBxEuR9WA3oGlf0f6YKBSAG80QjiYydhqq/qWbT6gbdS/Bnji6cHnxKP4da
s65Xn7nQg6cOrd9fsgrq2Q830T0C/AoS8cfhKCkFcnmNkw1AHKknSA5kM1xFf4xZP5oJGHK5wl/b
jzFXlu2brVu6eWj5NrlosqNfXpGGjZUCLtC7JZNkUvg7xgOZxsT/y9Ns7c5tg/dQBVIGnEVADgHd
+Kad6wPGFe91f0bNIuiY4XUWmLl8MN2xW9qlSMKc5plcduzyyuFznuvvAW56S4nxA3E5Um3sib6F
Ja23igsUbcwTe7P47Qtw8lPhXzfzYPAZ4FR0knwBUnGM5xZJkvMEcSKH88fa71CqCvrsk74GxoHp
dCd49IE2U3aff81oH2ZMDEU2oQkQFKpFh92EnBvqrApnBBuRlrUolYrH1KdXaWtjj+7/aInKfhNW
5Ce+FR2IeFsvQN7jjGBn5LXdSNAnaS2HUuhs6CbOX802TXLE5LpkFei87S0+bsYAKMra6QUX2stT
Poj3c451YStCG+MmNTY7zM8gukzqxC+aIvLUnrX1MLEypx422cXez0xpeZcyfx9Awy7e/nxI+f5A
iqDNdNj3MhIHSHSMFHCPCfKDbiZFJVnnr6noHza3ywFWaRRu1Mup7HA3swD3HtBVQY0dSMBARvj8
kj8kyFiLkrQHZZTPZRW6xEvIRDG1pfrspy+9MsxyrW2N+KyrFwfpngIZ04V/U2R7HmDH3w7vKtFu
QepwR26eFpGrDwMJRnvtHXXXaaKhtmZN1Xql5QOorJgnSLx1foXfI8mNTGcVAh6YmuuyeKVr9vag
Nw1m2YXt0WB1Fx4PVnOHu4utNiR8id5JskHY7BnFXANc8AKR03QUg9BD6oSgpVhtD42cZ0Z2xFFN
u+4h62CHC9bOX69LodNp4scSrYikm4ZpWxxu6lgERpZB//gbQ3vtB0mRuAz0b8tX1h3ZJkzb5yzh
+SXo5p0Crxietm2bdDhZU2fVmHzPBkkQGI52g5wHcYRh5q5FmB60L4i/jgEaFwmDSZwllRWHPYeW
8ygLMulG2kwwncbSdTrDZobdplamZ7PWKy6/Za5gi2ChPLFHpsEcpSXhy5m11voYr0LRRW4R0wcK
dsYbTILyjWx5MXXIkiNABFrqnHsOLf7AAKEmVtEQRsJa9J6qEzhBG2rCSzBD36PldxwgkhGtF4+3
u75jrAYBgYsSpTmZm5XftmxYK0iz0JU+31qOL5G3UrOfVgVAofRchF1zM1z9yN0eyVEMAT2+Mbtq
zg16oSnCevt6eVYSbVCGMpcnP45qKyYP0JxXTuB16rRvW4rO8cRSjsSbDsFzmei0eFuMsqauS/pI
0TUPD6h701CEMj5sxoJkAqaubQ9zSeEl4wM+RyKX5U0HeCZhpB8vM3Vo6euYxdXyL2XftyhFIwe2
lOxCjLczfC3RHqZ7fj1/f+nWte6WToX918HoBFl6Czv2J8HYR7RMOGVlFhWZEapKeDPjlHb/B4VX
arcLoP1GE7bnsUlGBVK6gL4iIAVKZ01BoF0YscnHz83oBmgKmDGgLMtJkbYPrsMx7NeKy83/g0zY
RrLYfsJkLKjILd3QoMP+W1Z4TXYQmtDFdtxSVvrxAOx+IByXYk+LtOyKZEwlxgZQX7LQRN20WSx7
QeAFUNPhLErLM8nrm3oaGBvB2vAe/3OOpYxinbu+1K6zAMJKMOXqka/DnFHg/WICnVjkodpnKltT
IW/s72QWpTDwmZdqYtha1K0/oHDSx7u83F790vNur13DI8m2DwHmLdKfUndJBdl7jl8YVAVQNVCu
Lkt75fNpq4ULiRvyUJFyZuNeeN+7pIi/F0APqeCoy/gzF5j9+3C83opy+2XfJRSwrDVgr2OPHcPA
I1b/RYtZbjQ0ONEDvvzpS/G7U4I/NfXBjmsHmChfRHAYZnUr2gj7luKLIYogyG0RMbPXSnEAKgHO
EBRCNranPkpyH6lUii5MvdSo+YKTr2ctVBRVDL75mO+xQftSU4yky9cSUVyZItVKweFOrLMezryz
B2I6oaAQeuCsv20xYbFCEEEvuzSrLIv2D8LMekEV++xJjkbuawWOv5dcBX2V9QMKUIz4LimMI5/G
Vb/fPfmwG7szOe+x8PC5l9AoiUUD+OvCaEgo2N8CcG+tTEp9uHy9ZQh+TLF8ApXQFsDL+1JB9uVS
PD14mG8vRJyc5KIkoX7snoA7mOxp1ZKTmyAcjYK/JTcTuSdKNtbTvSYeeoQkk/N/gQcriL2AI+jT
F8FOK30uOlz3MW9lauGaQ8cV8Fbn/aLgz0ytgBI4D2T5sy/mmlw7f1pGj4P3doiI/SVRB5riVjss
1PhwzCtMdkN54h5I6NgSfBTk9oMnSlsz3nFC+hUUkqfFTXn6i9xQlK7qhtKUSEpaXhw0/+4ZOhmN
jNGLnbubB9K8Odn809IyuoI4ctleuDpCR32HGNsHSKIyXTsr1IhTvi+kbpoOScX+rLYS1+HnbTzU
AFoNVw3MeETUB2IQf6rkc149iPqSOf2/g2zU4ooUSnle2EY4dzAsX9JAIvJjWX4kUk2lqOKevnVz
1f2iIFPjsHBrGWpHvOAkJPa+KjeMIF0IgtKyJi2AUhQ462pA1IAwARk/4LNOSxHCFscyKDX536LZ
dvfBoU5BM87NBilzBBU1CeCntTf7o3D4gDmqVhPytsLiQ1vsXqp2FntW82ve2qjpcT5IbVIxbCxn
2L9sxQn5QpJs6ZmedA9WdfDnDpwbz6MjbLlSVM9BCyJiI+Lr4cUiFjnJr5hXZt/jIjyLaPalJuLf
zyrs1owUJac+38kOfXfzxREN/w3AUJKXLHJ6ifNOXBbNxFCYTeswCG29/vJFq+6prvqN6YtvwcQ9
Ynt2AYejVMqVqwWctAx0aVN7Eqf139R7DtTUMpsgbWJU1bhHmlBeXXAzP9yX6D7bSf4SLmOCS8NF
DpBNbuSQE4bKoHg0PrMEEi65HqkMCx0ADzEc9NDzztPxHCfBZHsdqL/N49GxpEvI0j9HpXDx1x8G
hibrOTTGFVytOVLr+GtzYvCJynPbmRJFJ50evBgunw7+hbZhbM+dY9qmg6zogCWc82WS/BvBo3Hq
DdOCiQlX/T/YPOnXfpVs/Ep5GFS8hnCfRHOyIaR0bqML5YcFKFNDz9fVK/GsnndhWnYWKT9s90A2
Cj3iCE4eiZ2Dafi6yRkUV5Mo3wrX1NCCYrd8IFEQ3lTItWQE4DC2RzFJAtpBwLxNnqEWyEm1+GwK
Ehz4pCM6QL2VCzKX/CiK+bG8tBZ8oPn3oO/qyXoRTkHmU7MpDOFWF8xDCvRv0OdUv9gzbnevNi5j
dLhRHhw++dyYEJQW93nO3XGq897oklOuBFwS2+QEkM8mpTH19hUoOB1qOuaT6W6m4GSywUDNr3y5
jNyAV+LpJWgE5bp0VEO84fdT9qQLty6ndbuyFpIT41MRADqbx6lQ7Gkvc/gaMtyYoDY7WBkpD4XC
0JU+my/zOulh3CwMZCiSoiBe7F6aJceNFLLECcc/eYpd3sygSPL23qHK7ZJpdbMAxZAnbAYOEJid
sROo2WMIE3nOk81EgeAUbC6TPH3SFpFn7dchrNqO7LX7Xsi63c+95mtOz0Fr4xRienASJsOmG0LW
7DS2TbOfR8QMAuEg52etX0oMtf8VEUTh/o0pO+uh7jk2jUstyh7vu6oQsdRGOuBOVlreJrjb7aik
f0prkjHGdMvP+o2YOePiVVejSmJjLKAEvDI2x86yvwWoYuWZz4UjGbfIqLb5qufum98WL9/6vQl2
NgNoC45v/DvEQ12uwP2/bRPRkk2hdCbHHHEmmH5iyCFSvQ9ql1OF1hx8KH8eJlvtgnmzUIO8Xe2m
q7notsfWFZITXMyyZdCBN7yANuX+uZdGpzvmUt9iL6kBe3wuYqV78Ct0GwGzO6XfqkpMKB+1xlgh
AHyaGguDhZuSPbeHVVsgEsvv7H68WibgHEZbzKGYRb0Z6uZNDrBKrOn4XZ65QFoLOv65nM8ellFH
kEgbznTbXwUoUNbzUH/5/6VYyOI2H3II3EZAAFcl0grTVP4C5NqMVkLrZ4HZ3q/+FRgn1i+l8VJ7
opwzXCStysYECnCsYSJj5Qz8i6VuBEmzW0RN7bgAgCFhbzuzU+jkmjpGF9PL83EbeVOGKbIScIYl
eRjuHAkkouRuQ4NloUjSMbTpjpTNCQNNXRe63JJI3xjSLTiE6i0yEvc4jyySkhyspJTvlA+e0xna
4yytSlxBRTz5a6ydhBfYjd/nuJPiDICl7d0/W+XjqnWsbGMjhv8C998hLMGApviXsGqT46kys8+m
yKYDHnCgiXIlJDJyF/4WjYS41TnAATvZSPdhEK46mSAKAWjDYT9fdoqi14tEG5cCPa/q/s5F5Acs
nwCC/sgsKcSEehTEOo7iHlfgM2uIeVtek2beb5InS7KugIYWhJbgfvZjfXjpdWQpWrbphgT+PiMC
ijKvkoYV8OUVDOtPTQCaO7pUfGW5UCLA78Q43Zdip7i1+PCjeE7aLquKQriL3d0WtyyWvr3Z9Fl6
8psCu/n3b+2xR5UWqolpbrJlpVOVHJ7jVY/u8F5/fxf7O4CIBx+lUeOx7gY0Mk5j3CDs6e3Bx0bE
xbq+3B0122KDN8I8ckfb/j7cJ88fV0cjcbZr4iUXP/J7nxI2KL9B7FQbhEclk2LMer3JGJiBPq8A
knAr4lJ4M3ZWitpUBW6QM3JzyyGT9GsqNPfmhqBB/MAK05GeqdDWUfp2W541RbKZYgmW708jV9M7
0Wr+flKLwBeW91iBF1nvhZwP0eEBQSCKiCqcHlxR6TC6gEllPr9mu/Ys6vrZub8ubY4ElkNCVhvl
0GbKQ+/ax3Q3qWajHsM2XVcI6I640yyFgiKaEDZHiV56hFjziOfOcAbkKNS7T1BjBDvYYoTLiKVY
kMXOL4jSsgLYGyOwMpuDgskE8DU2DQw6afR36tX/YXKTr0gPv5DqF3Jmnhzxy/wgz+CSbPb4ZY/X
KMSDyLEIHZnPp5Facm6ZS77L8yRotBvOBnxfPs/3j0pHdtZN5Qjy0DcLIbwflkqF9jJps41m4HNp
Wl/g11LLOYy4DJQ9CT+f3+h6Csj4psH4icQFfwsf7QAyCa7lPEQ+8BZWWgu84TPzw836ivQXsxca
K8XdZMLTS+pI9xnEKwxMfC/Tl9jEP4DhOD8h9Bu06Ruef88QrwNh22CjpqmdXzF/gCiBbc9cxtEd
Itp0Fp/s1E29ra2PUS1jjMnbzqNFWsV1ImLEntYLATKs34FRpmCGgfDHSo4rw7hlCA3ZUP/XFVNb
EEG0j+WGJRT+1Uwj56bQ7W6mikeYvjj9HPeuL495WxChfggYSuwMPmE/sUx+QtHS5XHcZI38XFXn
CmbHspSLZlRfe8Q1nhbbhBfLP8HreaC6BUpnwXQYgE0zSnJJ/WxPou6nAboj67r5jKySTR6RBAEA
YnDpSrURpzGGsRM9fMFtIavD9sUBFSNpUhliGuwsDcwVEp5PKKfMiCK+P3S9nsOGwcBhZAXb8jse
eu+j0TtabmRXnwQiqGxZ5jdO7TLqZHZw7UEqd/LbmU0AjATbzvPmZ3mAueAq1tTfjJpJhSD7URv8
PK5qlFQWTul0CN5Ly462eIymRywTXPaSiLF9LT5AvQwDxz3LYMbO72+GludNK+pv96XofGzgrzX7
kdJvgEuF6+KIeKr1xjYp94Z6KyliCNHQU/oV6bveQH6aUK7T82yicytkJXNx47Tyda9DJadSX2Lx
bdvlZxaOd6qlsr3E73tZ6HIpwXajBYamoAMGXNxxR94Jve/IVkfdXZ5zpfSNibmnQzH7c/QtorkU
AEJcmUWqX6e8/1/tRZuD0xr8Ar+PNoGyD2IZlS/xVXVgT/KmfxcvxINXMtMzYckRLc+qPRnOoRAb
TZg+mI7sK3QYqjuEu3MmjpFFo186XbJgSLnZonQon/tz/zNrwjCEeARAJUEaO6635EB283QOp+N7
PJX/tMayhxBx4kTw1m7wiI4IyWlDOTNzIGgUUvil/by9tEm1jz+Pku3SUwD86ZnO8CIPSDj2MuDn
Fz2P1n8oMpCt8zl1tqchLspmRt7/QNtjmWIcaMIZgSdtPi83N0Zb6qt/+rx7FbGwc2e9+VSVTWzJ
0a7PCV0K6q90cjCcj7HD+xVwMDldBx0wfWHUsshCPG5H06yuUUdNgf17nctQpiCU36Fgap54AboP
JG3gA9llmEiu4nPzNZoDuv/wQtysmUYg5uf768U5Ehc+jJDqlaSeBlBRrPQr6sN+fNs1EZKBriNB
+2xaSFRng3W0IFVH5qyJujQx3BRUQhFgJlk1oPbaz3rlMT4M1AkBxrGiVZXr3m4NqKID7q4ypypt
r3IbexcaMpR96y5r3gJuSPNgTsYBjyOXtP5P5nYFL3gXuPvgR+4cOUeE/lvnD0nUJ/CJnIzUTAMW
Xw6JIt3Z5/f1B2qt7m60vRzAuFNYi/WdOuLKq7dWVMrJfgQJjT8Ez7UzmbMs+yiZiZKHPw60c7HU
XwmKtP75ohPFLJCem+Tyc0DA0+0P3vlmiOxI6v8WXDTsWQ9I0EhlBfMSvoqGQ9Z5Sx1zxzM08vsr
wWNdLrtB/Xcy3jxBFnm7iq24D1bFfHUmfGuP/KhuRkWMrV0RrwMOmLtZSIkgrWL7Xp7VegHaQIG+
kZOi6FHHK3B7lQC4G3+NiQUmyUYpl+1r14+rEdoDB/n0JtHOu4QTcW/JEEAG8elU5RyGSWXlIU2I
NQzKmHQTgfuxJEmyWC1OY9F55Iw9vsMqXlk/l6OB2Ty9RL1Qsx/xZ4REN9jzngoTrp1zcDK82tma
aQ0LqLKrD84jM1htASypv2fpnAvjbAbCMarcf6lJLUJQgor6tjsvkWw9i6GGQXUwc+HNKaK11xcR
F6BpYWQJOPS2g62HjcgUe9kg7Ez3Rtt2tvhBptFRhODlePNv7o12uXJwyEDXf2lIAVWNqg3Eng/L
daZnoidqTPZnYZDLG5CELlZn8uJlxBes2X0ZCLJ+opvOZqXOlIBb6G9qfCacSsShODIul5cm/0y9
7f6iNMlSzIq/5wMgEjIWD5QaU2LnujeE38qy7J/BadWj9hsvaQRsr6/hWYSxrH898qDu73RYo/mF
gvn7FKXxZj05Ma9S7TFlAEGgzKVfsLxKzbJZCKA3C0BU53ec2WWNCnvkrDBwuC36aEpefHszPvvh
H++P2WZcHJQaZTMGE9zmpgMutHuLER385AOFF4K2SxYiusPiZ5SAiuA4L7yrjkVKW7vijulbD9rY
03tS9mG69c86a0Ozod3FnFU8VG5Uyt9zAnlar7I3gru/IJ8ig9fVNIQsjDd4FCzpCenn17GyXo9K
fFKBkHQtAJHHFaQJG+kRpEMOJun98iao2VlluSXQHpepOtGIUHMOuVd82NqqYof7KC/T0pt0qN65
VgFOUo80sYJ7p6EV0W6fiazCcJZrVh8Hua3D5JPjxHTdncFLE0U+T4FWDlzTfhn9VgH3VOxURzAi
gHVyymVVx5qKgcBV0p+MphFeiEq4+TbZm4hN5k2t2UBeCGTf32xvYBAo/OYUwz2LV7f1JZk3UyZM
qdVEr+CFJiozjFDUmj9zXHMQYX2e9JcJPh+jaL+VXsZfUYTjqWj+HNkQVQEt/5UNSFFxf6st6h8M
HEzzf6PEIyUZk7FjcH6Jr7XjSqTb2UWc6aJCRlvC/oYsTuO19aAiJ4cS5Yj6rakFKIfdIUtlkPKD
FBbTuXMWOYjFH2lGDvOA8O6Xy3DQZxerlbtLchVJozDt8rM+Ja9LSe1Ywcn2DrFobX7j50ycMLwF
D0lSf0fzRARGTEiGbnbw4dNdcocU6wQsYDAy8dgn79lGykHBE0Fs1bj9aWQi5d3AaXBYa6XCuqvO
mUUnJoHEN3SDNUUfguOXNYITo9Djh1HjwLbhDnw/a/P+3L/Qd6c5Spr6nyfqHmLDURdsw/kb4eC1
bbxDG17EcmfJmT3JWTSxA3hDdkTU9c+kM+OAp2M7E1QuO6CvU/kLFNI8IinMc3zE++ujiiu413F/
rts96k6wn1+kVXbg2bpiD5eo1DJlvCrJRAaQrSs9V5VAB74j3MpQvWI4ajGBpHClBlPryu0sw8QT
jy+oBHfIX3KTmGlB82z8XG440XfIFaGgSLrkRVtqZLbfj8mrmfRVQxu/Dbjdml7cUxRkYr8UkXpX
qsI3jUXW2niQteSteK682elh/CpwIreX4u8qnzipT6BwyadthOCrPCsqlsWEOEsjJ/LERnfXYmmg
hJpQyROVC7B/M5Kc8pBl+b1z9NSVFL7rsWcRJO2fI8KFd9N7snbsmas0J/nlksg1/MX0zNsOiHcy
mi0W+FTME2NKYbif8pNpN8z1paCtzYrCTKTL9eBcQa6/wZo6ots4o9BhiRJ9q5Mho/BDdaf/qwl/
ACILGreY869jB3OWoUtMp3PivJuNFWJMafAfheBGV2idQ4SzzKf8tuP4PF6xO5YlRvvLv94Ru3Uo
mJVbUbxFlBts3zzK1sI4vl1DBbQhr3oOx4sNjEmxKk6AmJ6ezVtaCAYkvPTCB3GAChiFB8Pxq36u
NscOUshCGMG5OJ0QmWtD219Phbe89Ub0nr1Lk84ct9y43u2sTYN179nEtqo+c4lJrOvVpGjXZkND
xQdHY9LvL8jGrUwb2o0fhx1Z+i8FBFy7YySTe9vjRdN6azDf4xYxPE++gYMwaB9MMqhjdMUNfJrE
VnoGIS8j52/2WlaMfoYeCpKsZSpFE1tfF8/Ku58bnnwXVdvTAOtoAwRQCTjP8hgbPyjvRuzGdACO
oVsJALgX86AiNOHwZ/PtVZh5Z8EkNZ7PhaMHldNtO0Qq99oc6l5IUzweSyEmdU5IbHZxoWQa1C5p
B1AVyCOTkSdvQBhUz/4j8mofi6VD8PD5OGBg4j//dFJanKcPqyhvwLl0OtAuXepCAso4wu4BReHs
Bvw3HD+zh02NV8Zp/S+A+O1azDXzXjF3mhj8so56jGLQCctQ26aULDEP8VIx+bJQSKk/tiHRFDE7
cRn2xrudNq/BqE7TNGR7ZtKU56ZV5HgizvoKetn1/jEKQbaG43fiDdNvTJ/mvALBrTLjnmRXp+m4
SsXN0h1oPIcXdCWTKsDZPQBC75bMTptQyw0MCpvkfVXsutKeJehlRTjLX3Ma66VBTUcQsaOQdMfP
CfqaV88Az7OX275wQRspnzWmF0cNImxNpgvI2sHZtmTP8HGkCX+9mFlN6cHZZT0/p58S86Fcyc57
iAtHhSXB2vRfHTqcg4ddViRYs6NqE+Nr0ntUSbXNGxvS4llDQUt93C57Xm8R4ZWykSWNmFCuNiCs
tQzpYLSvbKdIGo2PKbSNu5KJ4RDkPtxnldeFpld9TNKrnCZ4M6gX7QHonnxwN5g8fB7ALIqobi7R
ZxQpi5wQnEl5QXCNX1/rW3jJK0qeMq4LO7d0eEoOVKatNMQDKb4fQNjyAif541U55a9aslDZV1JI
WV0qIwAYYlIeNK2NZbu2k+JWh3sy0f1bgCy+Azfw3MIiK7225Ak5gCDz4L15WHPONM1G+vV8m78/
WI4PMb+XQPVEqeq5aJxxAFNdU9CeWhj7bUaXT4+pYIy0+4iCU0ZkYYpBjckwDPTqPYvTiojuvlIT
Pr0iMVhOX/YagdTJ1eNsfuYyXvHoCdKl0OENzqHutUvtDfjGjIOpXa751RmAre4fGnbKtxZX/BXA
FgCbZ6aAZyV+jGwfvlCsnvNLbXYf9kO33lK69xvT1XBw7gHUPnTNrR4xV6lytAeWMCRsYDYVHdyU
jZSNY1xHSiw0N5Kzf3NJD0nDaABbZMVCRhMeowUlsZwmTIGHkRVtLBx/eHotD+8bPuURcUMtULEM
7iRNGPoMs5AF07VGdaY87YCQZOxKmbD7r17WaTcLxJ0mTvFDmpTxslAdTrMZeb6FtagMln18/v0Y
t/E2y38PsFnNBMATcT0vGmR0sY/mEfrRLsXHUMfLCXA1GbupVE+lVJpvHRaDvRCVHRTcOUv0PyUn
s20poB2BeR2LjIYr9dBg6S0HpMoQKoL3D98A30S7/7dqiL5yzz98lBH4TZsZkk6clUaC/fOnYqR/
gUKlnA1Q6N6FOF5T8XP3RXA3xCYX4C4z/zUPiTlElLeEsc2oUn9ZdO3UGoCjEV325OdvJ6OQT/bY
Df4ZYTgLSnZ4Ayjnih5QllkHKxT7WT4Y5Lw/iyXqJV2fNGpGoKMTvOPUwyjPCbFLR2QTC4fU5+IO
KN47d7ykJx4GWNs2K2nJw6FrbDG1I3Hmbokf7O/P5J0dcQjZVAjqJNWcWxOin6Ky1H+6CL5cvpTb
jWngVzxepGUCn6YpptYxW7A2hch15Oabu+/mDg/SG8SJWolNPElv26nspj1CYEu6A4k+RaTAgZpC
7rDX0Zt9V4AyrsmFQ6mqKc3WRhFK+Gor0Fx9Qbvm1xEd0C8hcRpN6LRMBDyhbL9Tix88vwBvN0R+
MgKwVxB1M3pLylcjQC2/2WCWyhoWVtE8+FbbVbLDACgn4Bik6AVJ4GvC79yiE+eTwu+/+cliC85Z
L8BKSnybTCet02vNCw8GP+F3LJa2eZ8FdetlAEkgKK7JgLmSn9XmE2u8IEMv0GzPrCqp1TYgVUsI
cAZexwP6VPPlq9z4rN7LKPQZ1z0jC5u1YNgSE7nr9WJ7G5Bz9VBz5Hp807TOLzS8Ac//R4+ELyjG
0PleuU2ycS+Uecm5h3hjWnJNzYeBm5tRWv8CXZC6G+NKnRYD/VD6FTm8/RIRvsmodytS97ybFdqF
+0sszN+Q8XM9JtBlENk5vimghXnpuI1J+WwvzcoZV5K9tocXZneab3zxuuPtu7HO9gYnCQPsCyRv
aUxZJLMm4uAMYqDWmB3tm5qgnQ6OYs/AvigmGsS6hPHtX+BTjjN4hCM6Fpb5bWDlr331bKJ9UuSU
/hKSlgBwYHKpsTBF9VGvGMm23+dfyK/0SmKzAOmFDzVFjy9TsoWvGFiyPOV0aiHbHzjum/dfk9uE
BD4J16HpWsvqd10Y4yfd0LklP+H+dgz3GuOFDk0+Z2NJKXxMrkc1o3ER4RuiELarX/B0bIOCW3B9
UI9mSGhOoafrNhZ5ew52kIUHx21k64nGWsyAfAOE2w2ur9Qm/GUOpgFW6y1/zlkJhknoIUpDPAwe
bB3w12HSEQYv3oWUO8mmZ6C/kiJDsFgsTAuFqFz1ivlm1bauOIYdZX3Gp6sgslxqKyn1jjtswn0J
xcSP/jL0mmX7c2AZ3344gx0wmQJyNwZ4yYt0eVeOWRLlgVB3m0/fDMceDGSfu7Z6exuknlJgms+L
F15W6JVOuSPYOhTTcBmu6yfI00aR8yweiKHp7w6wjVN/3sMsNCv0vNzrSxCeXh/5pGS11fErkgow
nLNu0MhDFe7vGDtF8+zLJZcIK3/gyn7R+H4xA4OUKrbJi8EpLPJXvbr1q0GVy2bBA6jmOzL9X1s0
PBOFGgGJlDP0NJWQu81ai5dDz9rUG9pK0RekBcFEkHhW7On7yUVqEztg5YmG4lZWojRA6pfEmquZ
n7+lNfM3gNTBAgyabemYvxT7K1N7HWBnkRCq44YSLgZvmAQaOk0I+RremxZCt/z0M50ELPmZo7KN
Gs/dliu65EcvVzZBwVpuBVVVJwh7sgLcfzurXJEoQj+/JJOcQx+ThcqJtf7Ao7CA3RHIQJaS8fwY
taNRIRFn3afZeeBnvSxKX1YgAWTU/gBH/3GNkauj4PNdG7JVJvFnjzVVAXyWYrl7BzhIwYiOmHMb
7500KZx1t6WLzGtEQam7RiZ/PJ+IwV0/x14IX2pFrqZ+km2iPin13vc/FD882G0Nr5vgogSB72Sz
Zg4Et2+4StwWFcB8amWX6cl22VCX3tvRunhXHjMY3nfCl1DiWJoAirTcod6HDm1lllGSefO6QR96
ei7XJkC5E5w2otve8O5wHwHrWY5JfysQX1l9vcxBe2icrmbTCL5crLX+tMLcV6ZprKJbudvXSOBX
fq2nolXpQtCOVtLaTGCpX9zW8WclDBpUUlSZzJkx3Y34nOqziwl0820jjnbJmHEVPh9X7qCJYP5W
0Og1LTXLzQHPnpYBgxSk6sLIWgZtFNDdEKSpXyK7FruiXNBj7iF0kZ9BhZhXa1VoVnkprsjWyUh3
IrhI2N/8WCzWABUPkkz+NVGzBOtobdiBL4ZbaGPaw36db5X92F6PeEO+JvwriM6ioBr2xtuhHIex
i7tUfOCfgbU+sjr+gLlDQdI4mrKtcROgO01LJ7ZRJ5nOe3j5UfZNWSP8umpa5N69evQ9uw8DZQkP
prky2pZiHxxl4aHgGfvD5iotXxMLPPCvzpGEBNzK+1Y2arB3oUqOWvdLi+7hDCJresoRVeUGVP4M
XWCGw3mvEetKpQgmL9xD4I+AsLGKoSwidIK4g1TsMg+dX30Sxx9P1yobUMgcdfXFVRd69sqvWDo6
4I3eAXKxqHA8fquhHetK/srMkDT6Fw11J+dxKsIJBfMgGIWmMlNdj2MoBZQan+DODjzr+HkbiDPy
+rdpiUgiSjEBKxzThA7BaZ1Arx/yBaEcZh7hvtcSc/40QH568/DJCQk7OF/vu6MHPv2Pvuxx93h6
BYZVHys2Ex6NknuMgCEI/98S8ADIUcz845VkU2Z3sJuYjUoZZ3uCtHiC5ju6JV1VR1IpnsfEdb/h
XiVsMBYEzHIiMS8Rl4Uf3/Ulflec9EfhPYJkO/2K6zz/vBEOkcT3IElg0etNeV1J9Hml+abj8QKe
9SKwrfJrdB0hbhoBTibEZepEVR7o22q6fq5ywXeKhf6guhItHn/SYLAKtODDau0CnC/aV5i0/g30
c4VU755XqzrryueURskx7tiSzJNCU0xhcnUxLLR9ZDmj4ZhwHF38dRUCw8/NIpR68vxD65SWcE4/
uG2r7kOahQw8bzSmaSuLbE6NNFqtDqKIl8OM9tQZ3NpNOfZcnbHmUZHAra25aQkXOCq5XKCv5Oam
N6DS3wreIlkB7rVzS8hYfxYLsjkK/unwiViiYnntUOjrwnwe1UerHssGhYcPZE2hzH1Q2VbM8PVR
Y7vJ6hVIYXFDgojxFQs2fwhQbIVV0/lfiW7vxwmUyZEsjnKmDLH3gILwHja6MtkBtEpiS5S6tC8M
qEYS/eQ0H5MVCrIt0GwCM9YWkYWchnHB3cgVqmehU/BEyOPxIhL6ACMqRYpGIcbcCBRRyRrjYTC3
1xINhGG0emKG+NYAJ189RK5QRy55e5EyWtFxRCKiOtj78vR+je5BgrzWmr4O+O7pdAzc7RJ6Smc0
2ttxqr3nw9YxwcvKue00olBZ/q5gvebtOK0MwCOFQoDAgbfaB2kgLFCqme1kdIh485Aiyx5QP3KT
JmQQ0UM6Z/l25UZHg/thIPkVAec5Fjo2uaEHW7lohwO2YC1GVvXDcYJi2u3FWtZHMJNqzr7oDVtz
nC8SRQ6Dgf6rDJv4LxWk12qym5+PynfXluWJAmIYjAKbVZXcCo/aIMGaI5HeZX7apZqof/4octJg
nujTAcRKQRWqdYaXw3Oo3bPvNYbgmonNxswuVAIuDlXLg8Gk0PVyeC8w2ch5rZYnyC9r8DcLxIUH
CTh7heg7GDShPuadl15UwxyKdbsERzpY96ECTuMdFI0ZMB2u8bgNLgINck3Wa+XbA9w6hzvCewJG
tLUXU29FQPjBf3257cmVrPUjtC5PI56ogBoS3/WbIxXIIWp40KIp5GoOINnQ3APlMUi5DHxUQXIL
hcfIGZSBXCG8zd/lmcnosmO0mhasbGIrk72FNHhgPqih8d6HtyttetdaflaqiPrQVHvZEIM5huu2
YS/ln26AHjb4EDo2yCdhkOzVrnAvL3vNUtr9bOlnrJzpZ1d3ttUjRrkU1moXDD2CqwYRGCFXlDwt
legDv6gu6quCheFtVOeb5rT8EtnklReAzk1RfTNIejXs9hO1B+6vfdW7rA7IhJkxPkhHtz11X4+z
3BNbO7HMMwh80hS+R6f/M96qWj5offaqqJgmmPgNRbAp+tQri1I2Zwgmi0zemRBrc0/X9suRzZG6
60HEoRAL8tV3T3nfwnB2dL5OGwoFrULQILudpSYpgkIw/OVQVEDqFYU7OIfzE29dipJq2e8T0NBf
NIxG2MmIF2u0tcMgEOwKjR1UhrM6ALl4vd5j07gDUXkRAOAkeGX5SBsPsb/3LK7IGuD01JJDiNj4
slN/QU80s+O+b4nM5ZxZgoadSuMw6UJagHGy75rE8N27+QBV+Ln6I7KBxo44LWnl/JwTPrS82Muu
QjSjrimSxcpRsTSf2hPzwGbO1NRxf0xyUaConV4vDTgskI6e0SBnbHbsLUHG8Gs7WiPWzSoAwTxG
qKleb03gNmrL34W8X1jSmkXOgXQAx0hg4LgtUUjgvqEUMwR4F1t+HtA5/2jqn04tUeONfPUXpOfY
6sV6m6bvXX6SyAdnHjgoJHAUwWderKjqNCjQVuV4pYfVb2fmYkrRScutIty2TDkX8shmlU+qRreW
a1mSG7ZvM9UYtFUTuF9Xp5xfAaqlscru/0DHACTJlXh5gUGEr23WaZbdkgnAf2JdR0eRWqW//V5J
KlawGOee+F3DtRdkjAhjOKBJYxMqCtkRglGZHzuQoMVk+CiGUKd26vePSyT7KWdXsUOo7yipoWDr
kam7D6ZPzR0kjtIS9CnAT55pBaNHul4KVHo3k+bwRheC0jojSSAloS1Bk/F52MQe9EBtG+njH5Vp
HuElgPPsi3HgpmSrboZVdvjoybhC/J9UKkGHu7OaA7eoWN4fxn6ZFdfTAZMRd2c+leSQePwJbB8F
OPQzbbYqGyUUlD8twkubFl8HKH0aBRii/Dkyu008NoM3QGOjsPMngIPtRXs2yvOTM19mGSzkiOAn
LJWZbir9LRK/0NpUD1i/Fuj83p65Abq4r+RPj0pHoHom+vL+9VZI/I3N9nUOqnTD/2KmMBZ419WM
rEL3CuDWziUfCLMjuhKxaHu6cnaT+ZdRW5vKWcTg5b2Vp8EMW4uXbXUNE7XSatMzlGbA/jtuHiTc
Bf3gE32vpodfIjUx71rLGXJe+dZK8WJGSiyRlGWAi1wK3OJFoKy7TfKq2NIx228lxMy83yh1n1jl
IAW6hBgHCa0L9O6O86+b9M7/HdIjYSsTJk3BvEH4fQzdBO3xniaEecVnj0iUmh6aiWu0luFwzql2
ME2CsJLXQXnC0QPjkoqtDkDAkSJiq2hLEJ47Ln2my5r9/3R6j9VkBwpkrFHOSpXX+HCDTKf7xvUr
YhzCsbpVHljelxmn9BjhfLesGatqIhhU/twoRTrBa3+RrlDUR1reeofpp05eQN92wn62eRBI85iA
i8rdwxhJTTWjl5buJ388WVfmXx+VB61mZFFO05sJo/hF99IFwxxsSg7x4AenfxhAcZlXB+E+1Ipi
qKjGTGp5ljimJNltBD0ims/XKQMTexW5OJtBgxzWMY1zGyRC30tG3YI/3K5ylBxGGVXWQkqU5k4o
TrX618hIJkED/OInAZguXz/E5BNmGJ1nNoJSYEyNKnplerUkD7sBAjjkG2FRLM1A8AOw3QzL8+Bt
41BtDuf4WFPtCuuFEejFgN8Hwh/UT4SxWU0gEBo5H6YvrPqaDSROPo9Wfc+jRqL6kpuB7AQKyUbh
4ZRJuys5ce/Cv1FpziGCLHUaR7GnMu9nYBISbkIHHXiUF/cvUbdcWrveW6buPfI+axuqi3xdvF9Q
FsHadL8cavNksivraj1tj8U8BMTJfQzobTzCRarhgwhpG3SF2CnknpWaC4ZWsdzHqLfbWPhTQAUf
SGPyY5/RkOzbtHT/goGb1BP+qhKwya8vqItVsqnmSOog/aOuwx5mDmhfdUp5pJUE74RdA/nj9ZiL
OY2WFErlm1/cAPpoqxobwTucD1sSpxm4v4DrVh1Vhi2RTJpbAUCiARB5RwspBIFFMtinFVzzhU/e
XAH2a2jfn5ZJ3hTlSD5Vnrx+dxvNaGyfMVM6m1RZ028uA20PB7kgfcYof5wOP2uRcSgTreMcnmxo
HZLzu2R10HgF/mAgw+8NVTBlPWEeGjysjzw4elMEd9jBY6PZnh6eW4RVAjG5fQngyTLrJmsHgdt4
6Tz0NBQb8W9JGjyLbi/Oz+Bxy5pUtkF4Q4yobyX1UYHcgFaeCGnTHVCXwPqCkH+bVRhb8QGzoz/4
20UASe91b1yRRHvv3BBQjRga90eDe6gB/tgAkZEuyyewkwEIPPWYMjSXu7HRedEICF/hHO2g4tXM
HVh2gJyhrETSvFj7rXEA+ccWkhfpoDHckrtDgGbmeRYDgP7hHcAina5qffxdsi/R1WSECtvSXrU2
u26VRKqFxKEXa6yF7UagHFzUcCiZ1azxavLghhaZleEN8hHbjxDG8ZUxOiE9ADvWgR6mdd5phnCO
RoCFMJ6+EZzOY45YXIckdBV6iht7EpOx4RM4gSqSN+36jVz76HURa70YzAHLtSVz4xZ+E50DMiWa
tfoA8bp+98vs9TNwQ9o+cb37s4ErwMF8X8uh7zj8/LMm5l5vRdMe8/HTz5rckXiFgctA3ugU9aXX
ujyjBEecOudESC362YkkwZzeUZbeHl+szNWXq/tm+x+V4wczJZHbcAcfAz9kFWpykIoSzL3qasjo
CdX9siugzW7F+MwUA8nWf3MSCmDNOe+1H9ckvZjg1yQNk3JBnq6eOQgtQn+2m2Ys5mhK4KP+4epP
O0V1PJRwOi03gAZkWDCLj07M20H2eYYpo1E32vb5NYkUj95YmkFhVw7cudVwBUeXGajlsGrN5p+q
2nHsaDPjhSixBavKIp5J5YLSErycTOIVGiO1hCJ40mdGjeydMwXRHXZoCpV6G17p0kd+sZJOCz+7
WxP4VgURuwMB1/G3zJ+8CaO3iW4xVUjjwsrkqAa4RW1r7siywkti4gcEJHxKC6MoUQiT+QA9tVtF
KOtg+ejBaATYh94s3cMXsldCa3WkVmZcELcvwMQfjyvVD+gXUw60JwzM/5H0QOVUoQtHqMz5BbVH
ykx7hiEt0vN/j1ZZAkJUmaHF4IBdYnAO8WldcrTfFbOOzdc83whhfTbbLV4f3dJEpodPj+Xw7H0P
DNh3O3vXoH/DyTkSqaKfPWeJ0rKMsM7EmLCvIZ0eGu+IWiHYIKbKIPV2J5pNS2G0ILYYgasKENud
9Ij8VKV4Kflh/7pzq7yyfCrUQkzw3TCNM8UoRxqnFqTPvNsjGjdnfrmvyJL79+Exd2K6ZfwOh/Mz
jrCGEFewjKFeLpKd1ze6HXATF9yKviUqRixwrN0TlWiImraMSiclt2JDRUIzLa1Yp6gjtRSYphCK
W5lUQa8J44KvkFE1idyLTAXkcIkqT3IBhWmHijpRDQ3CM2Oob6KzfGXs7A5EAd8FH7gkBW775FYz
Bvr4t+1nuLyjrfJoDAT52Yym0HFU9fZCcfgV3KTC8dgCkWJ0P9puLKxAkljk45yUKinirsxZlL/b
yZkjLiy2qar66yFxcpdwAUcE8FweCgx0r/op3WMxa4g/Vmlmg3OVSSpgfVlcGtx73QHU5wzfssMu
Hi5eP46odg7eNrS2ptTKd/6R+l/KMysGlr5xXOg08XAk7z2Xe0u3RRFxMGlYxlGjPZCea+4iRT0o
mnO2lNM3t3PrvD7L/HXtFQv+Qvggqbn6BGPfcuLlZ9iv/WeuqGnhtA/HDNUfZROUO5t4rlVSCkRT
BVmmHlG9+PN5J+9yJ1r/suS4nHSbw92BHMRgV7GyC3Td0SZqulHRM0j9SSr+aS3PGAM0yBNp3AQE
B5QOoZ96nHCR1/0x2s+G8KlM78jeGYsy9/JCdzCe//FEbjZg7WC6fC7wk4BQ9jaABNOKwbbWt6/x
/jEsWnEAec1tfxSbDwJTdNmzFBGzaO3Y2IeuQ93YSMlqZG+HfuUkjvrPabV7BSi4LoO6ZW3eV2Kl
rW/EKkFEw9e31fOm6EqGpjEF6sFw+vhA5lApOnZ8dSrIOxWzqD4EEfQqCCKqkLxKskk4130t6P3k
ti9DR3b1gfkvFNVADiQAfpHB1i4AHggL0D2xm0CBA+HstJumj1C1PW98qNdXAW+7PDEOCBSycw6C
TdPgPN0h4FG8z2ZuXOe9KEeOh+s5TEYOHT0Haq+yI39aLrUeT97c0rnpVItzwTEALFivemCbDfY+
h0QqnHnhYH/t07J/dT5F6fr1hdSGs3dxpiU7CAw9GsVIgOv7BhS/6B4SXvYItoSLXdmxexzHGRyt
jaKCgERzduzV/cJJzK+UnKV0R6TYMMnqskuWmxe7lwVg0iwTa+SBf/5FtIR/pa7IfmF4cwNaaDsA
wfrdLXVkuhOyYuM9zL0bU4heiYhwIrEZxfpVkmSuhR29AsVirr6enmbpk2HUEvO+r6WnZ8GUYaBl
fXd7Hs92DCkUa21gcwM7c/INCMoDzTSRSCaUUGwO6vFoTCpTPC8XuJA3BgvUzIjlABxf/Ekw3me/
whzJsN6/gbHPwx7aAJ3ttdmH50R2w674WPgxSx/QPHHDs9NQtNafIbOTsG0gl7Gn/CF2841ri2SI
IjqM0zzCcYtxmzGUj/rru8D14/jRtZ0DG/uxoozh9Ksvkdoko+ng35e4G0gw6CIhOyjAR89qSelz
uSvF1bf5Xg8OLtUK5andFxUL6/+NbprxDLiZFj9Z2wRl8F+mquknzbPv7SjQgVWrFNvGESYXaH5x
JY4THZnf9zGh/Y6dWyFbh/tNJ6veIb70aD6Xnic/F2YTQoMS28xBrgQ7mOszRewJM/5ZpE144vw3
kuUjRMM6xcp3Dk0AXdwXQ9TGmwGohM6nhmtwa4asYDHX2mQYJul84t3r1HMWsOkTBy8KIvLrZbLI
BXsh2gEzFyuLi0Qre/agmWUV9YsCsmDiA4uNLSafDXv+ufwsvmZBAmDqZZhqfNcF0KK3cLtbGpIq
871U3BQuV2kU8iIbQf295Kdd3p1BhufsFKwEij51JhWRLvGTvQVG7nwDaSKL13PfEN7IR3MEDhs+
lLw4Ie2ptb4JHMNm++TXP++iCX5CfThK4SP+dJlgDVEMwlgorsAFoeG23a2AAgU3v6FhJwyum9el
5Bd8/384hyTWw2KI+O9RrFyH9OvS0iau1mmhVSdH0qTitpk+zQGAp6qXpSBex8BPP6tTslpTiJhA
/mBouhhsvCCK80pov07VrdsHGcVnWRDLhzUXMc2fsi1blVpZXxTQnkF0pD/nPahPFEAZ7in9SxlM
hQMpg4WGjWO74KsuO/qfyuYY/xMsOfGHaj0Z1fi4hqikAevqGkanr9rYfCikojJDm87vubNhgSDZ
uIoqFkweRU6bmreUxQ/mXLQpQWbTimz06z3FNP21nZ6FakjWAM4BajQ0GXMRsZYXBNWjpJLP66pj
Q5m8QA7kOZhoFr0i72xMjNYa3Gzu5z39JjFRoWeqFhIRa4C9aT1Zh1FPUe3zlGE+r2hnqK4yTC9G
95PVRlpNCNckCk2KUa1SnjO+HLes+u2uARf3SS/4RPCkxL0fj3UIYSJ/H7xNGT+qUiE95fUaO/sG
S/hJBnAm1ZgQybISxbY6C5fzUE7ahWV6KyjvY0OKwGtvPG4+sr2ml8jmBB+94eypS+Z7MAeyWTgu
Y7N3yquSwVHTbaqJCc1FXxpQ80vYPP25ZZo/lqtzuGJsvRdsE5goR4YIk1VdAFn09hogjUCo0+oo
p+wMwBJN+OelumkoOXVQ3yaahyXZyJkIJowX5XuX+a5A5pCrLEPYh940gTjP7GTr2JMEB14IkL+G
6GxRWXfJWs4vZ1RPh8foIB6W0rfiVeJq2r+7r2hGqYzQzLkc2tDy2ILGbuoFDV3SGuLNsCyZEZa4
nrXJ6AKoUPhAPPvXAVSz40NsVMI3NHMY9i4s8b5MiAFkor2ZJSXDan89qCtIfjfLwxWlAiytD6W5
Z62hzFm5PvH/0qHisWVyV3LRmkf9QQ/1xvekVlaJWycxEYjJrGBLvivOpr0NXJS+Z80i1Ixex5x4
6anXwJBKXV847Ev7mf7XdBAjMBlZM2vjm7GH1bMxiC4ISvO2JfH3O0FH9QVuEAVbi2VnDlz7A0bp
zQVLi3kHk+077O0XTSKaiLnWdtajF6cZ46liP5D+L6q5hvhhwW1/JwarLUT8i6X4gztdsuAZPJye
SSP0lj1+dT8TpLRMoYYpr9VJbdpr6MDb7xhjoUp6s3s3EYLOE03MdD/w8NQU0FIo79gTmxsaMVQ5
qFkLaasNakli8gZiqHmQMzLl5Yfint6OhvJmAuS9HFX1Fq1wJN8DY7HC8eDGhkeC8Cyd6Z+y5k8t
15VNq2UG2hEfveqWFibxkp1bGvc+5/kCC4Pydi8HcL0GnZ6lYtlpfuSCnW3MnB4NFjfFH03yZo7m
HoTY/MeDR/Iu556WVchJs4+MHqlsq1i/7tCRH8Auqzsh+bjPpGy/gDEuMSxedNPbdRkFhm87vssR
oWv3zb4ocqN1ncsj5tZRQqdbtEoufxw9/3Zkf06uDhNb0xEJtzO+Zu3UO4CICAWE2o6BQiP7EIeL
6Gn+VdG1WWNkvVhKBzB6gILUJOdiRQWHgK7VFq9TLfciJTFasdx3hbiJEWYZeCOjaAmiNyKE3zd5
Njq1jaRMsOWRxCvUNk9KBygQgaX2sCh2mOBSsRr7ZOpwD235RK622fZ6OGBmnrBmfTOU5UyENxxW
L8KK4T08ETJ4bnUCAvwDS0vYN7slKk5ekVNV+jt8nU1oQEZSLfK8sVad2TF/1izdNjm4q93IOXZq
x35uGASgJrkPTLPrSzXSSfbiq+JuPiDtfTySCPVwCFLi0IOe5ii8cHq2en02FqVpeATlzt1Q1ubD
UhumOeUDPHfn4V/T4Wm5JA1xA4KewUsu+Rlc1D+kQbqdB3Qf2Jf0qcXy9qyz+HGRKRsBpJAUGRgg
swY++voc5UsbcTgMp8xR7brKqVgJb/X5VOztJLbzaauxdXrGxzVTazO/eFOPW8MV9w/yvHtpfp3+
Z5Rmf29RPBRyRf5Azc9ML+IRazd/vSgdyGkKwXk1PjrdyQS4GKAFhrxgsVQaPBuM5Q41MVWufEhL
6Mt51lgSXJf9024mewfvSh6RB2cPmtBWbZ9C0caKmtzXBzbhBDw9lTvUK09vWHhSSJ6Apk1LNayi
M3SnPWbMxpaeQiO3LCR91YT4A7zWb3rzwm2lPoL/DtdFe5HjXwQ9Y3ZA3CPQ7yCvyLnQ/dqP6JVq
UY+eT+KGJeDxHbZCRKAfKEBGDBlTMmMApHPFfezz+ei7LJEacMd6HKPNLhZHYmhUC98Dw/dZ/3Ds
/frWDRsMhu5TdbBDrO4hoOoNkm52Znp585hl4Je+Sby+AfP++C22Q/cCitnMYap3ZMvKW7uQCOyI
r2wKS4nEc9fVSkbUDDnmvtNkQAlJsw6OimIIrJ2WlUgHDaIymI5sq3CMOK67j8Bm8wmyf1d0zAW6
/QMJn8cnJVGEzMkuTPNPUV24JcRYQZlBjyMEvBCCDMRjuFLVFXCIzc36/nyOvJH6E6OAZWdombqq
Ho8+jHbc3BQGP4R1udC17ZgK4Ql/hbXyEhuZ0Obr6jjnZo+9NKFqRd7z+7rwCHLgutKVUIs4ksZJ
ypxwZngqFFLwJvlvoa48L5VxxjHOkld7olTYzXtAQY3TCL6K/ISHBrBr5WQiYFPIrNLZN+DrlUY2
zftq7J745B2BAIA7+CZyipq3HEOtV/02ICM0ViByE6E5jte5ykiMVe2jKSW3hHjVlpNgSRsT68kr
JpAO8HVLuh6/M//3fJUuuP/xeNSZNr9K9qjEJe5mFzrLbLGX6SZGlUFcJAlBcnun40ZpCx6eaq9f
/S4GLseKiAf9/H7Js6bf+BZshrspaWaO7hjDOeP4uhnHdT6202VhY69wK8EJ+JtdOMvBQx7ZKYoy
ArqKfP19zgFC6wNyT5ui/euh6L4d5hp6vFEmCXw5NGVamHdAccGzCFDjTxByAwI0LZXxmFhleHmT
MKOSGoISPT8CeTHhA+SAkEPVzXk5ef2EN2B37goQEvHHDqSIbIakRq2cwlhio1HxB80JqtQbHspb
h9mp9DCD4gBk69jiH6BbqUMJmIeuIG0AKG9J1XctrUxubZANHtfntIs5WO7Kq7jLRxIXNfs7F/no
V31q72iRNq5rgvK0bub8RyXW6gljsmyTdue4ZZZFlsfSda3QguSi7+6vESYBEF+1HKuYXy/GH921
3hzDn3qSogIrlTk5+afkBZrAEnj7ZlG5zmZSLDoOce86rq9MxiuqYKVxSQ8/Uf2QE2JN30hC9Sne
DgRPZF93sJDRwitJascglqyJda/E5RAEGxvyB3SOAtCJy+5vqvOx5UKfuLPNo47q3jQKN5TyfeWP
gd6KcNcl6132CUuiXKw9R8qobHy6PjOepkPo5IiRg8wYZ6A07Zb/N0zw+rANlpsuK5JRXGvBbmRu
bug8Ed4AN61sfC50oOjHvao/5sY6CHRcu2QakdcUBqbrwT2EsGNPLdxPhUhJYeXj8yFHUJ5V9W6g
t2kFIiwJvjG1YX86OmsgfxtetziUNZwQZn5KGzmg7UuUcgg59QhuMNYPwzprwbHFcS+GNyRlavKH
T6dlKcIXi8Uub4I5C+CaLmoU9Huu8xOCaagN39NXAJjgE5RZjEQpWf1gPIjvjno3GcfbitQ+3vG7
XTfMHNr+4pRvIyFQmG22aP7QnqMs4sRWCViyzGgF53sjIzTwez0hnyhF+taBrcwgvCrohdfLu/YH
05Q0HXdxlbHmuT3Zbehd24b9nEVlO+c22krkncxi91wFwIIRa3Y3y65SXiRUYiE6OJMaJULOLKqt
2Wyq+eam8FGFfDdOzrVD8bNKtttomxpEYasl7LtTiH1dCKo5XbAT/5Dv0A339tlrOMzp8eFyWWPM
u5cuK/aJuanNZXa4VU5r0r5/1flCnJm50Gz+cdk/GcTV+yMYFtFS7fs99j3SPt5TISCTKjFeuZXf
3oN5ILb816p0OiKVgDQDXVxSt0UdjUmyKBNBOC1rRpWg5rYn00nQIhVJF1CXJ6visnYCRW71/f2i
R7qiILnOhPLjbX9KMmqQ5ownZvAPwHcQlOAfo5bsPhpv0xx4TBSnidZWXh4n3gHX5MCOjyRJ67iH
tLJuEHvq+rp8DsG1edBqb4xVoXqRS/2OnBRUvz1eOUjyuUWvawNXXmtLL+MVZ56nYQRGmOxrsDDg
o1O4l2fTNoIarUiKdvZA2KMDMG+4+i5D2QepfUUB2tFeCqlq30LvJAOQE61+jAZQaXJAMPx5SVdI
onXoAb1EJbRJMb+kWkvkVHL43drX6TVMg3H/czYCkXn4FoQx4ncWOEmB6AmJ/Js5Ki8kY/yXUQkO
BC1N+NsOnSJh1yWCJVlfX4bnjmQMyrj3HgP3O2Y/lOmXunhlu0IYxx0GJ6On6p1IuipUdeweEOt6
H9VfiS5ovhLf1nFDvDdmbPwgvf06k0O1EIbHBpyX026hJY0w6wCOvDI0QTY0Mv9APjHvie+QdKtv
14BZhsi42Rmz+WZeX9A1RATG4sAjb0p/j5agrYS9FSs+6xTgbr7Yq0G+I8R0TrNDqKPOpBDMCvVe
1qb/T93C8o7RFOo0ubqKKv8nHoln5j0xLQeTwVOr9jjJwCmYXtMUhVJHzthcuruauahlOBOkZ8CR
yLpAErG4WglPWBapmIqKcmEvFyL4jqgjDUpEcBz2bvLu9zTEVU74Wy/50Fx6M6YAI+oaYOzdD/GR
0Qk9OA5M5qRKG7Ar6alJCZ2uahWQrto0Kfj9XWfaUMoqIWmLqFPnNpt6owSy79JkWtgq7sOMDeLH
qjqS9uLvnJLcGxVZu0yVLRiKx/yxIhc8Z5wgiQOlDTnaFfbluZrJQm46aS94Y4V9uADTdLMDyrZ+
pRTAwti/c/nTlqO3gAMPSbhiAwXnnyT52f6EfkzsX2fuFWCWigjU0AZRJxHXUtAnQi+jW5Tp6e2O
arUYXtN/uTgt7QlTFX2CdJ7yldgls/VHqTU1WnDiVayOXNMht63fCwD0z6hfr4mDF5DBhTA3Uu35
FSe0cATH4UnsD23oXRjZFx66HrA7Z9c2BF1z88nChxm+Z7Jljj0UCxqp8WXgGChxA02uHC35nSTM
iypQVTNjxKXkCRU6vz2jQwzzuOVQ0ZjECWNGlN5mdM7HgfEGyteYBmg6XwWmaPNiu91PzcksRyod
wgh8Yo9lt3h1v8DhOz48UiOZOZPBSn2X8tzpPM2Gkkwy3x2dGSvVDDhHy86r3ujOBx6adCu20z0Q
IU/WK+uYPU0Akv5lqvLCe9F8ph8+2y3zKsEGCVldW0wA37Tus8JYIrA8NGrKdmx6pO1TOrdvLP4h
PWBoJC784GjMRG99Q/hE+ACGPCxV/Roh7gE0VONqr6Pb8VPHj0nVCRrPZ11uGV5DLP8GePhjCdUS
RAYPouQwoG8PmnLU46fIwirFphTbjRS1gLFXivXorPBHd3WA8bxvfYEzOYt1ac9kIzSI6cYOEPoX
bz0tV4OtHXSp7/lWQxOKzW80ItPyCjNak+jQ/FJ0DbSpnehIw8JkP5vTk3/uz3Kczo334vp+lLGH
yynp2/SZo2NvnxdpOqJeaGSwMmli8/+uNouU8Tx75ayC8fjKCfLcIQzfdaY/58/t3j70ZwTvVzrg
we313iBSXa61v0vaWDrR8h4Jjn4wcQtvltE4ahsP8W0dWfa18fICPCAM4oXf5R9Lj6WczK5afI9L
xc1XWQFVso/b5Rzba4LxldKg2hkjpkIpl15z2643Yiuk5Uo3hLm6zadfrgWxdowBYVr49AbKBEJN
LPsbcNjw4p0OsWC9IZqA+ac+2hrEJjFW+fojY4Dh02THdT0ZZiMBhJwXWpCxDulAbQUs81MyQ+dU
Rn5FPa8K//NyD8F0ofVDb9++dCKzIzxUAI2Y7zLcw52rQa1FeBJe7iZKwke4n7BgZ2ooU3uev5zK
DWGEl/NZZ3SZorfTqbbWofazLt3j49eIqPJzjizMENjhMjjJaR9sdbbsFTvsI+PfzRw5MGFuusy5
Eb2m6lOjuVB7h1T2/rqmyizNESgq2u9/6YDBQtTMd8ryIV1gSvJqYsiYx3OKi8h1L60QWpH7VQZK
CttlUNBte6D1N8jNqAJ1FUs8gIgimc2m9eAfq9+rGWlQoHSqFop+Nocsqtkt0rydmt4kAdGPCOzL
fmvWf0q0TsN0NWThWWWCD7OSuIpm1miCCwTIIfywirKwLUmoDqOxLMEvqrTgr3G3uSeW67EUoEjc
YGofo4ORyYuN1FuJNt+DPgRALYz2aoY9bfTdVC5rQqql6hmylyQ1Dk+qTPR8Qs2Fv2b9XzH9IAFS
tARu2gbYxgIlhJoUAv+YfhHvfitlI+3Cg5g+hSot1y9I0zrYbNPNjZoLDKzkS2QGaGzjLvStTQOp
n9C5PaSMicDsWORrJYucpXHpSJLKXxO2Va2yFtW1VZzxF4n9tBeucfCR+ugLzE3TFUu3Xm8UkrLL
NzuGNS/ixoNlTl9mIx5iFhU3HHBpvx2y++oYnDz2VbRcqozEIlBPDjFLsrd2b++00v5GJQ1ep1wY
GfjWsPnveWopgshwOIs4wYK0ePCrV0blrEYrfNVBk2yFdxQ3xqDGUeHMVMuuPGuACVBu/OX7A4FC
2OLMa9iYX3odRQ7suuncknCTN6p+Ds0boSTgD/Xc3iR84ODGnsOSaleEZp/IR6KV4BgHky1tdopM
8VVQEXEbP48NXjCifrKq3LqATIXQfoGoqGJXu2difkW8vm4L0u9fVIBMXfRkTHD+wWoaH8Qd2vTZ
8cWn1+NTk8A6tJZcXHcwyIjJc3jucpOdOaXPkCU3axncRW+LgBFTarnQ/Pzd3bnGEBH+CYA7UHVz
vRS8AXRWhMR+HNT5DuoDx2aDBUo23QRB0Wirk++Fu4srsdYgnsDMJDe7qXkgXTVOi6bNqhkNeNjQ
5p5LLMLbZcIGd7TrMP0Pfu91OOsUWg/MlrfynIwjuL0ZxSaiMQi/gFr0HEHDmmvBS0f5DGrT5Hrw
KlFR5HWGC82zdZIB/zTzQ0lTLY6GvU5OQ3ieFMeI3R2b+mukZdLocYXSmadflhE//qebLi+E5Bi4
e8rpA5t6eNABKl18zf9AwljFygGGFOBMZ9LSa1JVXnvPCD3O2n8Uy6Vr7saa+AO+mkO5V8Fa9OTy
8X4wjMcETrnpwk7mUnlDRHIEC99DKqBbCdATa0nXhQgtPfDv1a14zgd8r0PsULL2DtBwjcdPyCJR
2dRTIxz2tZdfgouEIWWbk3NaApRMb6xULGudlpxNff6yaWk88yhLc9OTWw7fBaHt5/ZOzXwkKMfb
D9Up4St3q0bkrvfFFjAMwZqo1Wtx4A+NqkyFi8K6St3J/sitVBXEL8w9eQzanSfLNEwDBhL+qpuK
LIc32pAG39WgDRFywh4mc6mVWZBQXLf7EnF6TQI66c0ng3M9vBTrD3O/0l1q0vqXx9AsHVa7VS2T
/LiehWw0bRn84WbIUHlX8ka+tjOCqlez0kwUnALZ9zLisJ05kb2SCBdrEfEoTLvzbA+fFAcN9zsw
WJSpVRmzWxC3u7nFS51aeFcUCdjyMq084hX0J1DGPQo5beT8P5bceF8SKRGVVL37qQM393j6LeHw
XVcb+O6xCRUSHBekGo9jJaVaQwihob0ZyIze82iTwa+O9rs6OI2NU52Z/KfRaaIUt0LC/O9Cxavv
JOb5Ruu117nqfczJSOSIwRn9GNm+Ntiv1KAWlMJ96PST1afSYMNmHAKhroQouGU4pJs2bd/gSEG0
1fXdmc+IIne9Ca+c1K2jdUdyvu04v7As2hq4bw49EpHloyPi1OsVpTZd95lVf4DzdftXYnH6kqL4
lBGopnOBaR/tXj0ZsYAfhTcnGIV0OdmE4OfXdyO4hg0hJyd3XMtnX5miJGd2knszm+e4EKX5/riV
EUeMKPOxD9q12hq5bDXTe2l9TGXOIH0fQRv+uKYnfz2fjkX3+5PosqJbHB1r/macJJbkKR7k6gPF
dizdqJPmI632lck8Rhss9I2EeB84Pu5/gy5mIDti+8tevoeSaao6FaLFzDSLwSSEwM1tsc81Oc0o
5sbljmvrP+W/I7sXsxFLCmlfOBVHH/P0IuLvGeFeXk7Q1mLP4tcHseNfpT3XI9GErO/PhSR5m2s/
cqgQo94qO/NdalgMdEp1B2McSXnjKfK9sXBj2eKqEoz+ZprvFj7ZModHaPpzwPgfZf9GLdPkBg+t
1iu5WGoJCmuGkb2LuBqxj+hyiJsL6djaBrIr7kCyFUo0OkwO3JJQeUrqCXlYIzP8vMz/Shfvviso
rbOUeVCiYvRWU7GpuFLzj5s4V3WoW4GRJCk4T00sKBMgWAIFLMLhohQmWbThU9YXj08+Hlvy357Y
DHD9y5khNZJeJdQvV/2xO9po8xbxXM3NMfR1JkVDdejp++440yO/igmVPHtZP1tTAvb4pbfn6T/4
Kmiukl+au7YjmmI8hn+eQuH7+LpxAY+mmhcXuJEKU03CWOc/Sz2c/sG07zPq6eSDv6zxOKo/+Ith
e4jh0+/YcDNUZ056SRSoGaKhRQeJ8y5eeVJo6a9dva1HBFHbEw4QJcbA8jRZprF+hI3XUJ1tyeZ9
JkdU8sA9VR9p72ZlACtUdrrGj7YONhFe2XK6FVRD9FhCGwP7msvdUN7Fbz8oklS6sMfsXw2C8S9w
YCQ4OJ/its1MO8nGhjP3h7q0kKMVFWeM1R5xJbH7jAxTEh3qK32Pc+MuC5u8Eose7v67ptk7mAyB
BHltn8PwYwZGNCNI4Kfe568Vah/uc+eagr/1mOEuy5zb0adFPt2YrAsm5EYKtPl41vKq9+NtEjaV
HG3FGxGQl+0cRVeAzKMmJUGIexRMsqE36IoAa01ZAlrYHN/x/8S347Xzk9UMBURdFtK6mQmGS40l
H4JZji5slqFDronGGcbBGCVSjuGdDDmiExN6tduJB2yuOR8A6eYT3aJxtbZTLdCpGo4Wf1PjaHoY
AT04zbMUZ2jQp3ALEr+RY/fzHMd6MWf1BDKkrL+eCH+J/mZU1tLo8QfWjlJoJ4oxEkRTaTj6g5AZ
6fdogqc5fTw1YMTutO/o5oSQl/8S2/bAuYqM1+/zJzXB2VpghYtCpaDk/ZT8m7/Hao+0wVVKzhxX
0xE4nb6vJMm7uSfB91uzXP4zwhOFBnpIxREPpZCwJDVppc4ksvsy7ccxEi6BGrd2EHiPM5j1Deba
jaz5dMwsMICRuBUnMTbNMklkqplERz6Gqiqc8B9gCoQseOttwYJJHMuM77A0/jvI2iqR2CA/MvcX
tWTextTLhoo1SSHwe/0drzsjAuXkaO+7DE+WUOgEgufl4PmTTSfEZVi7ICf0krRytkVOYi775Uu4
rRWLbTvEFi+5pMcPa6jb9aLTx6ouJvo3wWrDlvyEIVGePOR4qqIJy7nXkMj4Ua0La7JB3dEOLUeh
nh7wa0JJBCK8udBc/Eii28dTuZdhWNAk6ssn3rbWaEdxTyPzFFKEczxlWYR/PZf0bpFrh0tKtIn5
UugIZVsLgTfqnLDeCTUbJRrhApY8sWpX7/Pgjaoirrv6cXEDpgWzTUSp/g8/nHLQKyJa7jCdY00D
UFqUFK+r7G4KPdHdbCq03cSFe+PuGyfbBYpN284hm6ra4x+dmZ3e4JUTlkXBodrZ6IM3S8H2B3qm
ucO3vMA0G+O3XDYk8iWupMw8Uqfy09HOkZlsPQ3466m9ge7PmAuQaw6AGMYdwUiO7sWK3doaLlof
d3o/ghhn+f4P1Qlvqp+3dn8RvOfBYZWNuBhpkqF2UN3/zkkx20bNL3ZvYDtdU7cVIVxNBVVpfICy
Nyw49L/zFaGvwvNJ/QXJMHgLf9P1CLyV/S8oxYKyc+XP0wq6YX05SpdXWB+CYvhP6v6Ah7+tUHPW
d/b9xnNlDEmYP0z8uDjqsQJmkgdZDSGl+/bwmKyebfWrx7OvBErGGK1+rFpvbWJuF3FPuhfxqzHf
PyyqSBrS68lo5NmYUJkLWktd6PJJ/Ggx5V7pLZ4xW9/6hBr1cN9UqhoeGaPwzZuCZUwVtCTfcNua
11b1aC1nuAoe4E40yM01BlS//da/Q4OzQJXQ3RHDTW+0uY0RjkFSInWFSgB7EAaqf5KMCnQpLlzb
YMgWrYUAcTKfG3WtBSvcvEbcYQgrZmzWiexNTD+clRx1tEkCciwN7C4RsnSMg2391ahEN+Ilb4gt
VmBZHoTVa0raNVSYMB9UpOn40cKK7CTqzXdKERkcMJHEWvfV+yKI0ev3shVhT263/4WOo8j5fMg+
Y8AKKMeExH1AbZ5/o19tP/EmlPcwoMCCJzo2QL6jMV+UjMh1qzLojdecNZb2AKhrQ6fnzBaXBv+B
53+HQl58vn3Rj/HAXoqEJ/G6ixUqU3WufdjQpWw3vtL3pW4WNiZAd6j/OUE0CMdrHnhH0WHkl4Lh
ztr6aK8gHe9zVjgX576MVCRaSI8pin4riIJITR7rtVk1Vsd6Y/9ts2Yf826eJwTbWB0n/j+9PR86
RRlIfRdTq2pT5N4tDXncl7j7s3H3MC2S4ojWeGDyPcacMYvtn3Vj4Xs4vKJfa1zFngyfq7adgesG
YtJN14ShFgQ1bjafHo1Y3uxt6RVDNWB9ii4y3hgQgUv7Bi2eZOr/4IMgJZIN/GHyC5TyPCX3E1ZH
6gHSlicLLgfBogyVHrXtrcRSGw7nR5oDqJWB37CxTWzqKDnEPxqXoKG7hMt/hih9wFtWfvLmDlyZ
CwiQStv7myG9kORr/+Xtq1WHBV9xuaTCaxgaxmGml6lx9yxA/b0K1tAqtWg0M6ZwBbd2+n+JumPv
tr+4SdmFrlpgds8BQQzM7ojCJ02kaE3jP9g7qlPb9/ANQ+lFv9Nz07oMrbIHupbw1jVO5NjL7iJA
GZKxuPyIyWScY8959hFfKQ/ykiIQFYG8B5E+JGkwdiMVmIyZQdb7Q1KJD/SzcB+1SLv82N42TXzD
RFuV4t2nauJHk8BOfbbfHqnp5lSPlabBfDjYHzM6mx7ZXb3tcgHphs8DMJz/boX3ic5P4sYgm7eW
1vwXfWWurNSvrw7IucNAn0BtlxEfuaHrOrvgTVzHped34IFKlza9TcoPbTK+k3t8A8lRzwm+J2uS
IdWwtuFvpoKvba4Wrob+/nFPgwsiSVZmLbzLw0rkMTjaCKTgdwhlnugizsy4mrAgMVUpSfEYNNbQ
gvD3nV46BRaZ8jJK+xnTRm6efxnaz8xOAzOIWR5NBw2YNdNoB8c1LVQMQBAl1zhRYak9zv/mfHm/
h02b5ZcWpBTLDytAAcAlB6AZ3OUd0afmmmF/clcB7Skjm0IVGAZMXyh4c9AhGIZ4c6pLBU8OfSTZ
IRTUYHRPofq+L6AlrWxDKTOmoAr+/tpciJ3xV1eNLUbAT8cCafK7UA4yFEZoWP3jPSaD9pq/kpZZ
MCsvsP5ankMFd/8uznfsW/JYslKu4XBeXQkDIjjBMVwCZbYEl/gw9O8+gvMHp3BlF44gPKNb+IFs
xweGz+uxhSYAFnaTShmmoXv5Wtb1VXH7NjtigzoK0oTNX96TNoqwonWeHRyJoy1N9JVkLBhuooLc
vl+2wy5HRHDGuW70U1mzKy2dUfNM/kbuJ78it59hNrk+DDvc472iv/7zEfkdDCdmjBVuQsh9Pyqj
tzxTccWaWpBuaZxiuhDKY3PY0WcsftHFE3hGgaXx5zwri6g2PvsKTKW945lTHdh+IsbKI6jwEQtL
q7ivYxGoNv/RZqRnSJWkN7QACWDCoTTmibQZl2sFqvMQLsaiskTXrBqt9QmbpuiNaYvKuppVYcFi
t6qpLCyFxN7oDvXsYVVIySH56xePyQQtpJ/M4IcjfSCUqS5/r9KHYV+dNy09JKBvBSsy383PzoJJ
Qsm7xNvIbObj9OjeNXw5TxVwU05ygNcSdpQb4/WgmIpvyD/KpsMDH8pUYsCsP3ylWEgSzyMomuQO
eeZE1GL5BX8WBY89XopllAa01O/LUv7robv2UTwXPzQWACymKg0LB+YTHu03xxXW+Y+t1cgmS9+J
YmsKuWPqsEeTXW+ZhleM4b4LSYnCZciWLnq8i7SLP5VnQRwcVoRaZVBPezA/EGBSus92sQKzfd5w
192DFUzLBicO4I6I7i+gtBAUsGgarOLzEU3ggXfnopVXYFYUF9c9GMNgYWds//2l4HXuUIGu0u+0
mUD6jsk8QCE3zHc5Yk++jIwv7zkFzgnv7G3IS4C19KG2KAGPkHqWXgx+0SxEaomHpzyHS7UlPZiU
+sdtKEJzPAZvz3gGr8bgTqQyYIhFIQ1pO62cxoNB8OfoldOHfq6IzQzFlzWmkg4lwr7j2f6QG3z6
F+H2F5vYVWphIONqgMToCN8InklRUDaKUezfA4Y+pQJ02AXHzFJEVZDszRyzY3HycRMdy+zs+Prt
44SNg31/PShT+jzdtDDVgs30x7yuCzQxgbystXK4KQPLPAoUgyA/lGqeGehfYwgWi2jjOa0lcGxs
jbO05eaT1ze1Cz7tWCIEmcWWzh1nRFxWJa4ctqxPJdXgDeqI9h4XmcW2ofH1qdQedzsfPBN7nTwu
qCyWNDkQvWjjiKLVMO6kkpI1qipiSRwW6ujkiwZ0SFyOE22c5uE4fqycRlVWrjPat51S1L5Bq2fT
5joA5eMdDvJopbh41tYbs4YFWad+rTVI3gX8zfGXis9aOUEctUP6dBkSQde3W0MuXNGwTjOd5u9B
dtv9BHktP9gzmevor+b/11YxQbpP8PKwqJu4B5EygaJpURI7dzPhDZeHD+lLfQsCB8TL34trPpbg
6iAgePUWWSIrnpm9yuNwwO+DWIgkgwwDJbcHEJ5yaJsCbWtNR3isqgxVkXMnI2sMO0OhEEvAnG5A
O+dre2bNRyLDpWnvq1aFK8aUt9J9DPphnVBQai27QraRJxmSo4mIxZ5xPUJ8XvGywDweQgQ267+3
2r/m87YgwzWQ7MFrJH1p6FHJUO0PGm7a1F2OAOoioV/hUE/Rr6ZkjkmM+m8NPDAfYMCVBBDqBDMO
rIXSeycva+5GAxL9fFPWI8iOFM3He+xjYyGXt0/d7LQ+PmHEkyZv0KBEzYyvqXnqwcuNYvaEYOK4
Be2nxYxDYl9Y4OgNzs/7OY3lbyal2JjZtsoRfjKtI8YQkiau2kT9nlj9H1dhz0CcOreSs5bo+qii
/1uraLfCheB8z/6mAnVg/f13No0Wwrbrk19N8uj+TAoqtFYYMJyZVUnHS1s2mofOhfJzTHOW5H7x
iMsw3n6TRijdmaF5I40ztRgOJe88hpR6WkOY/ZlXrBnlwJ5aCennCoomC/E4jbuvBYNEcZr3RgQ0
dKsvkKj0+hL+C2hbh6lOYz67jzW4nzJmSTccc5usTbCS1ctPNu9wNiO1oSzxaiScwDcExIiaiFzu
NbeS1yu/dKzy/TAvUSWUixD3vjjX0mIkLh+wdjlYuhuQubGQcPTtU33eNi5qb0PlAvwUcyTrLj5T
RHiSo/p7SNRDbV4KtdujJYAQ3gmV0Rhg7KZYtCbF8QkNHs9316mrzA7sXwKF4SNmDZ4aM+4GvSH6
VkD59s3gLOjPHm3s8Rkv4gYipj6/H+6MFaYWOqaYdlZTW6SnD4vCRhIQXssfqY5nhtFS2AUDbwc9
iyUg8NxQUx0pp9v7R5nGmXINusnPha+tLOyCURd4ZItfhM+DLI/w4h0PQSjqx1fMzVxY44ZtvtUE
ZE7asol0uBojEUrX4Pf+zQB/Ioy5wEIeYd2q7E/LmGs6yDimZ4aEsRwcftuiQ1zffUiR1CMV+5Cd
vLpEiLMC96upqRyQ8Kk6Rt/3HXkI2JyzpJAq8C43Wy5MIoPPDFrs3ENYFCd5/cEkDoz5fPVb/qRX
S68Ua6USaaU1XZ2E02qBGEsZpGQ1LxSlR54FOaR/vowHnzUEFFyQeC3dA6hRXBlXGt4Od+254yYi
KKFS6reEhh65dmED0elsytSZqo+EQImjMYYjsFBBQsVLPVQjUWE9l/6tf9QSaxrlRKvQxsp0Hd0U
oOJZF5rUhLvlDusz24bVc2b0hZYgKEcdPCN3/jx+ziGtWj8wsowdG/Cqc6qKT6ev2X3zyM241aMQ
P0ME52Ip73w6ltEg0eO6B3/y0KDb2l/3uEOBWUPJMxcugPzLC7TdhSpiUVhzyOsG9cP4uPBqRBCI
cgYSG6MfG+p1tSdgGRflnzLOICqb9n7dkqE6pd+xCqxdlVVpSYOKzrG8MHYRjoHcBgJUtGmAsP5w
bJCnj5Vek/x2qYHwj+CHwdJbx9GWzv2ho0JnC8ClGgeCgF7y9WAmQ+fESTQcGoq0hc/VjNcUS9VW
mr6XL//wpki+llJy61mExD3a6CJCbmsJYa1LTCW84CqMEClCupodDBRLPjLdPOZmW5/Og1j/WPCT
Hk+p989eWGgKPwHfMbzNXcPY2dSoyrDYnWbqpGV0L3w8zfioVJqkmEhIOwsHrr56rZC+UdYRus4E
8+VP/09UGcexT44J8Wqk869clCg7xxkD6sFi3q+ta/L6i52ddf9Z7gbjk2iRNaIIJQ+P4pQ9fnpR
yNInBxaQvaeVjJ/CxNHhcs29frWXQzvEv0u8YcaDqWkjHbVlBDnraXMerLVPdlWJRXD2gMQeGYjh
uIzt/XANrkTJ0GnBwoE5fISKJkRVj9no5n0WSMf2We5lPL9Li+2coT8hmATROZArQniXTKatqww6
QTzsDQQFleoO3oalLm8ALITfJGUq+IkvCPEmRc+YCfFLNbkDfjUyUagARGFn6RS02l+gCWPsoJeg
Yr+T37R+Hc3mb5BhQ0xtp7lThA2kXZUypmaTNJt2FJJIomInW+6kRYib4Ui18a29bCu98wo0mGNA
x9+A1SdBRbyzc0bfl7lNj+wM67gxDOapZAvx/z4GCkRif3Sz99jtLNtMgNAOwhLjG//brYFbi32g
J+XQ7+YnxflX7Nr4oSvA/T7EmhyeZqBz4BqJIjYnvwRpJI7AJEZ+UV4pJsYAEe+mlRQf2xnXfo/l
LlW5Uh6p01Wn9BzdnBUp+oMIGIzIfjAe9iS5ICFM0VB0kipHwqbU0h4zL/zmBYPR/rJXG96E6c48
ORMKOkGKgNz9CBMJ4SyN5dagFnc3SAg6/Naac/cIpZexP6ZeVsCKNLrxbHWeVw7i6LdXOVVvlMOu
HpLNG44+FAUCpBAa+Z+DuabqsWPC79QtRHavd24Z3/uDdgx8qx+SdejjDbgyoD3+qjpaCo4DziyX
x1xgli+kqPuhRL21Yf+eaAFT79rHWsyfAgDlleWExdHvZWCFjoDayHA2Vopd52+zsHbFsUqNxdtA
lzt0cFHp/NvlUg/HiVmqw6XRmv6zHG1R2iZhiW7BMeCChO1kj6FM2LwNauWURpMx8fTMNB9Rcp9S
c8hAzrGuz1XE20toe/KPOWgdiMnc8WW7JHZ+KYBTEEik6jEClQ8R7fGH/U5BZcc1seDRcpuOmZIe
R3PYjDedlFel7RgYCCBKIw76/9pIX6gttMU/H8ZyCuRji+d4xYgaJZdsgqW8jHmeNnxfLaBvuPZ6
FxLu8jmu7LlKhRaxp+BBPl5AwVXTKJJzS1hbp9saIZZAJpmG1h8le/T5M1UgrgEleeD0YNLThQwt
ulJTlLH2D0EvxYyJCqKmKX6+w43bUSrulYOheaVD3cWGYGtKQcUwxXF4SLVmtof56XSbApZ1obRZ
iqVmqe7VA0PzS/TjtGlAq35lOPJrQPxdmN8S1BWRqnKYKz1CDf0Kx+VDCZ26xuKaxLIEp7jLroOr
1YWCu2zZ1WpE6pNUzjriDQvxlp8THAP6CNSunMHTrSabQRMCtjPu/RvRMqwTr4OSZ9M1DDStHqH7
O3f8iNMqHE1V+3uLyP2O1D4uTCtk55lyAOJOkSeRACye4bN0aplrsQzPzmaPo3n55b5DaJOr+zyG
4Cho/l+2whmIUjQMZLEB7VihthOn+pc9eP9eVrE+eJ5E/TiArT35BQFF1btGxv9dc5I5i6yDXecc
Vj5meUXx9emGxqffSbjLtQRxXTZb7z9+rM37HbrCB3eJ0vl+JT5S5ge4uSBryJR2CNfAZhlX76TJ
iO8ZnccrMuEktvYqy5dOhI1Mf59GcD76jJ5Y24ye8rtIc+P3pMIcLO4TiflIZvI9ldIxmfQoga6a
VZfZ/pQnoT3l3nJTAeFsoIuBp5foqRkjEVa/xfOczX7WdkfdRqz2vGZZwkY1nfZlP5RB/H3kZ2Bn
25V85KSYGIoQEh+4EZD3YWRZG1gGXcj5A7pYvds8uVsAhw/t6jDF9Om+CXiDih0DsYF92Qw9oBVn
GnXD+loYHOMC0LjXu8yXzmhLhxUUUVcBBgoL86k36wfYX+0ylL6W/JECIHAa3Vxnc47Ale3WH3si
rgFHz7CeLrcjsu2Rg+OEZ60TiJaGrhZ3RchFrKP6UxWYhUfHL14mUIdvjOg7igS3tEkaaP89lAtI
ShJQMHUoBcGi6lo4jenOGR0qyVHxEE4AXcMayZUzyO2e+wWtit4frRZygAqSAViMTZKhuM4RrIcy
0ICRUzqW9zTpbSizafxkEx+thFDyHpSKMGrj7MuTMV6oxJcB45WNWJ0sSoju+QXSmIjzu03MmAOO
SXt5H+aU/IKCF3aJyxP8S07B/PiIytR/M5jJToQGAYm/Nf3L5xl/VNzDjy6TFCgPUI88XOBU7SOB
OHtTrXLXw13K/b6i1PyMx+HINGNM6qvrrm2GikvE4XIdBFBAz2fkbcqMaLkGixC9uYMn7xlHRjp1
irgvu5kYm/HxX8I457dfioifEWV2TV7rim3YOBSTRoIYQyTR4ie3DpNFpvnbU6XnU94L5h9uWX/0
NdgXUrhqycvysS/2c9hzBVaNnll5DC5BYFGi+14050vXkjcvwma0XHVdpkQObTNtnv5UIBO/rilx
ibcLjASXfZX0x7CabpWMJ6iC9NkJQGDzQAhme1t46ouexuzee+Ju3wXxDEHjnHZ9yyNtUmh6JGkP
jsXksaEyEROv0GOGn/0jj4IHD1wCJokRZudjXFNJiSRpIDX1vgOu+d64pRrbgs0AhHqXKvO8BtT3
bJ/P8TMKAlfyhU8ergHCezSNGmPH5jLVdDbFx56ChoMAIOzrDnc5uXMfsqGOIu0cyioC4vGXpy6C
HVjb5UZ3i4O+UI6mBRU4gQExlcLPRnDdBg4InIBvHahNYyD40FYRhrm146vYG237mGTsNoBLIwFQ
cy+1GSArVeFHX3U4sLE2tVuaFISfVr/HdSrI/ktTn5RilLAcvdP5xl/DyCO2Bvtf8ZSMfwYXZx6w
8RYYT4lmO/ow/mUvQ0+Q6yAIAlU2D//T4VVu38bL/BeRK2d4BxGZTP2slTtAx9nm97R4I9es+/Xm
xiJldOxmjKPRwxwjt0v5cLwkF+ga3n9VuZHBJ+yqJOFVbVI1y4hw8DlAwylbvydMhZl0ev4Dne5e
xJ9Y4kg7aj0wPSRSVzmB8ERyJYFbRGrU7/BUuSGC0igjcG9769uxx7jL3a+2kOg1gMtU5rsU1zjr
H3sJglXhsU3JljSNX3W5Bi3o6t8iVQBEODuUi9klHYnsnq7GLZV4KBYfh9LN9nyvJEaNlC9k+DP/
ruGg4Qx1KKXgLSaha+sxxXcC6vLxG5bQOp7F49/SjmtKX5Bd3NxhY+Y898XLhDhTUg6KlD4W7MZv
rinO7jwT1++IyGI1rQTwS6TQjPnejSUw6ntFL9xXZC1GsRgnHnQnWTiYJUa01QReHVGzFWg4+GdA
5tMrqbv4ykX9F0yYgc2Le3g5X7vzArvO42+Lhp7UmcRRrND25Mz3Nfl58iW1UVHtXARh62ThCrP3
GozP1rr2F9ZYOWIy3MJ+nKgx8Y/3byx1hJ9/irfLmCQ1Kik2OXlmZsldiAKGB1xrMugfOS8BqE5/
Y5HjDhpQWvlqbIQ/6RL/u4TqMc26o0yvQNEjk8jBIb9DOXA8iqkIQYx56EHjKlWz5eVWMesWOQdK
jq6c21/oErUe1hcvD035/Xhd33UIIyULSbmbEia9sPWNVMdp67VqgEjLzugl3lCd7FWUozkUFhd7
7zUN0kqMXxvbZWmrzVChjhW8Eb3AxoMKlpB7sgMbRt+IGB7ZzGLDFI7HV7vJTyBonhTY56O0nU/Q
DeHNL0YLDKztuHuwMEp/aDGAFMbkYErMjxIwTIrMp6gVQRj+03cRv6ohCoW0K3Kf9wc0JoXsgShX
mLGuPRWLNOZbBXXDInI9USuVVU8lMMIL8j+UoWY1bKFTe0DmG4pkMmHt7KXTY2ocgqfmjKWdic2Y
sKqizDzDP36foXDcBioHi87gxeY1+TOR051ydW6IAjjJXHt61aLDdLc0YAjn0GlYWPr7EhOA4ET/
um4ABNraFsGpUZxmIwaKWgAs2IH5Pshz8xZHVqa96W1nvkTOfrknorSa5y9Hu5VOizFf4yQ1Btml
hhAys4QnBdFhg58QMzcSQiWy9FIvaMpE7FtKBDFBOMKUmVSzWT1mblqcw+IvCG5AU5s2IgQI7+G9
8KtqypipLg7dk+V/DQytRG42GQvCU+naWB7w19dEXlmfUHjtOmsptV9xlIoyg2eSuDCi9Pf3AaG1
T2aBtjWPsPhNQzvmt9gJ4zJzuC7Cb9dfuRB0/AxFYE/06/E5PPr+5qChotyFSKFH7DwR0aIfnqDU
aNdQd6WXv8SVQCgk/lm2sQQBRtwPmwG29w/XxfAYdHA6dq318l+tSnOz3sWQbhSdIlzmwkfW/ITc
PltG7hIVfjKNFGSHbjk5MUKmqQELDuQkdJMsWseshF6areDLn7Su0E8LXBrcBwc6+2xYWkleaGn5
u9ie2EGb9lMcGOeReQcpz9ES+xEl4hpjkohCU4CU9CkcFviukzDdevhoAU2INb5Uk2L0dgf9u8qr
fyxKe2qP6PsVLtv0dKAJI40NAf2NPVQQZayUUlmDzcVybh87UQ3drItGMAtMOFsabC5ZDfk/BREB
hkjDnOa4NzWnPvxEh18+AIwXvYFkS7Yk0JJmPBeuhgQAgdFy8Tym+Qcpy1xxOdBHDbVujHKUqyOI
K8qq4XxNB27QGaM26EUbKsVhEz5giNaEINleOsDSWqGUMuAXWqaHKuDtsu+rnUDHkwtFJV9+u0pv
yMdO5jq4aksVSXbatZsWlN2LU6gAjpIL+r1EUD+6AB6K9a7RCt+nNP4bUVdrqgNFwXSyS2UjVY+q
cY+mTDv05bZSUprflo6nQC7c2z9TXXt1zm/VntvvIjllu1MXNomZ6ouwosOrd7J4UgoilZ88M23r
noy7NjNnsTO45b7+h/J2A50ZEtZCmf2Lo2MSxjwnSwLfjcgPhEfO7vwUmUPjWVgcqxvtK3AkcxbL
/8rRYpwc18l7K4bCJTKXRKjX9p7cmCoIj7OjG+LMUopKfUX3T0p0G5dXqL0qnMXdOHbcxROY54lA
Zteo6d6QPFU/kJqypLMMmFpxiSZG9ItujA4OGNT+0GE3+qluY94Ti3a+5yOo3LyEu/RG82LdVRVO
Ob0q9z1hv605refu8ExNhQdSZj0xxcvJsFd6jDdug+RseFbnCxNunrcMCT5+RZBsAqXpcMSImomD
2nxlLrx92RXbC1BxM+WdPuldFwOMU+fT3ujyUc7igaJf7YAdKbATOGtwa4sXpzJsfCZcX4qdFP0B
jeMxFCxN3Y0p7oBbGNgIbzTBGqXtuYXtAf+fkuVHG3L+Ud2WUYn4hLY/IYL5q6AUPIy7NKC9w2Qu
K9zImnyOzK1PP7J8Y+4hoEqHjNKmW2DLxa7ylULLRm3AV+VvNhusyPCAYPTu7Ljx0nn7borreAaW
ImLlsThtk3U4c1P3qLxyADLdlMGHf06kiQMRpLAF+Y26WNfWmSd3BKBjPI6bapbYUy6DTKzEpzhZ
9wrAExA+9DiptUpkqkYphZow3CtbSOhmJcCudTgnzDu98zh8o6B0RAhcx6qotQmeSR7kQuNLy5f8
k2cHlV/OPLxvqN1QGRr42L9AJqaM1I16quuPRdkHJG50SijJEOug26oZfjELwEWrOqQez/syIZ+k
gk6KDJbL9Ud7gp28O9MgEk5u6ae4KgCGc32kU6PacSTd10GUqb+exXHNq3P9dwU0dEA+8eCi7t+2
d/lUguL/r/1fecxFDbGPWpvrE33e5ZL2PNcP6Lt/gQrknWTvYb8lxwxqN1XpBxSPTTVP0rx05cjr
bbXEDkbylhVwzXeKCxr/BV6WCsKTGdS+yfeYYgjWpXOBfg7CwZAaQQqORewXRRgzH6mp6XRNWvC1
QJuTKGA6Ez/S1tgQJGqPtQ2AbmgbAtcGyrn4KfWXh8kP3k8/gBKfoXza44pblUa40tqx7LH14FPO
UIsfF98t1stfIBMG2kZbdz+u/kmWgzNCKb4cRoyluVomLTn5Z5kfNBgvZyc0Tj8UAl81pTizeCfn
TTVClOuhgRJrAWyRp+NbFnw8rbwF3dS8RlM3ZMAX4LxLx3GldKO47CS7Q2qvjTeEz/RgRLs2vdqF
hhV8stJrMyukd8MDSwMxGAsEe2kT+EnhaMjfjxatIyL0N5k75LtH8lKUnTB9gU7VuHIZozSMvXu9
jKUPHbyP7oSGqW0+csfFbHwTfJKZiQyqQ4TMVyO4zKnzojzgdGw5ROfj4UwKwpEYu0kBXRyYR/8m
gJWsUwnMuwkpy+SgRf0AUwrDtqzN+JnpttPrEiW6HuwG5jsSWWzISFtz7B6ACtKsD477jpZMkiTi
v94n7lrVaCz/ip9z/u/olaN6wWkH13ZrGPxp6hsX8ZnJqn/FaO11jww1VEZT5UBxmfnGAMsim1oY
1VwJNXVITyylzwQAU1cB1qCxSlI9Nbj4eeDUoaL89yrANygtRntIvFSpmtmDKh3YBT07cqyCb8ms
SRxmo+0C5tW0J4/yY65uuG7uvUNhWYCVzrhBqOjCjsi5t0nHaj+uJ/KkO3vtlXna+6khodWsHf6R
1B+9n9xW+mPiDUIWf02l8mYkzLcyb2X1oiHHEyZeq8HfDd9Awr+y0A4RNWmlPCR+gSjxxD4QKUCk
Bhddg4fkXDV4RuOK8RjDDZUhESdfmHXMrrnlkETRxFNZSZXj+tcXAJAgy8Fz/DGdrKog6yIgQA2a
XFwfdPu1B+T0B3TMrgusxhPaQnNMn5FPqAUHAVzX3nMM7tdchB7hFaJqObNU6PY1S6mniNtiSVYQ
Pcne76VwQQGMnBWZWpxFHTbXQOeUTYjh919W5pyxxrX5JpkOms08+BJL9nSrXQnRqsset/qAXkPF
coRk1WyT240kM4pIPJIF3PSkHdeoy5hK+UYMddPd/XJDlx4MSittgaO4jjH1KHQqJHu9TNEhtnii
nUQCg63tddEZz5NIUio/G7SDIuoMjedcNd0YvbaWC444cugap13IvfsiDmGrivSYZyXxVoBaLudD
X0ZHyZyROk0eznyRp9HBa7dNPmobGiQCGJfEdjTkxPNPaWkAXEpXaSXAlN6vJu7tMFEDRswNsj6I
CP6tZIJqaT60wS4wl+Ofjw9nm+1ufp8/ZC+O7rLJ53wSU6EvuKt3ibBP9J/FJ/p5TO+RjTR0EOFg
iO2oSWEsVzfIKEROg28xEQODbNGUp4FZrOTSC+tyDD33Ecam0PJVr78AosHjZ+cQlSacgxNFaCh6
fZ2THLRGZIvA2VG9VP0h8CUEfQxGS8VthqqE7fS6JAaQtZ1ACGqCXcjMtoS1t02DSpRWRT/GyXoF
IZX226gFEUCrxy+ovGUr8jUQxeE38Bv92ZLatLkzfPdb4QrG3KRVBwnP5LDnqKEGrm5GWP6DkB3m
/qkRKDlgDViddwtUPIj72QhfZMoBagSPLa59RNRCzQA1NtSmtgnOCe9gTTbv0M3sZvclmzgJRLij
bi1H6FFe6set3iZPWqVxFmD2KAhZNcT1WgkRjeOTfXKzRHnY83F0ZA0gjuMXTTQIq/0Ma71F2mgA
tAX3tJxfKbv3uBnXtimuU56S10V/o/biD9KfDYuoa1fb477brnZ3nOQ/YJnayGNL3xddRzCxJI4e
8Kjv/ObOBIsrL8gY9zoCLWgGlQMPkkh6CVMVrMdycdvyybgMVb0MjFjns95S/HJf7HGiI11pPNSy
iHxCOWENrh4L7ma0XPhsZpBZo98b6ESbNSNqL7z6hUoBjF6LeY2qvDB5naPIWzAlTEIrxfljf+HE
XmbVtwfXEV6EgthCzsMP74qxG8rNFp4CEHppr8gryTqvCQ769P2oQgNY7O+BfRZFrY81kdbcgpNW
8zYWOyfwEoeag13y9G8iQ0i7PoHCGEVwK6+411dmbLWF4IP1grk4Y2Qn62OnGSA5HQ71BoEBaXSt
icPIM0nGkvP4IJROKY4dNNKLbWgFe5r8GV4MRlLO1VoV9GeiwuIpMlIyExhnD+L3uvRn7co/q2qm
RvE9aRz5lm7JKBZJCSJ5hVPqMujDqDc8Q1GU6/wftv4QEB4iVdf6cUCTZZm2hWVDG4RamYi7txrE
DUKAW1HyYEswESk7NAc3WBXL0/Ddw4ten4GvSpWfR1zKs4sABOL1RdUlclovHgpgGppFVyUfEHDR
+NL9YfZB30hWRaALgI5DvF6y1o7jKoJvzBzCDQJ7fm7R2lqIb0OnsgzRKxwWnSIoqQL8FsSHr2Aj
mgZ8asL+uygyBpYhCyZk/tr4Zaeif6FNIqPb0yTEh4g9a9uMj2PVawkgzAezwHr+cOxi/sQxKPrS
MYCYLFT648WfUupWGwm4rKbjnC+OlUTmru12SBPgjRAHoruXGGS1RqBazph8pMX3dZEKx/4fFwui
7fMct2pUyZYvuEi3JpztIqDafCZBZDz5cP0BPu/UGWITxxEF2LLV8TIN/VbqofEy5tjPX9oDocvw
VhvlytC7IfNM+cchhuEQZSKtPXb044QXBNA/UFoK7siNZHYUmr00pN+bCySd5ezCBZADaOcqz+hl
PBExJOqBomMFObSh0JoHmIx1JjKAxAQ6P3Wsa3pWcsYqHBkG70yfB5LOImTlmOfOOUDydZ5+gnZO
1ZbxmBz41n6N8dw2dFGRBtGY4zQPh9E1AjZetmKgAkpt0W1ulpyXVBjwwgN1Xl5FqQqudcum8EJV
DMYErUU/cJNbMOD89S8smtCpVvhEDltzn3hyciiVaFlsStqxEMBdHHHtUbw28oMakpAblhxQb6R3
2OtAelF+pZuOirk9eJWyj29O0nBtxT18VuXrpNcdyoITpwGTHiaeat7q9ce1rWn2j4R7u0htFCx8
WHhWAlexeuFiN9XT2UJaA6p+9JQsYut+p+lmSSP4j+/fuK76mpX6IxCnxeBsjZajmo2eV40e4JXO
T8ihmPLc9fFtfFJwVj84ccPWn3DYOLSAKS7vO5SewIu6SNAOuIGpGozIJMvTc0p/Lz2owJh9k4Ef
WHu0HS/xBsPBoLtVUcCeuXJI+mAqrbCxQyB/kBabafn2omyFqiL0HHV7X3n9hTz3y3DD3tzbyFsB
XT6sBfZeWYZmG+4iVHPrJ18eEtmNvZ7kVXsgObCEo4eCZ5I9xbpn1zA0sKT1BrGrdP3vbHXA/wfX
2pBahn3OfIB9H9yNyWgBi6Dx/0UOQ3f8mn4Pf1jTdRrvgNYAIZv1ffDyRx0v7ui9nM5Xki7PFUCr
fjy09CJyW2dWAOoxlRUEYfWqPjT1VIe5yYFU4MrS9Y5ymyMYV5Th8kBuROsnPjXDsbfbGezCB1Jz
HNB2VhzGSqjDPtY9VS2k5l/hb/6/umWSOr9DgKW7ONyr4hafLR/SwgARSR93W9xzgy7tOku7U4y6
cd0VpzNlSnADlrZ1H4SSAT6SNt1X9wLQzpntBGvpRRilhRiCjNF7kemBs7ol7GGmmHB0WCR+4zhq
dHnWi7qQbt7nE56U1sIYF5Jca46G4hjsv/PlxVK9BDr24hRCJC5JMYuuRXi7nYpCQMKxma84q+Yq
7+aDYSLFKlzGXGmdEd4InEICqt5BijSL47zoSSrWpimldUPcBXr7aOwPz2IEZyCSzaOOON9KBmQi
eC2/naFNVdtLimMd19BRQicoPV8NvUoKYf1MofraxIVSePid9hz3weA0+3SAVZrgHSItWoDV+N9k
9brFi8JDeVcKkyBIJ4TgiMlpHBoVkSyVf6iFcBaK5jUWNasMOiB9LrBkYBBxeX47BpJ5eF2s6rH0
2vvLrYvOf2h57OFmDHUxLrKJ+Dny7KroYLP8YcYF0q4n//93bzqgKqksZQOCzggrzhN3n2oNxrdp
LO1RrAV34vkajDew7IGo4yojDaAaCVa53w4UfL/PBDp333+Gl3JmJsBtvkmy3Bv+eKT5abnAdnsE
KqvUUIb3MqzmNawzt1Zt9LwMccI7r9jP4fW86uyd9d1NGrJDn+t0bc5/d2lHfy/I3hUoaX1+A7cZ
WW12LtlAKm9sZZQprknGi9WDWdlZB2QjFXUcop+bnlV0I2imp2C4+4s8xpsdq15S/o388et8QbIB
JRqVzUwJhSQFp5McRq5dzFfbJl8nIFFd3ZVrjFqaMo8ikKm1+/Pz+FnY2FEkcewSLwxkbY2peas3
5det6SGfrwUalszN72160hFJ0016dUplzVrQDVlNIso+Eex4QnfCnll1k6P7C5MJJLFdsg78MYOh
ZWL2juod7xawwvuovcT8RJjWehE8JWk7qvyFSJ2fzu6tmMr4d+tvpuJUE3ciXw1UnGG6yYLYqJnd
0Fp9vUSedh0evNz6NOkFJb55vFlbFzfo3IxiYqOMhhYNTOfZBRLKjNNPIDnHUtuSQfGKY6i8TK54
lpiJwbEgza+OeMH8NRvNanWntf4TeNC0XcUVaHaaa4Ssm2oWwEwIaL0gnMDCfU89u7sFPmEVnW5s
G5PNxFT3H7RNbDmTS/QjF7ZY5oERME7uFksZ9h1gsnB/ljy/IWuhg/d8HAPJdHHc85XIn1NWq0oi
ZfS7HLOowk/cHSQ2apx7oJO9/szQTRB+AaitmyJ6QmQbUeN+DVY6jVcyml1XHLD4mmgj7exTVTnq
p+hDfIphiR6mkNMz8SXpd9QgQKPZL/NIks/NxEX5nmZt4QbIxzrsQNyKMenMnmY9+Ww1qZc6y4Nq
DL5cFnyDUT41+gDNNiE5asoRmFPuD8g93SsFyUaIJwFij2wxDpmc/vycGaIAOg0hUFlHnPuVsDeX
bvuE1rXbchXZx3zUvjTOV+qpEBNoJ+mrQus0VLljyGuo3oxE3r4tMmceqGyL+cuZHi9g53oS+kNw
q+LbIZgIfd1pqnojwmtp4gsd+/r4SqOV/+BpdXrbzlhTtwaZ1vMWETUJ2rY1jSdfarmPkZ94qYTC
dUCt6ZzyVDJmvZ3b7dBUJmNYTFUujhKQV9TQkejf61LdKDc+CxoMQeKMl7+N4OcLYd9zL1tmo2Y7
izUFdmx2fvRdSvYYkIV1Y9v3z/6q5y+DbaqCaNrXHBUuhvjPKpVco1OpN4+GFT5qqfGcAOnsEMCk
NSX5fFnhEUvX1EO6y+WwEDRx10EwUbR4oT3bVa/SSThlyM+eb7DOMSspnEEIDB1OdD8rvJgB+hue
4S+flU2eworiiIxT+rJ/lWnc+p+uL84exMAcJS4rj9jS9U8+3Ga47JaqQSIadi/2LDxqFdKlTTkh
vKJhk+CAnTdIPdzRzfw0YM6fcopTsE0wepSaeXXFky3sGGZB8x3VQZvUwpn/coU53QBrB8s/h0iv
vb1mSRdfJhUiO0489i6a/Xz3Tj0zwdXD3X3XUztinc9dwcIqHGfsZZkt2CRT0+Tsbn13a2t2V/x3
P/J00JtoV+UqpZ1cL1ZTY1NJbpl0EGe7yD5pNxsylu9qq4GHN0SNGIWWwDoW9tGymLdAROAmQO9Z
/3+C6GR9zNIbVek/4qLcbr/1yrKG9m3zDiaAZu9tjsyqOiTCC/g5wTcMewpCKu8YYXT/PsfLfI86
YrWJAQK4/R/VN8NCCXGGhiJNrfrCYFT1cG9sp754Awx2I2Z29BI3PgdPCRzVDT3VZOxB3ORJNidv
iPu5FutkGG0untFpjMCUyB+5KuQwRKg7/W1t5PPCGt/EwJ1j3CBylEkGhVpd6IpgHenS8MabiRPE
dsdKdyQWV7D6lyYVH76R8izU0/wAyomYk8/NK3CzxElYBjmBmEleWpgDkHDFWVj/UT5riY7oLMBN
LwSq9rKaS6CGASregXALKjT75rlIGvMmwL0jeb6f7ZUqV7xs/YPv9+QzUfkWZQHqnMEevtUXQqOT
JBqbPM+1mI3Jd8BzVHtcnI3WHzzDGzjAsD57ttIORl9tvycRmlN7olEiuBCZixfnuwqiB4Z126Lf
mxEjqlIIqy/sPLEQyue7/eL1OAtK1eqtvDydmWADGR25enSUHfvsO0zHqwdarY7DRkfovK34Mft3
oTHVscD5GV8QumJqccbycs3Zca4N66AKGPXIM3lyJuHZNCS3HrbGhOdkhP9QtsAum8n0cIZLqius
IyeUPV95eZzvVU1qrOjOLtfDeg4vq6fSEnEuIcTIue4GsOAqhqpPdqCdSQZOYvpW/bdETa7hzO+a
HhXTGxqDoV2e3TmcafO8+DZG6kADppI8sesy/8NFC0X0RQdrLGmPeNlUjNpmZ8y8/rvDO//Y8x4Y
acsTcGSQEAZMX3vUckTJbkE8WDRFPYdFygJWB7lsHEeSQU/DgaWVw/MzQdvjd+2Fh2dwL44dEvAL
H6mAgkKOu0ODjrRSCrZY8Vrs4Dlypux/TF7rJHer0sCtd0XDmxjeTqWCBYI6YUB6pVHdrMN1LsOQ
yDUUawp9XXE0ECcDQm+wKVf3VTVLoooHtApEKx0MDbany/++pa+4BGO8KIoM3UdQ4oCQ5C11D/Jy
C4gdvZgcVYQUdkOlddjQyRp8cuC9j4ezt+aIsvfcEO+FZxopRNMgyBQ0bJ0yLmDQQ7OAXigRBgLe
e6Kw2+zCqFYvVZ/YHeMphaK+BhzBld+VWzTpKPiIQ4mGE3wiE4QOLo8Tj6WtJpGhX/QjZNGvjeSm
gXBljHl4xnqDsPPC/nXPvg+t8Y+nyCPjMZ1dx6MZNRIjZoKgDGNwQYrZto74Wubagd5w/G54hVC8
VcZPMlzVqmy10HOOB97pFdqEPWTOjzTUcnY4JxHhNlgmCws4vJHykERRyRhZI7dBCA+dtaZglSSL
1KovmRlGp+CyXO2wq8VCP8D/LNEBq/99Jve9E0Gkf4BSZQAIJKVzeeAyGCNx7izYHHM15q5lu6/B
BMwUbUU0+09cVPwrxr+6Qm5A4FF2WiXR5AJpPdX/UhGvfSOIq73ooHBUVZD9CzH5Wca610oxUiE+
1hS99EQ0YFFdh8NmZdWM2S7feqbGRL86Nub8/2YPaqjzLP2MMitB/rEFg/MYN8oA6h1btHWtMrs4
qNeDcmZ8vCjUTK+Z0KohV3QJLhlbT2Sa65uIT2CWNv6gdysFxG3vWxrNOpyMRsr0wu6UvrgnthTJ
1G0ezIEbosJ40M59W0bW+wSHyNteEQo1ODscx12GLPpsBX2xW6ORWo7ZDU/K/6pqU7SRXl/t2hsZ
0cFFJWk9Rt0uoQ05ao7jmdJKf4pv7QXmxdM60DocN31yq4Hn/e/uHFyMyiyeZ830CFEpCx5QqNlG
IcVPB++QvQn5uN5+HNbfIslebjlXjvWhC/7uu7HFR0WUh3w0jJKl2ZVisZdQgnKJ8sHCqdfopF5J
xtqwF+5PUDYrxUDOT/Up2SFX7OjqrqXWAshJQ5cG1ORqfaIyn6sEnJgqQifDZ+qP/tf/8cgKx4mI
Epo2j+Pz1ra5ARhBDh/GcoidUGGNFTprPqLNiS9KdoUuzSaHOT4SbpfAIiV4NMVtx8MHsphrVcvn
KngdLsL08ZOoyrCtKh+/sytLuB7VwiMN2WaJ5kgGMAa367k8O9X12bsdzYpU8FoT4q/EXgKuqTeP
TbM070yG0j6WjDxei7IRDaRX15YbFpAvSFjNihOqKaxrPRgl78Dzg2UliqcP06+xIdtql4HzDffK
ZVCams7D0ByMDFoY/444IfPw8YwnW/siVN8DWiXs2raYwYQok8ce03CG5nzrVJOEKHmkjoqdQ0xf
YQfD5OQ2Iephn0rSw9kx6nbUqJ7VQLHJ+X0OK3Pg3s5b4gMt7GiJfwbNTmOVgmcS89u6hzEowD2b
mVIjlOueZJxvLYeQDqGN2jpRB9X3+wfNAcGRDiq9LByw67n9eoRPnDCqyy+6gVbrpUk6DORWEPEX
FngJP1ZCPr8y9Vm/EgVJEv3yhp0UY72D7h4c9wkSIkaECYkTJnhUuyc5m79Y1LM9cSp+OsW8uZZE
4LwuWW1hAe4sHF7b4aKwxcMs3lxvLkAtB8yoEr7de2Smnw6Lc4UHmeExUp8Nf4HhzTGE7cF0KSRV
oAai2RaqomCyzPJz8S2IGgA+6Vt9cn8ef+P/z8m0bVy/jREHLIlZi4ZewI8vcgHSQqTdskP5Ugsy
4ivlxQsVScqxLWooEPfcnnAdV7eJ23eXV2P+e8Gq6K4ovDrwyyzDNCluK9wCoa61yVNIClRPMbZ2
PnSgtmAETKOJQW9p4Tt/1K4H6TuE/8DBlfyaYFtcyliFUdt9Q0kACUrj3SREwDRTtCtfTU43o9FL
fT3ERkvuZOz8ZGPjCx4PPzwBphFBQmA+12kNvZCOGh9RleWEtYYdCJRG7/DGVAPoZ1rHkHmln0WW
FfVOCJnBvS1stivJo9qG+2FHgaUwMQKRF6swudUF95K6o+twaukwZLC/c/qL1GMXcidAfSAvrtgL
mLX3en5ZhPnQfmtIQUZpQzygnMbCmTnULBTvWWsTV0Ik3rT8EmcEeyfoexLjBfMgys/90GkcRRT8
JMAD3jjdzaT/TBeLu+VrxPVHMiqsJHpkJHG9tBK33XUmsjw7HHp2ERtpWINkdD9SB6dSvtj1wVm6
+2TFaGpFEBspD3g3AfYMlDuyXU0nXpfRKTb+JXNhyjLfYrkWlHa9XSqs+SfnuUvok938ATAvOVt2
H7CSsSe+plGDcKRQj03w3Y9+rJlfjuTZCL3RUe0Vj6QKk/7zLwWOWYG+BPzLfJpvbUWFg5Sbmfz8
eaSp7HVxGLY2Ih5tn+KXrGPqdPYOH0UItUMGHvtwgu3TmOE78Ms5WOvyNoZxcSnPzHn+984kLGFm
/UJcQ6tg5q31A/7FmVD2EFgtwk64VjbcYo6aainJJMLkm7xSCybjwlNNCpLd2AvxTh7tWQzwGWWl
yf8IXnGn5pBMKIg612bexf+tVgAbrChnyEo7jypOiyDR+gNFR0jBxlJ7xSleOKu02/c/dQrXD7ht
xPD+nLXHloSmpEWHJuAGqTMb8GayRPP9x+/Pf6v7hC+AMXo7msVKHTyUP+agQ6PfGm+xB6ITgNL3
ymwowVlS3uEZ5n2ka6ThzaJC7BFYdVLZjPfX7K1VwZEeptaegJlY5cb2gIo+dQHghwWaRWPteIvQ
DaP0tvUYAQoCqnCAV1M10Yng4XbBap+T6rqcEuF/miOXgcCtl3ocbS2q/NnbbZFfJAVtAYh16Z/f
TT57N9wI7l6L48MDqx248qU78QwTvJU0INsOhxnTASIdfgkaKLJ/sKCm3cHS2rFN+5far+Ay9IL6
8rnkgDcItngZzm60lXwYSd6Tr2bpxFlBoM1FauW5TV8Jut/ZqOaNMz+HNw5H42GZhwz4FCFa8eTz
Cq1kO+8DGgF2rHKDBBy4GOS4uyoHBua++n+34b6kV6i9x+iniNjEuRL7w/ylT37xmFerKV+hF0Sk
b+hI7DjzcX0s5UKXkfNtHGEtGO8nlurga6WDRcj/iZ7Brd81peWMwJyu4rDEOg8mp7voa+2g8+3p
tuDdXq0VP95RSwomLYZ8afOTFGgyTOv/UJKPIIIeLYlqkzOf7xpzrqHYcRL67mcgVPoqDXHkZAv4
gkseQvBUtbsbsQ4bCC7MA1EoPD4U8ae9QDdbL1xF4+IlmmBKuFketmMKENIKyblA+x0SIEo7krq4
tBmOwnhAZ5PmfpJX+BLFSVyrsMCNDqAcHY+o27HOCILnnwolMAW+mtwe5B6n/WDge1by/MK7Ip3f
lHuhQqrwv4/5zs/gQ9IhS7lMj+M4XusZfZY8IxgbpE72lAl4rb53BJJg3MWuikGzTpWeANTUdCWn
3aXQWZLywXcRjeGZZ8gLVnw6q8RoYsBwk3/Q2329dTNxwKaYSZFAPtjTSQ7GmSzkHQBZCN0CB6nv
5WEuOv8zEmr0yatXw/DuXx1Ie3tQxmeo4jzmWD1mv3aQaunXi5UnetKSiQFI9YcBc+NzOQFWj7Vn
Npg5wD/TIrbWqfp3VvQXihgXhzkxsB5duh0o775V1tGGxQgCWy2Uo8nr5muKBrkC1RXyhjRyHoLy
6Q1wz6doB2L5t8jZMxgA+5YtpJ+n5CAEKpVxyk7NrR1RQzcZIuHNng75tGI+H8lzQiSIGhs6P0Su
6U3juzu17B7uUTMAy3mQYPOUcU8Z29xV79F1K+rFxA5j07q6kG0+VGBm25G36rOghcVh5UUFCRmz
sviB0EHE+OhhU0p7KZCjq6pmHRFn9YQisFo3APwF3W+XEgrC+A7j4b3e8O2rCaJVmyra6kXZDNWT
DHNqDuzKbO3nhVfybxXI2j2006Zp7YZqZkgCubmmVKypiMpzH+8PPR0BABFk+AAYrVl8CVNdp/2J
GHA9MPqq7oLapSM+KCc+RdxAUUwJsZB98HW+rWLEd6V1tZpU7rOGfjsqyaojDNXK6XlLft2/7KLU
1O5Z7yoN5IMS77KAEfHn6YwKDHEJg60g1nTRjQ+xPFVI4uDffLlMdSDcO4a4n7gyjZYoVAtiBSU9
VSSqhARAp/tlAEzU4Y0RfnWuu5qP6xuwNrkg+yumBUHvueUnHnMRbJI8Trb2d1xtyAxJBKV4qhbQ
Fy0nOaYxD005Z20VSt3SItZQ4RDYhltBLgvgeSPDGEMI0Xr+Gng5B2jYoo1eP04iNLp6OoNJp82N
26w9F7JbOnz0A7ieKJkP+/mxK78u39EqNaoD1jB2AuHLq7aMp/5Leu9GMfF2wKfjB0V+LsTZU3m3
jG8QZcQBmmAVt6GFQo2bCw3EVvy6BMomnuWH6ojK5H8oLfkU6PRwOBETh1b503OITbdbqHvhRp0o
vC65S2ymjH+SIJ5Py3oE3xKjE1FdJobExiSd1BPAYvTZtoAJoB5e4DFHkvR/FIhpbbD0kWjwwS3w
CAUcXkrj2fJ8pzxi6M+E5kU+Y6n4oCOSov2wW28G1jeS8vb8SjDssnbKAVj+WLm6OSzA05ey0a4R
1xx4UOdH/TEyHOVyM8epdHzZVxxp6AMdGet6hS+Jwvow7rmfQdg5yzAQeW3+fO/angSkJ9k9fNvX
gda71noLiDYxKceSywLDDWTmGOYmkw7XirqKNQsQJPjfNTZrQjxPO0Yqc3LsGhDwO14P3sv/kbKn
oMUwlNKoSKeMQgvomGEdMb4h8bpLVlvgRV0CGPPwT5JWvlXoRPTTtvfbSYpVzfTOYsvCDRLmiTq7
Dl1pWO0p1sGixGdwGun4ffG+zBdhmYIierzY1fx6WkJ3rvAsEu36cOiQ5BehI0N+sML9FGngOA8R
Yl2vlGmd6WMyUiKCIyvd9sG1XUAWA2dr09Anz3YhAlVr32DUGyytCLpvWKoHlZwjTLdhjznoT4Zc
L+CKSqEvNQF21cAXfVn7QI2CryidC9/W3mu08MLgKXlkyYM4ZtHYITcYuKRQ9fut2DK014ZHIj7z
T56uk92TuV5UHhq4FTW9HlJX38YvHh5xbIECnXlBqPUw0FGQllSdMjK8/Do9Yg2IY3B00oAzhuXF
yIO8yTacnrx6DVCj5suqh+4clC6HPgWE4oVmcoxlU8gHVV0irg/J2VkO1bp7refAx3ft12u5ECWK
Sm0oPbTmfH9ySCCm3VWCbrgcOj0z1sX0ITv9jjbqpYyThRUD+afyAePLeoUVaQjtMsixkvJeBfAJ
gQNenHXZGx04Adzvw4qn7zKkb8SS7Pl1kwZI6UzykY/kP0t82CWvtyWVNpkabobVsEGUousYvK/Q
xGXxJFvHvP1ECPIW7TQNbqoXnAKD6RjlbF/7qmbN3R5gTj2PZp6yBZcTWjBBkT9aQ4JqiftCtdW2
Ka3w4jjjN147s0hYmUiE9w/55NCAFJb2vcTW3vCX3dkPThZwRLpFj2n9APAeIDr/b6IVsQ9tUXWH
L5JVoMId8QWqad8NTZHIdDkw9mqcnkvcFJPIyhhKHjhPdnuefk4qT91B/5v5CIr94EKMecLobZpA
GduQSVoe3rFWHi3P/IDKkgJHKb5mJaIwgYvXXsG3fNhWhrHqaWXxazhEh/aT20G+3YgupP2Rt+IC
pCecX2xO6k5mSxUF9tMhiBq3+Dg4WlJIEQjpSpsivem3o6NGwWD0BpT9Me0lNSoPPIQlZ4QaO2hm
DVdXnOGIW080YAKRBi8NPpL0ShnrSplXmPGEufigyJQiG4U/8EedhA2YKo3ERutv8XIWoUiSMrzC
OhZnLJx/SSNMbpzWgZlWNAlBbUixDEzetIzVA8lrLF7rgkv7CRfpkRkKVlnwGGORYpstE1apVHD4
Br24lvo/esFUhcBcpQsB7pnTUltu7uzJigLGGS24JI11AzYDR5kiSCLuRnpwshmCk9pg32D6Mq4/
19A0YLeUrYe/DpiR/qomBAuq7qTSNarF6INOtVFVtoOqzP6MV4ra1UOVqUJVAed/vL40XmZfKME5
g/NzL9kzPVRDpIJ1ii1gxplCcf5Js/mHgr6dkMlPCK09EYqVwUZiF85yBk77EeDmd+fG4WmA7jpM
MNZXihanhSZihcCxaLOqnFQ8jlC4qqA+U5A7RlBk/huxH26/j8Hmvnt4MEhaV0L0yJYefZXFLhFz
mlfDP/gyrc1qfTBS6wK0XaFfYz9FBT1N3bUOYLHBR8AdGjl5J+iEAOwda6G5xXph6QoPhGSoAXIu
qpxrXJi723Fcrgm09epNG7P7zKUUKoLpxViu1RApiHL7Tu9BbbmVh/iArOSAT2uF2mrYyfaPq2GI
XwsxLdrLZe/hfTjhiJ26PoicPjM5Y2BYnqW6z91ONHrScshQgpR8yWxsAKWtIVEwaAbwy5P1Bpdc
V9eR71s2Q/LvIeluLPKVfE9nuiGOG63qOY2voTTFHcxB3rOCO0YAA8SW1PkcAkTb1YzG05DPunwy
HLCodSGymj6RAkHAuo+bgFHKPI+e+wlKUfEApl9CC3z51wWclU+YGh3ruvqaTGocccSYx30JW8JM
H00nxdtOMr1eGhmIWtgZBSgEgH/qkQOQTjyeL0BEZqHJTRjSXkgWwGO/GRJaG3Rwv4B4lYwWg3Qe
GgxL4HKfY/6KezK3oggnxen71csnN9BBKYLdFR3FBXXnFHlgJsihkoLSjsVEt2Ts+RaPbfYcEF71
RepjCzqjfUoAEYiceiXxY2VKCYn+QMls8EyLyderRB9HkDMOmbfSJhTm6XMLac4MlinvJR6zel3J
bRzvRZbrRS2hcWlw5l3cZkn9bKJx10wh3We9gQCa36TfphxuibEkxtE3QatUzGW7NtnnfPe0qEnx
fYISovJ98lpXjEaJ1YRbxPkWREd3ngn4mfqib/kDFu3jS+mchJx9GLh+9AkvwSYmndqYGqSRER0t
rFlZmzm8e8qcNDyvMeRHlmPuXHnC7dxoJ7fRJtuxtJd7+duek/bERYiAfp1LJ0zsFx/PNyo4KVdd
jBQwit9qo2Egjj2QtnoDyHDycCfzzIHqef0TK1ReCUzl7J+qONB4+dO03ddfQYtyaopguPQpEAKI
X+ATNNuOHqM8UhFG+gmutcA/xd7gubSUoCmiIGTpe90N8lgwaIEqQ6lQULPKlNz6dd8qj6e+jnCw
0ob/g4sEBx83etruSgfG60hX5qkNRsCNoCVyTcnNfgRZJ02xhJ8dU9LRAfqC1ct9UcKEyrNOGiEZ
twwD8r81eL3A+uRYj4/WITDn26T1KIPu+3Q/C3vUAw4flU/8j7VC0qnRp5ZO/Gvw0EkQrulSeuPh
n+/GRaM8+s+6Se+rrVJmx4yXit56nzE2Oz8OqKLe0eIMOgBLarpL3b5b9CrU27GThRKmaH11k2C1
eninmYuEBAetNNxYk2SBRCnL4uWgrvobzuIJRqqJHZPQBVpvxmQp7xMI9qN43GP/u4TZz+ke0zah
+FuhLYIzljr8a6c7rR5wtlqs3VRg97ZljD9o7EwW7qEhL7zCJ7Q3ooii58Q729R33H3Q1l5Ght9K
Co+C2wz1lGVoAcSL7eYWNdfXJUXECJLwbsKOZWnC1OoTZcjR0Gu8AV0ftrk7GQ/IzvW4KX/fQTGB
gbYU7WVDAEGuCGBB6+qmK/ssrXC0tb1JWZAqcDqJA7g/UsiGuSXWfK3J6/+SkzpGffarKxLwSgSw
bzcNHaGyS4RIDcc3yGQyqhBYPKYj86XXlAM9Oi7lEkYOeKMuJvU/QOENUqKDf28Wrau7p9vaMT41
dmC2T4a3nmYYjc3NA0JCIDgdF8tmwgnU11TZ0LZAMXnm/vEBdm3CMy9Rg2VzNsqhJjNC1dX6MYz8
eiN75UWKDCvIl7fkGbR02h6v3+Y0O7Snta383edsWKzjbizAM2M8+j4gt+VXGtP30QcLpADcKIH2
1oHRV51TWEFF7XSHvoNKj17dAgKxWA02/624srvhj0SesGO1CcqRJLGC3PAoJv/M6EEv64XUjsic
aOAQOFL2Q+FfE2X6NkVhrTlqbU4eXakODhqJj6ESLctenIiVxIUlo9YxPXhTs0T/FwTRBy6WuKwZ
OIOYrORCdI95Oklm8kkcZdCUUAal8pm+r4srHRKt6SHz8Ryuk8UwF5xgFtJJetcQcKZl2lSlVELJ
t2VPb1PC7fro6XHD9WjWEln+FfYPfAXVtG5wQiuT7gsTvlbCqML8jT27nHME5Q6xdzZYGuZzMTJ3
aSPlt6EaMab3dt0vOP/VNL04cFXXemu2wjXsmTuw7yIHI7jbrAKIqT0VRTs/fnanrI/eSKT1EAjm
aFFjQgEJqqhH/Bx6Ya5YeTaU5bpbwrGSsJq4jkNb8Md6A5uV25CzR5U3axOydozhwhiAEq2vXS7R
7lHu7/Go6Fb2yn7t08XUNfap4u6a0L/iLP7t2J8ooQmW9ACav5cZpoO9JCTecvvl86ggjwk3Wrii
V+joMDm7KmROz1hyhOVN7mH5tZX6WP2F5LP7tdwQulBPoWe+o9p6QJSWEBB8j1EO9bt9tUY3X62w
qWZD9deIIUY0BWLJuPdBmlyk6A2RFipuCE9+fdBsv7JQjqbWzh5FSsEvxYqJBfso5OTpRbjLtaMg
oKsMk5VsAjvgbHhobtgrerYtnz418wDpDXgnnZPS2DG+KzqRi4sau8t5msr8Dign4y3IaTyCRfA9
lG6FIFJAGF3qLFOz5j+fZOD6Vhy/BPfy0x/6juOQpSCc/p8euDSAC9qfDEjfsYrhVv9Huwwi5CQ8
++p/oR5ChPpcfZyqYLfkTosFZKU35IzVdtlLyBvE4hLUws5rbYWkqSk/TWZeKKe6jj9FLADYn5I1
54r8HgPv9EY12C3D0QTVEYcwQLpW6iFHVFFVZyEh1MeYNa7sxHdsUuucMv2qRiMG4ArnNrLxClrD
ZtwAw2nXM7sYGxx2W1r78geTjLNjEQpZ+bb0aF8h5TeeWa0nNV1lBctl/V07zPRUNxuzlxEs1M0p
z6nCBHfIo0GH8sR5Y/RwVRipImkmX6rlsY3IF+uK1UHw0fZ71YOXoSs4JeTX9MHY1LEQyEzUgLZt
P9aSKAY/tOe4NUSJu8EwpVU3SSjEXojMMOUaspA8UPAB0U21IUAi58phv4azF/1OLX3SOupIqayu
jRErdCKcdumZHTRtLMQd0Amxs9uV3yFVl3WLelAxb8wy20yzQz5PJShSm4qHY+XMOuY5YOBXNZD1
SUl61EySY4+3PJFG0eskZvdOMh1Zq8I/ZyUZu6KN4wt55f7MhftPVMPM6urli3ddx9ItL032WGWq
/Mhro/q7pBqVLDBZwNC6z8cSkTR0eBzSu8JwIAc+s4gtYl9Ocfa4y6dUCSyRLOsnBmUU3/n8/kWC
C2sQO6jPZhc1U3sZSRecUCjDixtaY/GL0xB6VeUB6+ZW/piMligXRWPgfZJpS62SQ+RHJ6hCYbWj
utPWyu1Jxky0yUwB3/r+iNnFEya0+52rnRh+SdDU/RZTZ89+LPa5Au8YoY/6K0B+z/1idXP1d1ao
xAiQVl0foF556IT6RIC2YPNIeJxH+OaBaWbKT0H0EerVs+5fsTfox/OaX5I31rguuNdGf9fx6F9k
QLUdYoNS8WnynmAzDyImKXp9419hLkm9DiqFic2jDpPIP7ly6edYGBJzosP5Ewd4Q3e2hq6ufn34
ctJHt46EBMjnMJ2Dj+QUkueY0xloIM8QN1rLwW/h26iDJ87Z93oZ0lyaypV15MuNbMrtClYGmtZr
uV40uAEdjA6Mma1IfCIoHaqapqCHX7LxjkImS2CGxY6/PQTnVcAu9K6QEtoQGV8jcOp+tZ/NDFCb
x2NZpmVwydgP03UYYzf1a02S7LbiibcYv+Dd4mr6uq9AnYW6AnxwLSYGXo+wueZwu8a0CTKcuJ+e
JO+ujkAk1IZ8Xbf+aD7TrumQypWJ0ZBTIPZjZPxRqfFL1mvmPVoACQccNQqFanVNB7Q5Jt0ymV2V
V/3nySjOyNkAhjiiNIS+k3g+EnhczQ4lrPOO62OQxVqCNZYqv63ExW1+4gIM7OLMQxX5rDJ1moAi
kpf4lIMi9nCmADvi0GoC91Lwc6oC5PSkjokmZ5Vl1dS/AyPeofEKIAsEChA80W5RJnuB3R1+RYzV
Bt6ZNuYpIwRZJZoMpbOissi284Ert5/jHP6LpIABqX1lnX4mGMFab7LBdq2m5uGntY49gqqGYYAZ
lCEAjP53AdKok5DGjciydtEC6x8cGNJlIsRfJf/i9eLN5/HyaQz86bqeLuqVPowUxyueNtqQ289r
JcQ2gtHszh/5QDVeNiBJD4pH6yPfiCsgypNsvz+Wa1zGwtIOK/j0vAaLRfL3ggEwbhJXvTCsQDIU
F4+vukI2XG7yotPqvYnk3eT804aapFcnAOKfGQuYmphsofsfOECTZIA2WF0rHnGbQc7nVoqqnAdO
O0yVyAtbMHUmXwQPglU00op9V+a2O0WesJrxz22CfGJosqU3Xh9pMeq4pCyJv16dk/d8PFtwtJXK
T9yjiQMqKWXJZPMCzkHhctelq4bSJj8ZUZ21IjnSN2d7BwW6hV6HIsZZZepdYXonIWp6ehS0sEki
cTvzilkZ1xfP0etYactDMbN4eJbVFJKJihhDC0GX4PYj0q5xEh0jnxCs/yssXx/qLU4+MiICIoOV
a6m1iiWLcOp3c1ENuuX8ihyolxo/ZVcCaAuqBUurufwfKNlptYRdWCSep+HsJI6H4x61u9R09pmx
EVfZ+eBYQC/PhhF5/lPsOaEff+pl6X3jDneBYdZFa++AlARFGeXQC6W+xIZBwlyrwlOQEUoj0sIE
VQUXGi3IFClXS+i8edz4NZgxJymaPtM629xRy+jMTgCWzuTe0Reb4946cZ4Pehxjj+e2j7cDlvCr
ilmd23viaS69hn4oWkWyZ84Rt6EmUBIr2XVKjV080J/A673Q1HeFUpgnbx6Ql0Y79Cx6yETEKcJE
LAK2JmNVgE3TuxMQ64CsSmJeGRUCkSXzTFdzcg2Jf+cAqoPyD7GFyaXVXxaeCT8nQUY+iulHnPz8
f0bE9gpIzAFkhRyr6HnE6QK1rr/EuI3ZrTCb2otDdWbCIE7AauNIGGxiV9eAIR8rXBk6I3sqm/Xa
ilKbGvTTOEwpPSG5OJctozCz63DgBYqchYP4R9mSy2T8H/TE8cCC36wiS6msymaqeViMvjGQdN6V
CITYnBa8bS/UqNnVjnisKDLKm9Bqb+0vH+44hu9Q08pqdjU6pfuQe+RkcU3hij6RdBRrTNdSvWHw
vTceYH6wRr91jVLkpPXvr9wyNs+m0EGaR9iKwKTTRbP6XOeV2fDLwgtNYQDaINl1UHKugo6LkdCF
fS668YEvuhrt8moG04mcqnLwMx117W8oqAm+lI16fIuQMLdpaCzDOJP6CBP8I4u0+jvXl/bZUAQU
iwnLrMSsFoVMmjIUvPxk1HAmR01w7cih8UyM+6g9Pux2tvFMD9ep97mP+4rf+HuVxx1lv/2Y+zUt
uPJ8ZBR+9h/RHnABDvpz5rlUQtkZBCabSXVccgzE2bD2nIzh+MKPyoabO6/LcOH/0GbLN0JX6bd2
lmIHrrskWSIEVTQ46zd6TiCNVqm+vP0SWmGaeF0tzQKzmdH3IXbfE4aGsAF8bkgVpXqzEbYOtLmA
gY24ZOmtjNQn3CXMCIDuH7nWWlhg4wk7yy4o4M0e4/5wYb//FasceU4WUvawvpENH8RqNk71v6p0
Fq7idrZSc7VJIYlDTpSM9PDd8rA29YFZeAjorJM8XWCRHDWKXOeUs5K8qqM6RvPoIUVjBaIBMCn7
QqZMDYh47maDKbcZv+A8fK+IDxwzzNP2jGZUN6ZaIZjV4jeXYmarhWIulwIPeT0NFYoOYUuABIYj
CPiFwy4yZAMO9B3GTgEIFQL2MzYWx43FCvTqC2BTVnHnCBnyIc7diskrUmKgawQzga2FozDKH42b
QiZxnmtBbYFrEQ5yorxdwDoEm+cXERHH0BPgxcCOjLdFLiLn+hnCfuT7Q50v1CHKKDLiv009mvS8
K98nEGZr3Si+dSvq/anD/Eusw/ay5cPRema9JwQCrempyHtWtIlPsUOcO3Ky+ZbxNNElZyaeEmws
648wwfBvd84Dm2nIMrXZ6IrNgn4R4uNmjfU0E9e2yLviKmUk/q5G49gY6/CpMP/TB+6X9a8DyC9g
+JkGVWouH7iezKO9kihTWbNwCwtkg1PqrcRzBl1qBOtRSofTpS99zwPAROCfiJrTRH+Eg30s7SnO
GZSIef3rSjsIQPaqWYpcJUDyqzCqc6JCrB7ACIHNp2V2OGdrZcMs+9oIkFIJ8MkPj4hP7yPBEvWS
gpKU7ueLaBvVkXkdQhOl2mhp35zdHLq4wfL/tDo9InN7r0OjiBPdS2lSV5voovuGqa/l3t+KUYsG
AYXEYvKaCZh1GVv3Y66B01zcN6CRp+8jZhHnvYOCR4DaRp8CxbUYQxXCZFimDnJvJDOU6o/egXm4
Qdcb+ytgmCh/Fn1LyNIdJOqmRIXJTllWaNGU9lgY9jWVIxnU3P4plFBsvwnb6u8m/9FXBtCkFefL
X2o/mxSN/E/Gv+Y/C7kFQHaPkXqfwo0IuMbl7zdHLj4B15wg8PQ33cQe6z4qp1QZzZsFnZxqrAe7
On4nk9Ewz07Zx4PA/kx2QGPUDj1Jj0kYLxTJFTQBegI5BqCnEtSw95B7ptsKLvKbS90396iwg/wV
wvJma0nAZ8gTu5p2ti4PqqktZlXWsWQbAZla3Yr+gkaPiw22oCY6Xuzc2pgw1Wt+y0ny7/pxzMmN
vTIoyArGpZwSJxde0aZzRnoKXAhYmudbnxaP4nX6JMKUxjo7btqUxwdgF+hF5PJaM3mS1IApgra8
xCXZKcP0BVyhM0cNxeOnX1v5oLFqzENlKuu3LC6z26s4rSQNl75BaCWGUMBE4pa4/urRVcK8RWLL
JYBHDcwKZMh67DhAscBk5yPAHnDoMAkyocEW0NdQsOsniyzA86XJXKLwJhHVfGPa9AnW3qL6m/Tc
wahiyyrtVl42v1AOC5/8f8+3c9qI0BVGxwyvY/0Iu5BuAUyUWfVEMJlEGs3i3MoJOrYdnTTPqreN
HgImxmLUyjWcwR5mDiHYd8YqIDXL1uKwV+wxPHV10vMD8tTRQIxUoh8KQKOiZ6c84uPJActlMBGo
6RSMobvMD0Q2N8iqUTJKYFYMhJTKdpS5HSvGEfI1GvFC9ASfjoDOmkEZtOR/kxpt5or4Fvus+jq/
qQ7P/1aPWP5We6IpaXKtawVbxcbdDHbuLIzO5WSftXuPrTj0iMVocuSgZ9terNyxLpj5SrWF8r6k
hEjJeieNbNwDPMhhmQ2Tlpkd3CaUkT0PJoYvkx1MWpJiiZuZDGSmMCVKHQ/WU/CjPC0DZxWdAkoM
ZAaFm1ySO2HK5NoUt1JBUERfgbmS4OamBho7vto6qAv24IC94oo0Hp5oOV7V2dlIvmZSRXfBProA
34QEJ7fCpjuLyhNQx/T8xQzNH+Z0wHTcjC6YM06obatYuwLxoujDYnyyCqs290YWWZkwXBNKYfQR
n3ENIr519xlK1ni1eeqLBX9yQLwnvppOUZL4F/GUnv+Cec4VZ9ylNUMAjbJqoR4WidHm4MhU3VdO
GlLQg9YNY76uRcTsX3ZHVPPl9kBhvk4njU9RdBHvpzMmooI3HngGqDM4LCx5Ho2CaCHcYn8xTz8l
W8vFsOs4L3VkuRIODQHg1aPkfsVZ+NOflx7vTL8zSAANinZK9eJqxYbBjtUz3TZAUM8FRb9/eB69
Kb+/WjeyNQYE5stGldySl4eBBJVVsodO4jUeTaJpXTbPXAqcdD7pwoZNvDGfFPQmjEOgBWgTCmUy
xUAxFS6+S46Sr6Dc2c9zd//TpaoKveILk3gzl8iyH6If+QZLgBjYW1H1QOb7nrGQ3oDpY1rN49cF
GpTArp8zAL0N4HIgBlrcmQUnkFiFRBewpHNvMV+j4xsLUw4yka0saogAroqultsEhioARLuJxw5/
1pAkRrcWAGkVVgsNRyCKhOlC9q5D6xkzy5EwGRPvtGgbMS0ojuV4kb7sAkmrTDL5DO4+w/onj4fw
epZ1viXavKQFYtjV6kyMP8gXcXrmfKCOwGkuj1LmxDUtsuFo3cqUkyZqsgTRnPV7AzKRoP8gsE3q
Zy2LWVeb2eDNUc7N0RaA+u4NDTdizwlHonPcfsL4bZGMfHphUq7nl5oEHJRL0jNJZ2QmHtZw5/Ze
6pNlXnzrGvoZhIwYIKgeFzS1G5F62OG07diz0h62E5ysssc3qRkhQHDEgPtUoe4iwWLPJESyw/+T
W4/45jE4xfY3SAmy0IXDDaa67Y5F5FsvpLe53E6iow4jEeITHPhAfzfrvIBA3+MVGUoOaN24PRJe
CQ0fy8/wUIK2Fr2MpmaMvhwLenuvUc6FdMCSdXu3ZYdIwLTFiWWR1pvt3bQjPvHytUS6Klr/9PKf
RK6WRSzCmV+lM8feyCfu3sNPPujKxFmMDlb4xtMRc9dKVdUc5Hrn1aaDNUVCWzycxMLAcZmBu8D8
zHLTbMSh4od4RT5F/JqBtoQXp37WDvB0VuKhf4A08wjlUPLsot6SSYrYo2MlDuAjNpLf7OJN3b9Z
wbDYMu0Mu8tMyPgCQytpT4/MFDa+Tkcmh75QpslL5PFIo4rN7rgPCBl1wAUbQqmuLw8Yu8YOiVAe
AcpNzVNN2/pa3hxjnu/V190wXrYN+KBGXdhehKE0LyM9bgA3P+rn46O3qgZnkKjE+C01Dzmu7JH/
voy79ceqAh4j1GnlldudLZlEUP1yzr7TqfIZhXvZ69jkbbMqZhUG7zTvavTyaZNKmXARi+LX2HZN
ELUReAYTxT7sL4FupTjSD9VlJ7moVVm9zKWmD+VzZvVxCNUYaMS9Hq7OcMVmezStvXhUzbNcUIJ3
r8rlauNZy56hE6CrdsIUDKb/n5+JklHRndmkSXbEzNFZNqk7cmvNYNbnuyWriyI/SOyD+Pnj7G/f
jGzi8z/qHZuIJyRvMurc63bbFXFjCK8jf7BEqZJWo4QkIZVBov4NzzZIG5N/3jD9bIpXg6yaV+hE
Q3VEUuU1MiskKpwrp5477ULmLhZMWAOrLZX3OU4FhnRfLgN2XWCfFYM5A4mqpJMlnrmGXYxetPe+
sf34WdQ8UEY8FfOVRHKz6wGMPs0XiorYA+KhsmusE43YLbreEhDQX90/Kknzxrw+wevfC8NbU3Aa
2FfoG5M1BYuv43BtaVG5jSiSVzXETKI3cqWDqAic41h3ib6mAL4X0J41RW4yGtfSvEnXUjJt/syl
900v0x1CZ6NBsHCnq5jQg70nRj0JOqOwhBXTQlFUsxIfVX7rO8J8HYER26/4Bci7H5JDhaWKy3XG
xeGoNrG3PjAqeVyy7iphbKEoODTeI23kMwVfaUcQ3wwf7OZgk0UpohGnsg+3kOS0vjTYZR+iFPQR
jMkFSZL6lXsZHEH1MpR7G49PFdAVllvC+Uupl87FjI1z5keUsh+NI57uCeSaZR0NJEJFfDNcr+su
7SOIAEjvm8lGMfYqonsR0YaqLEkxtUNlGYV+MO15uLD7WKrwzPf45lGaYtf8+z3/RorRWFeb1emv
ckspHjMJLbw6Xng3VMDZZXLNsOVFnM0KipA7s674lmuGCQLxRxZ5G7Lq9ba4v65jQtxUVbM5LdTH
zYyB0mjRLLpxQZXn5zUtuItOE/W+BZpf9J6W/MVfeHKdulUo3aVgdLmYC6lRgpWOTSbnQjvHw3oq
9GFBmQjaC9YWxeGSV9WKgb87VzeOEtDjCKYez9GXhqM4Ny0M77deCYJBbbcFKvwaTQUJSWsK8H6I
xUTR9BikNoob23UsL+XiyH4oMe3IBRcHETvIiaFJwyPRzRm6yY8z4PzX/nJnGpIND41yDgphZ0P1
kACzfWxbsT8f1hYuMv1xDkuQUxjb/Fvnah05g+8gvKPDMQTv8+GVnquanQfxA0a+dLBpbgX1W9pp
20xN+BN8IBqfpniMVT6nuDs/IQ7GuJ02M0ZD+cmgBsKVHuGoLV+y8mM23NIwfwI1dNGVecAxhk/s
KUCVUGQyX0feu6Z6jcngX+bKVXuJADmuHfouhh7+mEoGfdcnhiSXySyfGjSG6CKnSz08R/w6tT3Z
P4B9LNRBeP6hPmQPQh6Onm1D4AIvJKoJJL3iYM+sYvpU9p1rLJqReetYW/qeezpXLqI43mznguM1
gNbcZmWk3/C/DPpHKnKSEnCCCM0lAkUtWoTQMF3ZxBs7C4wwqAteLgVco/L05ASntGeXRL0JpzCZ
WlIVQ9SJnyK4Kc2EBRWXzXoGFaFjtczEu7cR3dmNfkmLV1ryvR11sue0q9XDAvT098uPF8sxl+sW
xwVp4gbgYFyZXpwMZQTwe2J8SHKcJaCgd0+DWWY5IJumMFp5nkcnamzFXPOMV9SdCsyheQBKlzxj
BL0kmai4fAGsg9jf59BTOy6bp2E7g9/d6wxCkOUP+Ffc5CKbgjUWhELMsqKCp9kNUzIONJy0gw9b
HJ3QQmpMZjilibZ+yQkDQBFhtnsBT7uc+JruV4Y8Tv5tICRnsf/qJy0mN0kyfx4XVyqJFGe2gzYi
c6Vi0mb8VyDzL3jzXqtfiQS4UN0PwMgzGma93lbCjF0q6R8EPqKmDBVZRqj7rNIZfk6Y0RtjAilM
6kkHoQWoSnNTriNE2mN19NS9+AWsfyyc6NTTUs0O63omWUvVbiIWGnzEymdyiB3RHr2IGeQYeLec
iJOAUFIstgrXeohQDTvKU6blIUhIEgIpcKqdMnsHDqQyJ0Td0cvLxPWGKz2jRsj1W0rZ/SnZ1prD
mtk5c4q4tTs320dLNrCJiAO/TQrat/QzRB6n3GSTsUKwjWDIhwfocV3mwUss02iZI578mXFgczck
0AE8MoCjgvEnoTix9lFgrN13a+Kkso/+ttrehdqadPyoEzYLE8d1CaY8US0+AzCIIuMxIU2d0Mr3
PQqzfeOIs+TH8Pm05HcELDCB3apXv6RKRqSpKQ3F0JUuIETanqa4mLuxyZXX5IGl5OeyxNBxePOL
kkJmLW+GPx5I4z+0gF77gYnxVpCnbEbA5AOjMu4AXJ9u0OKBSbMSL7o/M7rrFguvng1NLDBhX0N+
gcJLBGBTWdNba6wWb8a3+ZP5zdc/ovCGfVNekOC3uFRyg80EKinSSbtlEkeAIh8TVcLmUJIYoN8X
MGfkg47CPFgPlAJsSLJB886nkqzpriK1xuz66qEDXzRfRmPetdpournwYIlLofxufubuxLopdEUd
a0L4FSDNHRYNaSI3AXmZpug9DcE6lV6Fhs2GMixnX0Oa9soXnV98ABf1h9xOhz6mzZl2GhfW9MtH
iwGtbLFeyxQjoZG8BlNZTjcKujEwJJJubvkUkL5UizHVEcmgKinO26eRH9qHE31wJAcU79igAH4E
bQd8Q3D4F3Fzd9IOBZqr9qp24i+cXoyigyqebL5aFY+CoyROgeUzC2BuxR/mBUKizHw9DFOZYhCi
9q3b70pZlOTwSkaHBsTrL39fOwT2vTIqy8DerrmXAYrbhWc1Oa4rgt+nTnPlKugkPGeu0d0S5aS+
zwkstx74kFGiEpTGFTm6i8UFi2W8iRtu1P0ZUKRSmaM+ruUJ5ZkmFavG4ENk5bsRO2hTK9Hh1rnG
pboyz2arysMV1R+nXW1EVIquQ0wq9dfKnnSY+82I96HHzIepnzCLXn2K2uvQEZEU1x515HqEEsIn
fnGKmYQYcBsuLo16JiICktKw0xKIzqBCfpufmKsepkrHHwzQP+hi0AWdT/UD0Q4tupo8iCnZBvvB
aOl6FFCQAouUvDLrCPI/srX1+uwRSSkaplPtHEMCCti9hp6sn9LOkmeo9GujXsPDSogVcGLBtCE1
TsdQD4byUbHHNfRKQA/zFpINLzBwUB+urb0LvdC7nYvLSdExz/7R2XeMa6sWa6rLzKdK1/CWxLFp
wUl4IZv+lC/o4SCFu7derXTp7glWFRnOZo6X9WnM4HErTbxJMiL+Zq1K7Lc9+LENtXxGucmTE2hD
bYJvOf6dzheN4Y7qo2o1z/x0+Zi1AvG6WrEJWy0CyHM/L+A6iIHmMBAdNYPUcBFXNITTSxdPd9MT
00QlVpYw7/hq+FqoIsNwpXQgICDOUqJYjktoSyjOWOCdlofnOfYBAKCNU3bQdnLj+UsEp2mHkh/x
YnDKikd1IYKjipZKw+wPDmTu6z6EF80qGHPlByqm+iTcfmHOvKj952LoiBVa1vDNwQxMMMcoI9GF
ivSoHFMms0NwgfXYHSTHPzGNYlyArinlM8g672X/aHhEWWWn114RCilVv98QD8B7oRHi2wjC4BuA
hAYmqxD5DK+dyUaPcqtXPXzWm/NjOuk4/GEJYvtFOJAV/VpUy6RWpjJVkRd/lMtxbQuOPZPzauqb
YIHlMcZZfbKal9jAUaAiQzzkoGskoBraaisxzzRscnKVvhEalHGtxkR7l3IyPCmt5oo7/Tazi3xk
cmOk9xK9O2F65aFmWfNu5UxUMJEJbnRk8AAyAHw3LHi9JyaGUkd8K3wCpxSFd+pMx4/X/Su/mPN0
PIqcqu04UmYtyqCV9gWjm4IXCB87MVBl51/+Zwsb9NGlI8vBn+j5oEIuYKD1xewsXhFJE7yHVFhZ
nSigymDezAkzHE/gfvcFBOKAoLJLrflR2WZO9MYuhQWyJ3yezzxXoysF4XQFld0XqADhjj5PBjWr
MrsUFqJkbSRWcldYTwRo4Of2tiYa0++uuG8L2D+4NIUjkSJEvaYfjQJcniA5Khq3d1uOIGlc21Vy
gNRUMUV+c9O/Cfz79NJbtxa4a/rrfNTUWexPxEq5XFk8auCQcDPiYEW5ajd4Hv7nuc68PdrjKm1z
8mu5UlfmbjRrjYZij2e4gmeIb4k49NWeErVUma7Gxf/EumKA0RvzpTrw/Z1n/3+890IET9Vsq2MZ
Qoq0TuoZ7xh5r/dfRqjyzNyBr/MmxNM3J0wabmDwblmQZdD/Hgpcsf52cF8bySMSek/lsF6ITnYG
+f7BWsBGJX7htB3wjxR2+w35DVvnUr3E8dqGg1l3J4TJoqhFJ5eF9QLmXAwA+b63YfRow9rRZ9L6
lU9YcUKck2PBuTrol050fldOBzuRI1pYoZSMYx+jTx2Fb1ahrEV4A7kn3VyfEmjr+M2f37JaL+U+
Wa01+1mmNuxXLLAbVhmqkdRYjxM/9B9x5kJG1Hjf5HvIXik63ADtNGtOuJ6UnPEIprPXQhsiVrP4
+O8qMrzRjxChyiwGOostvWoAAViMbciSDDY5fP3WYqVumnDri1IA+yykmRlW6U8ufPLeT5fBdAiG
Q8+9QLpi2Njhrx/mKPq3qJSO3dXdnDwXHOnYbC3QTdEINvPBPvNyREnvA9wYOSKfUQemRKip/v1u
8/n4ITsJllHHythvhubQXzQblEyheS7AIao8Clk6JSgq2VWeO1ZvsGCAg0Q6mlHY5pZQ14kJH6Pp
cWvD9HBJxrKXsF10qroP+Y+EFYihq4x+7nFnowwOwvmcLGbCF9jQWGDJ2ulF08z7mMIRwIMUG5aW
mRf2M61/j5OQuz4nK6uDEqhbCtvELt6uzsQ7nEtdgiEPRExJYOT9YfbX8AlLMWTkXx8C1+iB8ET4
xNWUsRhgwXwMX0MnHZDkoSch54zNB+mFGexelMT0ELWxw5ErOVBOPJxNnu8uETPaql88ViE+Ng7e
yQhVgXKA2NkxU6C3Xx00tIF+jxF4gNkmVfrmvCPnPCI+hURCIaYoCvai9pHjFHDWCxseVnbPfoT2
szgztYnvNAY9Vfs9PREkO99mi8FY1La5Yt4USvy/wcKDI0rqEqeH5uul483LBKR/sHwcgO2B18Ps
ums0lgv7v6rBhUqL+jr6g0Srrgn/6Ez79iVEL8CW3cKPWErgHXwKQFAqBt/RrPJx5Pw0ZZrn3qbW
t0PqgX6zoZi4FPDT6uR8wJd8igj0VdKteZNqkEX9GK0iNx6+X32vjbQ81ingWzu947YQxHpuUa+L
v6JwPdrPtrQNPr00zd1JZ+uXRUt7/e/JFVWB7GQNK+2PG452ZrwHxoMFn/lqH3+uah904G9o+6q+
36x+t0+pU+WDRPjrq7pQKw3kbGXqCA7UO34b9TDBaeWvkpD4QGmBqH48dcrvHldtcHaVpZwkp2Yq
WXdy/Wcq6+hwftK0J19yvWe4fYusBva5NcEzxaXEy67Zu3W8WRncZj0OOazlZdR6EXR8/Q74L/lo
49PIBokJtZ//6DtRXiaTSJoluWzpLYYI/GwxR4SW+Z/JF93COnyfq6fdzGKRY/xYktYv6atDSJCS
LFReF7Y85H5bx0co4uCr90EfTZkJToc7xgyT1VqRnxZP3bIpDGXa6sqpH4ulijPXVqalL3FS2HKG
kEMdnNkQQjUisTTsDr7aDYPLLq0cy8u05sqmdWQsa2CPm284qgG+eLr0tt1d4y+tzG5ISkADSiJ5
wKokQoO74b2OzdixD6GhI5ed0kk3gU7gMk1FCn8OVwe0x2J7JObXsSBaWH0wXJiq7ypmhN3NLb8+
KmLnG/HpkXWJdxO3To/GJMk6tzfgDvfkuFcA6Ug7FQiKSzKQpQs76g2bq/hq4eOeCHa+i6xp3peZ
+vcI3mujjG3ub5ooqqSWGN5ohUUQjplkHkrrrmlyLA6KZnWdUDHnqpsexAjfwL4W4ijUX9Yg0hKR
iF+v7xPPWRBoizIq3yE+Wkh+sAKdnFVW3MCYZ6VyrYrPME9BXJEEMj02+ueDm2/en+WasJbNowmN
PxjjkJ0TjnNJ1ORsP9sbagRP7r/1BAz6omye/RkYc/tyZ2cSJ1ZYDXpFqV2K3VZLcPjRu2xMgX/W
0PfJuQ7bxedPGLGPGPbBdA9kiugQYuVUoSPWRsJlgQrFXnw9cQWtTwsJhagbAFjjS4xlePMEZNAb
eBdE6MmNbc0SJcz4Ki3TGaa9sjJrtfckuu6SY/Vie3ZXiqMjimj9TUnIMwlfD6xeUcv7wTg/7rbC
ST1BjLrAjaoZkb+HwT3LRD8KxbwbdpYvXS9wTlFy+Hv9RIyoi5tCzOGp0JvcR8IVfUmR4mt5kfo6
/Weisagns4Da7fPoKVRKgiBfdmbpeKyGixN60suOiywY+FZUGPv2KpoWLP++rBKA3qqLtEz714Y7
CTMCl3mVyCxxiriyvchsnkzube1FvczpDcZkxgist7EZr1UAvYubO+8FQAFBtfc3x6QIfXivAbEl
0+svwbZ8Z6LVMXON8nDfjO8RPF6fgNTdq17bX8c/fTmcZvGZLjNA3Srie8P9UdbLxDrIga5Y3Tvc
2s2EPJVzFr5np/TdzsXkEeEnO7WYr/gWyqDYXggaQVsrBFAf6hLSpZcLMbqs/oFqTEalKPtmo8nQ
Shpt9EsOQXCR2BECVSyi1XrrVvNt8qXueOOIZC9ULmy9p3T5l7EQBfjFgfr8oseDg/yAzG0d/1kR
upH7qPWhSqFWNq1o7kuAIowoSxaUUIlbGDop07LiHuI5/rqmFWTv+BHZj8PEOYoiHCSg8G7dYLK9
giiOyByVvROJEYqsIvEnFmDApj3fKjwgLlILB6h2yXfl7JBPtQZgILUWEBhe4L4LE4UUGjrsUmFU
++5k0MQ77EeTu2/W2ptNZuC+OB6JAv4P4yIdzEAaq3re8wpZCzYIvH5iU0ttXGEv0uVN+JjDlV9u
xn4+KP+SdQpBxu1jTyHL7qSSxQBu+sEDsyps+UOrn9K7y7GyLLMORkB8R3d4G56sbxjXmiEPgxxy
+vBrt/IzXK3sGkbfV2OCoNY9PAJeRRcYO6PGgaOv/MKSDdX4Zj7fm5WRueLz/yuTLC5IZJXXlZAq
Og5zuEUsgjR2N+y+uzwG+BS0AakryxULzLuN1RzJ0LmzsTiXqyQ9APWFbYvfmHHk5MkvXYJLU7Yo
AAGyg/Las3S2DGXsVgonDUGRcDGM0V6UwEQRPk+wquGfjIKn2Ry6p07LYQWzoAencaJxx7qSEPqV
QbhyO8D21ZC9xDK9ptpn7KReuYPsRWxSbxCc27mGPMQ1QlGyZpBOB+UTFOlw2gKVS0X5aURyO/9F
Sa7G+o2MSdtwvsjy3ZuKwCMAE4wjHdutariTwtn50VRzpdc20qzJcKCyYJ0OcirWMmSoiREYeIec
dJKYYJURVe9mGnSCstn21k0WT04YOcGj0ySaYTC+e8m+TKUwa6ELn+9m2vqpXEub+10Y44lqXETk
zyqlS68kIXebJZ0Dl8gUW/E5utVIGn+zOi3GZpIQO0NEPmihZp2etiGnh2Ku8P3odBmImhHIbFK7
qZeRTWIfetAE5w0qpapo91EhIYPtwH1aQWmhbhafq7eZtpGbLW9zh6EHoVRtJUzz0vXDP0gP9cdi
iDkKwEbH4WoaEwP6LO/2C4viUEwfPPB4SRsRoAoDjq13OdiyHRWwOdWZgfa3vpmLkYgBL6p8fuE0
BRxkki55AaO0U2rEx8J6G8cmTTU1EnPs60ZC4V2dgPmJm+WtK+2A73MCsls1T8R0++DzBoIWa6Da
wC5npTcQKzF829v5nlM02RFC2G4jgvEEFPMNU7uadnv7z2qtI8IiQvVkfPCuSFnb/ZP8hXyck3BK
MDIgUiYLh+jtm4E6fMbHLuJkz7IF6Z2XiAgejVZdZ34DcJ1nJdvwllEMdjSgA+SZgKOCfclgnx7M
/gkIUZHMkrsXcljpmfeUaH6mpr3OVW/juG/M+4y4+0K+JV/ERiG20bLDn/ikPGHkcnRMsau8xSlt
qQ1NS9bZ3hWhyrVE/KIahaK/dkdaVrGGK+eKZK/AZM9zhLtXW2V1w8vgwi1oDomvDztPFLwZ4r/J
84RV+ba2khGC3kJE+XUesT6SvP84RJvlILBuV/yR+1VNLUrZ+/9dxZnfC6BE/whhWWbUXenv3KPs
t1lW+d8IfqwiAZv+4kmk1tFHSwlpGSdzYfNPPN2LSXyePwXY+Ni/x3wlTVbLDUlaYDei7UaKt52o
4VgBPB0uT2YR61V6u5jBDY94lGnIO+Q000n6f1fRwI343wT83uSaAMXVXKCxxUqN+RuFKLONXyi2
wJ+V6VPyFGdoBQikGS9160c0M7JRtJqwjSJ67uErz8RgBr9A4CeuswDIutc12N7dLmq2dai0eutU
lbwXikU0RlkCm50w4His8bGEILnlUknH3JSONyEyFndbgp5R6bBYuLZEqJnW81ZJe4JL2qq0To9w
BuiJTtFKAViwRQspKaO/0H22R08ifIk/CC9mkRUbKZsmAGbdh2vWdON9Spt4cRs0kSG6tZ6Tfwyz
vrN4O2IYYqg+o2IjdDZemos0MkiAB4OtegPxFD26kkkikiTu9W3bigLwPo5wJHXa2dgM8/N8Mgv5
Y9GzzRWhGAygL5fvnF1gM4DuXe7bPLXKlyPTp1vX0xatawOFFV9KNHumn+VW8t1hGmnCtEMNXKe5
uNYdAorQjExqj3xdk+aaAIsZKPNTcX1iHqg3A3389iY2uYXTIFmtGhGaIXh3x/mncY4SThTcBXEr
S3/i/OUn1hRS7MGxrIQLtv/cFnLWVSuUVyp303S12slt8JV+OX4Kk28/J0anvpGAzZ6DwyuuKCG0
CQr4aTHlDh3VBoOvoVnIfXaWpGIbadkNO/TiCZDEWHbmqewRyIG7My1zbGMg1j6e5ZFuH2Oc7lWd
HSC4wHa05ZMdKuV26KMak3xGAeFvFxF23FyOOpGBtiK6CqtV+cCWM8UZty2XIPo7nZgAvbZc+J87
V9jnrwzwWlabRYznIj/3QuABhBqZSplUmBMMZVc5BR0PqELacMw3t5bEZCrF9VIchOv1iyurU/o7
CjWJ5XsEZgcSye0UeoYJHMHv/kfSV8540X6LPWf1tCNO0JsTjGcHbR6np+VEnxZCVqR/4SbEKVjZ
bNCe2l6pUJLBxFgCzdqcb5wnPIyGbBPu+fA+Tu374bS5Tij/Li2VbzepbZABg6Sq+xJssdpc46ml
ZLFXX+bNheNBvDvAChG10PumyAo3jdy8BU3DuQ9RCDG8MBC3GtRs5NIF4dKg1lwZrHN4zaR8kItF
0HSuqvet1vdVw+iLZufygDUqPneAdzXZZbmMlKAl/kaqnbfIEou6ngGdLOxhY3E1OBkgFjMkGnDz
gtu7Cy0NI/mO+pvl/+6p2E0LEFwJOjEKom3xe2BEvdvxJItl7Y/V07f3n6ZKXEEHGncouoVN6Zj2
9pMhpXhXfW2Vsi74OPrUUYn0G7iTst/ZJchjVXEjfe5pgbC9ZPLBKbDwjL+OJs5bxNRVs8UjJHDd
aelw2lcgo3VFKsIjijzbIota6YUlr6QJTKp/SW8VqZrRqc/WRYW8kGDwFdZEcCxKbhwv9PrGn5NA
t4+ehQhL7vmebZpf36KI/mpIRAl271UmdRQ2cU5wLsQ2UIbkb8LE+cZ8KOJ0s695w2ubTdHEhnXW
1Gq/XrLx2UtLK31Jg5QX6j4JMyRssreePNmURaEhX2GmodX8bqxgCGSnLhjtgDtyX/r6HEvzWhBS
FLENSFEJNTFr+5wVuUvfecVTFKXeSEkO77Lcz+Wvn6hp3Y0G7ZrYCMFvPHVuVpS0rD9vGpoXE7/j
hHUgsTuluZi4yYU1px2LK3Cly8D9kQGYbC8b/tccdglLSWp6SyESl3YPY+SW5bdd81CjWU2H1qNk
TB5CtFaFpqStHDkqOnsmDWi4V/pGQcVhw6h4njkyrzDD601n3B/bEl7h7oxDU1HiG1+daoLc0lhO
l7fElI6ol8diwf7s+ItAeVnDKosDO0qsMui2yR5FsX+17cY+Tz4ewhLOy7BOfnMY2H+za57crva+
qfEalXXyBNpep5uXaxz9OR5mGe3sCl8L/v2G4cxCCCZYMjlYRUSOM/971fP5PEglXQZUfhq64v7V
yPt35EeJDK9phe/Xv8xm71Szq8R7B9PGqrxoWEgUWGrCXl1INSdV9Qvjh+9c5EOYXCIZa+F0D2SK
sXvju+9W9WJaTJKs3qedOIP2t/QJunMS+TElumTXIhYqVNbEQeuH1uLk7oJe9/rt3VfnbHRvRYgD
szfNIQCffqjIufXthMxO9dWzmCYn3NrvoVmncgSqtx7budHAG8bXA+Kwe6WZ++RhbiuTxwgxKA+z
6oYSTF4UXo7Wgc+tl7hOvifsEyUTFp+lb0ZwtB6+VizUwefIUvqKrraA+WfEWhPLvWPiCDMqoSCM
7lkv0lBfcLxTY3LWejrmmKUzUMy/9kx8jMMNBhFssmeM4C3F13+y9bDD1rp6IrOhlitVT345DZ+/
Sw3hvjS/O4Td8nNE42Cj/rAdeDIHHao0iipGUAfMryPa0P92DAHKrWRCZXiXWXVi2KBN8ZeDJL3A
ujJM3niu9n4ihXdnIYciWIkQ/G/qa6byZAXtCSc+WY5bT6YQzBrlXrwAes0QcDxinlFfMNsAm4iX
QiaYgURWJgC5wtj9C4IDA94ouPqig7Z5p3qEjv9UdMIkKwMcVKDi4wIrddd/RZQC+6cXK+D6mPh9
4KV9Ji6klZ8QVBJ/tuWiy2pvxq0Zwod0XCFBfuLy3igg6lmxVnlvj9M2u8zUYjwjmFQ72yh9YlqE
0Ux5m4maRz8mxrkvinFMRVFG6qH4GLePIbv5BMHETqa62K4RtJmweMZVs0Ps0xoP7IdKNP5cow6c
1KPHyY+BLfSpaOhpW+OEkM1z22ktaRYa1NDTd+9jbPpYlMSg+y6Do7MOMUv2YVdhOqd9zb07XMGp
zOu8S2+uEiihMzwlB8bSgdMULn4Z808pu2Tg4eXXw3QvEG/JWleQsxmZqChvv7M02FV3jb2ihXl4
Leb2tOMe0V8c9QnXiuxxAzwstPiMy1LdureEyVoGWDTWkkItfpuOz1EKFv8nzmf+ZixYP2faGasR
9Ctr24JJoPLHE0nrXNA4HTwvnGWJcAK6pA1zfLxWlR/4gk3eDeMfK5ZCy+OetMqScV+mikS6ocGG
5A22YJf9PYKscC4aol9srRYC7oYc1Vul7jk9qFLI1GEoceRVZyo8qONPtcvGBWhoiILZmUYsq8Fm
pmktC34P/gTvzSimDKTRC0EmZlT4kQ/q094VSQcPphOucymajvk6oP0h0O0DzwuUQ6T8l4LdVjf3
hl4mlLTwiLAZy1Ss3X49EShA0B0KUhD7fSU1KGBTS9hVSazV2gHc5BsC9H5AhPMKsFN+weID0vBu
ZypoGPacP+/Qy7IbTe05cM5NtDLzRyovbTy3ghJNXfn75QAcNaVjTgq5iWoC9vlglDCz0xDOjy3I
AY+xj0D9Js/bSoifx2o52QW/ODAR6LvNYdfFWvZXt0XpsKFX6Qpso1oK5uKuDUeWJ06tId6PvA0C
exPzDnCyrOfhBv0VDXblN2hAKKny4B/C8NZa9pauHlabJrncPLFzgJloX+PPFUPvKenJAzwJJRVT
5ujclAYDpEm77rN78gbE7T/uvPu6YFybpzyM5UHNtct1tFOP63jK/3UT3pIjOVD2KZZfsd+YSdB6
Ah9xzNr5q+H3rF7LUVrxBUFpkPsyMepWUXeHHxjK32vXBk4gcXMSlH0eMlAsiOjX03ZWPnFZG3+c
J+98UTCGLL7am8pcxKckz7JIZ1urkQOwHh8BK8fnNwWmW2zrS2UVHqitQPsJt45AoHseJpDCGJOD
K6IYGVSig8aOBzxG1YeBhltFssE5SjnoYlYCeyS0SIQ2JcMBgQVwki0TvyzIMj1brZxJNwE5QmZU
YAnQ4VHMZhkiMLwfGHl40C/KHqcpvaEqg4Cwm7roF5a829xQym5KumQGCkj9pfURsnVJ4lnBMvq9
cOqNu14HX07+F5p9vHyKB/f+t9OwCJR8epOphi0sURkpqdKXgf4z7LdX/iaW+QwmzHjiJ/qtvBtN
SUF5VTQ1DnnuoRlfXeAtfQ4Sx4esXY+sgliXyEos7DjL3EU9mZWsSBTk0jcg4AhhZg01OPIXE7eJ
+Y33MEUTQ33eYu6/p0YHcBQ2ZBiyIiSSbNfKzA+i7XyCkR2+ZEttyPDCVRIwOTnZWKfzg6jWcd29
0yqnIgENfCFVElU9Mnq2n6sQIbck0KAVfVUH3uHA8nGh/AR6wQuRnp4OWjX6/XvQ8iyj/MqyrDSs
szkt6WXRjy1gPTLSel4/pv7GP8Q4PUCoQIQ1ZIHVkrCPWiDNKDRfSPihDxQpRhUm3zBiY+5hetXC
OdxWn+v+J6pTgBGGHy9pFaZSvyeF8l5Wy4/3M5OOfAbOIEIQkIhRJtdUa4SwnfPIu+43qDgjgSr1
42//tZLUHzxvbu3ftjePFkNelzCT5m17UON+BWNsdwf88vtYOwHzIz9mm+JgXHFjxUVErqLWfV6r
rGSqHsvExWkY/a32l2CaYFBdx2q1L2LIUFWAJwd4OTjigBkC+DYMJg+ehb6gPm8cKYitikt7WTDj
FP98/+JEcCEZVt8xydsd3RugRcgc99Zz91c8zYDgZ42m03Qht/I3FvMaNMbnUuuzW8uEoavG4vIh
muG7+9W7clVo8UAeAxlqgl+YZHlP+YZLFBp86lF6GsplrAixVnhYWpk5C8gy9xsyr/mU6K8x+jF8
3Nv2B7R8L5jqdHjVqzrwB8Dnucfb5osPDQtP95uYwq6w+KrMQcs3zpJUnKJYg5mXWGADwdI2VZS1
l+rt6+ypjiC27dseHwJE90JCPGrcp30uEu2ZH15WEW+LFkSoT3gaDWS2kmTauEpU9MyfYQGveeOi
3lR+lKyAtKdWvfIzCPllU1e3opxBnwwbbiqlr9BgP42oLzYh40B+XHlv/ccBPJU5HCNiFJypTEih
deyzPsmGuvJukclsMBZAM55HMJMWLtzuyZ0MxxUo27jufM28O/0JHTF7I0RwwFMuwBzX0FQBYQjK
IrXWR/OA3yavzXy6Bvm2oX26evyHGz3uXFkWcjVvuWjA4lAcy2MxxNEcjXVsQ15N/WC0coOiP7Z9
pAKG+U3Ra+DzVNl68zp+RaURxZ3oN4uRpoq4V5rqdiE62F2u17JGvs553iDrd++GDDXGvW7Q5j8Q
7Z1O9rtxsglJLGs5eOh+8WWCe6+nv9nqrzmyMt9gqLApCix2XX/Yo5mgc5a40t9mUPqi1O5deG9t
rEKpWr6tDiDtOMOO0fpA/dIyb4zpwLHtJFMaswR6oKgfYWgOsVbHBo+RQx4nSMOKVdCyE+iYcrWm
FkxUefqSqjGB7aCV2XYRNaxkqV5YQnUASycAHTEBhgitS7JJeUxKfS4/XOpNeLUkbrp4uGHmxKRM
Ysc8A6EO0XSZNTFM5b0QsxzMbvTjtdb9y7PjvMSQ9fzl4m3iqj1274HSf9WKKE28lMngPIbvnRx8
WJjWSSp6S6wU4Hco8En3UdFz5D7yB51oSnsCKAawfbc6MHbPYc4HAfFe+YUxXB4q10jE8MZsKmKS
tDAs/EHi9UucjPjD2lsaVK3Cs5/3Mj5rZgNNbAgYnoNZI5AV9maR9sUqIeEbMJAvg0MvtVw1ZqZl
458cSHrwmFMMGxprjITQcK3kLZBnDQVkk3z7E+Pl3oEaLaFcIopi8gzUMeBuXbGqG6UaYypjDlZS
t/93sMvPADG7Q0HRv/pOQ1bgXXYsFppO306M8mY9Z2/0QcL8PsdVnYCkAe8plevEB1J7amaGhxrJ
p608TjYz3G4Ez7G7IENRzCbbCUeO6ohCaJT8YSrQVSMRDLuWtbaHuXf+iKIjg4KKfRi8bxeYqpJ+
e0AJqiPgM/NGsGkDIfqtuuSBLa6QuI0n6lotvRIFbMa9CiZ8nz7m7zX/D3AaUAnH5TQBR4wrlX6a
hXhKSxRshcI6/c/G4/YNFsV4mTNmngDApGAuPOAobzPUTEbi0ia+PLHtovg20H/F3y5qD/+yF3us
Fpua0N/HiEWcc90v27x+QyE/+dgFzoBsRmlbRulT4d9ozt0jeW7yQyToKzW/t5fPNuNgDosFVdJA
6L6DSqhpfcpSYjsmFVchNkQuy590MwJk+4muVrEk8QDL4RozsIBYrYRiWHLz2dfrC9yIVFspl5a7
wgEg5Dc62EhjGNYwxjPucmhDLplvhbQ8QwyLdfLcFJzUpY6Dc8pksFbNtzdkXEqD4bVrsf8h3SA6
n0QwlQNpVGftxmsm41htsBbxpkCQhmu+6m0DEGOwMK1cd3i1o3/mo1l4RBcf/CZ0yDLY+8fPJEPH
GeIs4UCclRpspj5QQLOwiI0Q0BtPU0V4PrHhp8RM59BIIo6A6mKzUWbJ6oZsn+oHXVW12qT6tRT4
w9dQiOP5jDwK8uBPys4pkHmUx+SGkX0eS68z709rJB6wYMtkD5R4ITDzmnlaPSTS9M7Pdxp4y7cH
z6ITKo/6r7sq0ZY+Utypr/sJyJ7ckdVEmDzid9vQCRrj2qWTeIsi+tZcsGpYP5Gqjxu2EellJ4NJ
g47rtpJhfK1TR6q42GOgWBMZ3w9nE9IF/k+NuMjWCVlkwgjpQBodgbTR3lzKjtN4grwZL3343KEX
q8vumHjtqUF5njT/3pwl4GQMlJdaHA6LcVAP+jeGtPYwhrhJIusZ78/y6FvHxRPX7LVyORy1nKU2
jrMtFoLtPRXqMpzJW2/7+T628ICKRafd/A0SfQf9Y3m6Tow7qF/Eq3L+YFS/H9cWXA6TV0cnkQUa
cOSu9gk6KEpJAQcXyJJvPPTSwDfZ0OrkO7kJPyZCmwGi0wPrwx6Dz8/bu7DlvJQ1nTF5ih78H9SB
z/JMrV/OwF3CJ+Cpc1qT3L0VZJqULT0IdtgWA4e9ziERbvIbkaR+JnrZRfFTPXOJHZrbj0GpMTqh
/iaDHiuKM/vJGvYfrXLUz7zQpVV+zEILfdvFSqetS0deUR3wm+tOqj5wniEKa+Lme18ASurwXcEO
saqRv6BxDfSMV5YLmainsIYYB0d0xQSnJ/o+g5Y2Y/EdAWdTZXVfoS9riEnFFELKcbPmADGFZMIt
4UOtCjRV/OmjGv00rHFLsY+1CHi7FTcfXyjRzN/QIFvQcEt9C3hC5kUCXtcMPpR0eUR9V6pbnmmC
VY2qKhp489VnUesoCqa8aYDmZwttHo6+/LVbYoyqqvrQRSIZY/w5wX2gWVP/qKsUDoMVtP+OrEdj
KswcYiT9vlOE3YuIbdU6slsNKUJucXjJu/8rGZw38i8AGGWt5IhFYgsG9YVII+txhJHc/MQXU7mn
X1NDmm68AR2ljYa+NAdN4x0n21nSNKzo4vZcojPBmWv5Ii8ljP0/CAjWltFOTRcawyK9RXLR7RgG
Tn0x6mV7LA2S5RBV7J5305QYmIzR+HYXrukPvniD+Y/B3zpLVvbivuecAtuoRp0LawSuWTSyYRWy
GVbRaMJ5+SeumiH0q3laRok2lH2Y2UvhdkW7FTY4yq0L/R9K7EAUyvX/5GtRk28LGBMF7MU7g6Hc
5RflAZ+1CL1m9i3KDUjguGlGHefh/9m2mGx+OmPwVEQBXNyYhf4hEYq2ZBsUm5oSogTsF16iZtVX
xyBA/4eWbsmPUhFfXq0xY/3kKcpRM/VzRDUaVvZgKt4XG9U2G6qTnGsKI0f/JyW4EZGibR7cfMdo
I3AzwQ5S+9HcSaPzwcC1pqnQPFtufMUioHqv0bTRZl/Ta1xfhqO0i7GeKlOLw+jlVl+kp19iCKsp
aMUg6A4/2UnAs3kFv7ouFTv9yieXpXIDE9QBc7OJzayOfU/icftD7pSfyA/OS0YR6M/NVqCaS1A7
1Btzi2XvukJanRMKEebKchP1aNbpEi9WWxB/XBESYaKPEkRlmz0kTqk10K5c0vKTAih8wcJhwV4k
JsjNDFdBw8Yr4zUdDWMpolKMUEkusgQIQyf6IqhLeuJI7CXdt15cejRtoDNNw2XQSOFR/acZBXzG
05uWdU56poSy0kyQikfzVp+yIqXXClycD+4lCSAwpCoIcl5GDiG5iMmuc7mUygh6z5eLxUsNqOiu
OgnxZkm13HUt9m/sSBV7f1Dw6UbFhdwVGA9OWC1mRfq+WB7QGD7w4s4YPrZ+5kJBPfrLJBoNHjen
1GqhzX/bNjDpCUBSIF6j53t+jr47qYziSQf4v5BpfoJXbCGfo9kXdQxRybil6ej1SyDpDb5srzrO
LPrKryqzUX2vjZRuZYuO1GPd+aj5051U5K7m8tv/Z+0pRZChXPaXxrYClnnOo0UMIiAgH2mofyg1
CZ6tmvHU0fncKv/Hm/NTxCPvPLQPHk7F8y1h38O3tyu6N4L4OhofRDd9CGLZsOBL049AfQC519Uq
EVrICjuVedPzcuq7ks2ItAiqF/71E/DahF/buhmwLQ1ZfYnES4EI9ervjods0gB3xbi6vLHgXydo
er16ZKSCIyEdiyUhTmIBEURU97/gleO0YTzyCTQcU0Tbxiqey76yIDTTGRRJoo/AIZ+0rnX6W0gY
Q1FnxAT3ZfyPwoy3MJiD7yb25RNd5IHnWn9wh1U9kcfERQnfKU1Xov51JV1hZfvmeR3MZswrCGKD
INTPrg/I+bB1hmPbqYYRYD7YhQpfPB2wfUelBJwOKVto1/wf3/LpPmWw02Q5FcrkdEpD0psAxuFB
noWs5cBp6DxNjQu2TW+YdvGfT7uX7qZAeUPQQzP0+v78WD0z1uLOh9fs1ocxdGbfWNlJFmrksKxb
8qFyr/1JojBBt/OvlsearyDHockhVYaaRvs2kdlPsWeenY9C7O/xlrhPCtjGo8T2eJy7IILESkoy
RWlG3jQANxdE+8mk+TxvI/T4jWQ5ptVGRPp5Cb8W6EftsuULxI/sY1lr7bmOeUbfwD4Xh9iAJq+t
2j+a2x9Fint9R+m0jNkv1Z7aVgzVaiFlpQ3rLqJH1j+NOlx5plCwjQlp1pHPA0PqoFZasSty3ru3
Z0sGAc35En1myMo4TC4MlI9vlTRDxePRiWMucWOzsRtG5SzM+UdZkJElScrEprKREqtvfkfBWrcD
FrvsrFBX8gdYT2VGfUdzYq5zeq8pyqPJpd7/v27Zq8pW8dH80EqnR0ejLzdW378ZGA4OcgvQRmjB
bMB21yi455iuY/uJKTXC0rgqrS5ZueJecv+4GImcurXbieVAagiMUcE15OTGxKMuBlIHJENBLSpp
+fnZoinN9939DTxECHQKnv818INmUdURsQxrj/TsH9iDdkO2E6PWb7btGySwgwYBr5pS5speKukv
Cvu51wdC/Tm+tGqKqBOJIPkEt+slujilst/P87c+0PPg/FMIegGFSBsUhQ2QHka2HlJ4ccUg3kWO
GldMgi1vqIQdm0Gy0z4kasz61t764DpjZOtGzadJmGm8cqBDB9nqLLblGWjOXWcIVtbfeOMEhxYJ
UytH3HCiaOKNeF/ee59K7ejIRtzKaPiXuH+Fsrf1I+A5b0LMp1GKhoLz9H4H6RT2ymom4927mQWs
LjlbGEnAKxivgqSSkD0GyisKsdPUbNio1wvPmnRwHtECvLlPYeE7AwYng4muIQIC5LAhdUQQy7Aj
tiIjsHSOduxRDgWahA58L75ou/TLocVSDi+fJ9nik21A1gYT3odrK/p9gHb5O8CMcNOrydfhX7oJ
cEwadyCiNO6GG2Ob7RboBnJf3/ThpnCr+0f/lTOMAorpAC/Hbm3W4pVoUGwdT54wWkI4T+vO0qr4
4pbfsGY86xU+3NsD/vweq1+e3NTSaK2rn/Y2AKAvLqCrJFsGHUcXBXDuTzcMb6gS6H+1ZVyrTZfp
4lgiuAaw3O1mcXp/IR1uROhfmq/D9oDHqvMQerkNNo6Xi3go7UysE2z179RwdrtaGFpLmQO2aNmt
yqVLh5uKCw/xAFgS745ecddcdmmO6aT8SS2Aq53liDNea2yZWxDWdRzdg95O05Tc6WX9LC2REyYZ
VxKjUU4eNzyykYGg83M8+B1qmEBXPufu/1RW0gOHZKanSNo83JdFPjiKau+KW98khZFGnNUgb3UJ
11738ISkbEkBvIwBM32xLRfZ/sGFfg8iXtiC9puKBkyPUO1uYM/F1RGDVkq9PMqMye67NQmUl8WG
0BqLudS4gOYaEp6zYk6yAWAtLuHQ8aOsE1Qpd2lw+Kqf4fDWQpgfa99rtF4i8J59dq85SnI8Hrvw
6O6bbxG1SFgwx5muFosFzLuua72ypiMJC67J05uDGA7ZhFOnIxWmlSWi9zWXO3ZFQB5C6k0GuKlp
F2TJPwBLpDtubUO8/ZRcFbA414qdgxr4ZQl66B4GcafHB/oElcNxDHjzU6u1P1VVfc4ynaYKKGeX
cD3PB7uqhcDVD4vJHo6zh3lJDfz44wcoI1JCIk1MorehMKkqYlSVOOejcUxS/8ZHlGJNUw4FL6kW
T2Aw/rYA4GXmoOQgUg1sMwT4XtYp94c/eY69jqiBho6loIBMyGA3i0rRnQ7ZqC62OJx1fB03NB87
sQUgi0SriVj1Q1SOqnxZb1aJwKOtNXqixbTNYl9oaf2Hb6NIW8J3EEjuSQNVlLKFpGhvWvAODcmd
2yuIZnfh+gkJNGelmkBtsietBNGgedOv4iIS9t9JMrpzlDPzjlwdTS93kNPvI+m0EHqLqEqeyb9T
0VNvEpZ1TzRXg3jnHLPxlzQUNzQkVvX9G0gy5LHVjRm0IvHXGwEF3rqcrmgeZ5UGO3SHfOkOswXd
CE00R+Xka3HOzfxoPI9HB9hhYK9WyH7RYrYN3njXj/tmJGKQZp6VPnhSYDvYJH5T52peKRmBULCm
G55gCB04lEnSL3+ZGauJXy4S96QA5pFfoYxZhaaiLpKstCx9wBq94AcrnRUTQSz0++Gq7FVYnFku
7PeJqo6qUhZgy6LzYI74MbBlmTgP5p1K8ZKBsVXxYPwDphJTiIWvdRtKoqP5Hy5C+zIlxgxzyPQK
0rUB8CYb8bxs7EizT2+L/I8Cz/6RYhswEQlWwgeVuPF21HZuaediXofwq2MaF3qe3kAf8w+1WYTX
wviBxXJOz2DRi+dcn5v/ayCkfIRUNKCohHndNKx8ow8b5j+NcF+EjQUUb2OORDIAIZOu9ig98ION
Hal+slrxn2RXsEmiKP6vjqqxz8BOip2hoOakZWTkE2NUxW8pDYLN/7LEnDZJbJKs1wK4837ALTak
wBZhjYZ+H2Z/azyBgx1ma1m3ymqNvKW60EsHoiinNR3xhVT2OpBMRjNFpBqXrlNIzZVY8tC7MDCj
K2bXJ93OEZn3VOzCxJC2mDujuXnbeZKiJov1/COiQcXXTTQxC9fYSf0Fnb5wkY3OKPKqnGrQfM++
e+lQcwFI7yPhstCN9g7oGzIkqL8CDCxjSc3nAZ74cg81k/XsM8pNIS9LAZPZdmKezNfNZNrC+iRO
xXobI8c93jKkDzaryru+xmoYwblAJiPfYDdUBLtV+MprBE8m3EpfNRcwoz+idHWxqXGZmL/LPw1J
4gv+zQqO1kVp39XWPdRno37OLz0cQOex/YqJ90U4pIoN6jIPln9x1YCadok/V9QUVerkv8Yx6SQS
ORyOvKO04cxPObfIxeVE4ko27sla2gJs0/mkP+NK3xoyITh2kf6h/aLNz7HfcihQc4vxycc1zLQL
eQ43R6AA8U1NZvYFSxvO865VmNxbXFEkH9DyC5MyozbapTWuUI8xPNUBP2+lQhTsg+mIRVpx6Zts
m7Usjmwm0SAMEN7Ri0xT3GqcuDSfPYAb6R2J16ktnesHGfPjgdeHkhRKtVUkd2TV0gzIJyoCr2R5
z2p+oGOIwIaEgT4QHt87IEA57v59x9jy2CHkfk+1FX0SA8vU7nFhy3FHDnmfbSYbHbjja4B+Pl7d
pMthW7P7dEB+LEObZUkp+doIW+IXw0usHlCLPGIwG+IDHziwycro6WdbPQqzbdU65pjeqC8eeaIA
GrvyVKCAJn6qtwycsuRCPBCfUO3S4Xo114S27qQgL2LvlzhBL7/cLLHs8QHaJMd4hIDS3/eckGDU
+MtswL99icFT7cbeK7jYWLZKw3gA4tDFzcSR71oyKvnGDEs597tgPQ3/9RWcyI9v1NZXvcbNHj9a
yztTZSzTbe1vOolnhUeCXqoPCO8n3+MW00uiHTSEJkbEWu6t9kdUUoaycjY7kusaBW4YYpGLhgMT
j5yWZwo5gFnMPYAf81dAI+LUEDFPQTNWz1DjggQnhFwJ9QEdQlTKkzuZBG9IN5ScxFSQHS3zT+NL
6CVGwsx5pKukH41/jWr08yQTg2vxOIp1VB3PVIHK+odusDWMwZ4OdrRTbmisXcYC9tfrsP9aK6HI
V8F3ObpUe6zxOj7PbivojjHR7y/GkEvO9QW/5dM69Lycojra0uAX3CRqMIbF5cD598ZxvC/mwd9q
NdTeRLbO+7VF6AG3w3h/PWntKxVOs9QRNv9Q07GO8O0Us54RI01266H7EV+tXrCt8Kva2fOZIOlA
YfJn1/R923QhLYJUrBb/NmC2W6q2tdk+cW1VassqvPt5SeDHZ9DAsxHbWCoDY3cvZBuOIMbiJpYw
dnXFqAzddmb/e74NE6tgYUliAhp6/Owrzv1ypjXS7RP9XJHUSXc/DjxdXPC+sordo8WHT5bf2cLJ
EEHkUE8I3zeqh+LA+rkqRcJzGE8fN2Ro2czletkks2GCvzopdB577BtaHkXzIqXgj+e91Emp+Uq7
OHZU4APETUTRPDxuZZb1YC1Bq+LO3IC/pHABYbRkTvSdLTG4xnYwYOmVYfxelqpS2rLRipXXTRg2
+Ry34rkcJj2v+CQf51LxbyWhAbv3qEYlM7H3atPeWNwncGBvoocdi9LtZQz2NrVVRK5hmGTRIMhB
5LTd4023ft9vnZE2LgGfla7qeu2HN38QkmDiv62FtzPlxaYvwMXVFjIw+swCoHehqpNQNQGWDTII
sFE8jsp1AF/ggWl7NNhyxtO4nsnqoA8JOYgqik4h7Q5OVWVqgeiskI4Pej0EfmvW5nYcWsQ0cj1p
MAiJ7gEKJXO+O3t7r6RBlCuKHMqXfH6MDPm3NedGp0wL5SUpcjqQh9fLkKyFUMGN11ENypnTH85l
AHpcB64iyr1gobU/SaedXRFbEMgVJec/IIEJDT0+rjruLhYUUZ1HEqwxLwmnkwZS/mfonrIew5we
JV2nDgGVa7wy/1ei/tplOLr3OL0RrhYlpmr9fbZFkH5vZhCUbTGAwoKha5Dg4j+Az+wAmC3OwTmu
mrr61LMdGK4UoprY+tHQ/ZKXM6TwYGshkWrjGjFsqrdf6VCMLNwT9dI5IfpqC82XDEEX9FDRTfxt
iydKy4eOZJCKJvcm5nqvdofIbz26Aqb0owpBsEKg8fD8oqCU7QyvJccx78FvFJ4MxQY37AHqU/+4
UUZ2C0mdXdH8iposItZpD9w60YjaJ73UmxUTBuTWzPhvazQInNCpELeMoW1aZeFlrc0qWttssLT7
w2O3iYzIEpY7XdeSil5IVjqk/v6gO6Npp6e8mXiZnLzLewlaGnOSIhrbINT8eIacR7Wauld9iBBA
z7z3Ebapp6xd1o15ieZ9kdwrctP/qZRJ7QP1hjdG5kYnxY1c7NXJzZTyT7/tpf2aZuXlm5izEJCt
yC48bv/4V4TSFItVlE8DBvvS1owUBgYCpX46KKmEfGSCCQwaiKyP7WQ9Gmzl8HzNTGAzu9uijjv7
pAM71hPpHVcka6x2+aW3B8ptjKlfUndg2my7k+LHf1RlXXUqZywcDHuGQPf2fRCAETr9CULnOO8d
F63fAYkpnjlx2DvbTDBVViIrUNl/oDTV19xF4Tj0PqBuIy3X7JzGUZcSsPoRcITMWD+3pNMNN4Xm
5LPW7LA4XYoFiHP+RfxejGc0gmGbmIVuynyN7BV338mKKblTm8XsEtsXssxR3N7ebUJZ0u4xRyh1
+6SfXKZ/czDDFkkHR90j0gnk4NW3SISA44yx+fr9zVTNOg6dWEqvIE0F4rLa/0yqGl4YgRFjQYfx
ToySQEFkhFaMWm380XDkcMvEncYH4jdcmydyCeCpgG7qwlkskzq1Ef6uG/78S8RU092axrBxCY39
k+Om99Xyt29l3ARlvK59nalhGmrJImVFnfkuvjWvnT7Xqs9iQF19vl5LOkGCu26zu92EOblpNriN
u0X/sdq/YdTTruORPVd6WHRrYHWdp/IFGJpOq1GbijFtqv8sKQcGWF+4ffqrK+gPSUnM2PsgDLix
im90Ot2DxaoO3yXU7KBOUdwhVOhpMeAbueZgpD/4ZghDZoyX8ZzpLavz5WEjpupt9gL37BQDEZCs
XpOIaDWdaoQ0srZ2uiT7zt+z2EA+cVtzhb351DMRFoW3wiCCN8aSuRYd7V8YxXnq6SviwPcgVSne
fozBBbtkryPmZ0oHF9VzSqAvFIs7/mplqumzxgxEfRk0X681zbxdr2ptkKS5hxq6RgXjsfIZ4xXO
20x/BqSZYm+rhVAHOZ2dfCts//9bst07YZbPVFIyOaMINOn9ef2AoXicFBFaPSG2Eyi1p0dAAUDZ
fKOxY/bUaDdQZE6Byx9tuEW6jO2kC9BsEipjpvJchit3XhJDJAEq0RG051OfZ18cYKhGUp3U2Zvx
ZMp9w9yacCXeXVXYj6VOhaIZynDurhBvpDdT5aIkzijhnssfcazKv69BIl8ODUq4Y3sZyPPbnLYd
Yj+//Kck3EepxKlI67aUTpwC25xwrvW+EJJpFpGna/ZNkm4Z3/+m3yx01GKUsPEBvvceK5z4QrxC
+MFFqDd29jauHYvyz7x2VBeZk4mxOe9oYzMkq+CH+CZ9fjDr2TxwmyDFGPeBx95X1FWFCaVi+jUi
HMT8OjzY7jHmUrS0Em+ewKsdq3UKmBJ16I4nX3z7NP2w8ceeKrKvSPvvtjfMP56EyJvl0FsMYP1s
ElARH+Qa/reRXsGdz5HwQRRsw6gg/Wbp+riexkM8/iI3Jc9iFZIS/gnWQEuH74Hnn6rXCfhFEX8U
VVxcjAXoMmRFrYP+pDjuPC5drReXBWOe1fb62s1qBlJvRnTmeqaB9ntpBvtQimx2q6GMS3+IIH8M
60ahqhe+DV5awB3+0ZFIGbKgdNrWcBIwTI26bVmW51rzA7+aIhr48+NxQndMYzmZl0GYGXkn/9PE
9CIzMxwZCjvMWnB27HfFDZfQvKw+DWdUoOa2qBvHjoyMixcO0WkXqxSJLJQrwq/gtn16d6rAGjqH
bDxCiAvljO4vvXyBiJaowujqtUs1cI4cuOqpF0wA1/RIhxDXZtXVRxmpcc/2FbaSc0EDKDyRT2O9
Tx3XI2nATGqMBB0cik795F8mZA9IUhlFRrpqfwimS2mMhl1/r1x5RbpTydSQkF+DiBnXl0i7legg
XxQQZhVQvx12KGzFmJk0i+ktz3MkvD2+aQsMmGzyEqLw2FRxwhtZ8d2lXrsIloxnmSzq6bUkLxAE
XQK6x0eenPXp3g9S8FZZZy+CpCbTiyheVvLnMsFgYIsB/C2lpgpK7BG/ngoOk1GSpU3gXejhUUWv
QHkFp7Jbs16+4Cs4SPzt27nvwSoOT4kxcGGJ6783sRtJUhQVR9w+HN3vnQBxcnAUSY3b8L33NWgy
UQ42YRkTBFMOk+fZ/M3h0oifpakgDzFPoo0KObg8q+9AOWufIQjLcegWQZtNwSy1S0U7GotBYqiY
KI7HNXhQxtx7WBt9jO9Xcps2XNJr2oou95Vwqljnja03bD5QVzptVV6nOjO1ByD2fxn1Xy/m8DM7
JSD1Pi/TjjIYMh+dvTSEYk1li87GKPvBpGewMUC7Rgy6+695ohzV9k4vyeSIr141UnaWkzk4PuXO
tcIIALL2I4c3uDB9XZDm+ivca7GYu8nwxT+JlM1/L/r3CMqULE49uwCMXBccxbynV3f+0vGjuvTM
Z5vCfduz6fCV5v1NIXb2BEQ1zKvxO7h54rPKRvkaE/02FX1V6MaGOBneXK4Jptfv6Dnet49T2YiV
Xtwq7pPQHr7ESnrHTFWexGszAw+oWarBnLYUc/TuxsSvGUz0keY4LwkdImg/rKU40zymygJiTLFS
PNhYkKPLb0WdkRiCZQyYWQnZ4i+dARsHFUVbG3SZ+Net7p1K08WrpphG1F9g4MIj19g9/WDsfdRY
RfimrCP97jZPzrKsnfctia8IpI8Fm2x4I1BN/BNANYNn9xqb2EK1KmnyQH5SuOmBen2M4ZA7LQ3h
373IemquEwIK5KM2xgwggdnQk3d+8lrnnANEND1sVF7MOy1mLrNlqxvWcBIfYZAM8Qc++OQVRRuR
6lkDGwIY7axWHly66YoaHVnVpXafCj910GYhhU7qLPpfwa27OOqwwKgswYHxldQf03tO7yCaGbzG
q3Vu2L8RBBorpV+LMGYrlS0eYWGJeMU1AZPbNkbKTm/cstkvxzeqECsCR7HT9bQQNrKvV+OC3tvg
RAmgg7y52oJQxQGuKJlWy4y/dy2DphVSqrNshzI3W3G7XOymteloVoK/1JJZ431j9lln/VZakX5d
fzLWGVF31iTpLWvXI+l4347qTUP8P2sp4LkGi6IgWprcleiOcTBLpaPp/+MtILAmrQvsN/3Xg48H
PGdxpMLYZubJUGOLfRhN5Y+mG6HoZgnuzzfa+ZuzKPlKC3F65lhIrCq3Z99eFYV5vi+8n1Ar59EV
hSlz+7EOE1Be9/aHXhnlw/mjpP5/CF2I84IdwCTcoka+qkEacjL+cTrUVV0BiiJhzx3iMz2FytMe
Ry/rZ2lzkXHG2TFv2Dd5Rjrw5dL/Hr0K6AlSJHUfjLPPcwXYopKkkB5DEU++Oil0JCddkAzfiF5t
qFm+sw3ROA+rK7OLrlH/XWLs9tpM5Nz1VWMZBFroY3J0CBxUhwU5vsbRZUQGSCbKmb/sPJXfNJ/G
YkcvJk2i+4lG86T41TEVStbL6y2e4EYIkvKossksLVRXrowgjGtjU1HyAaNTz7WbMqpAdjdR/zfK
En54btw3Y9CyPxNKErIfy4ClnPh5x7P6tW/IsFyWUDgHKaAVKd8FBGNqifYRuKZHsGJoCOdjghN6
KGvFZKZiOx6me2qIpNVhCIzxaUsuiUgmVv5Tp6aDZodLwnwsdcfWjDiVGopLN9Qz1KZ7eC5r7rbX
oPY2XstnMx3Wk4fSUrwkI6f5pJPHevVEG8k6sOv5TEAUvy73QkaOqr9UmELjae9vYasXZIjzsncX
TpRIUVzHDIhc8qHQ103sskB7CWf+cxQFkVHOGlN453dn3z2leXyTteMohpwhVSBngBqVbRYkREOE
6MOodA0Z2fp6vGvpQe/TVW+urHpzQYvg18AFyeEp+ZvTuzcMQAbouUrow2G9V22sKSJga34/zxAe
E5l8gwiYHPqbbet0Vrga3pJbqx40pDVZWHvGBgVWtOjDglM2MCfWrh48rHEh55gLtnTMDi0vnhED
NpVW7iO2EDC+3bgcLXr9XRSk3xNkaihIH/M2zyp9pjIu03pjUJ7XlRBMf+P5dqdgnBkSZ4NaqSlz
ztbnSWu1KTQ7PpkqD/hlVZogiuyxJqsq+MUd4B4T4qayOZYnkaPgdDEW4Dpz9fz8GMX+z+iQ5ZLY
fGZGK7QTwIhLBSX5xzwW7Oc4sKc0Als3w8HK9OFTUUPFzZw+lNgOsr/2tg3JpNrIzRz8Foif5sUD
jDaFRIctj+FJsewZ8NhS5hOoAFMQzY4/7J7HKWi0RZ8kSkVigMVCxRgeL00dtp79b4iMXgxEhXtI
iPPPl+pS6D6PDTGbRSivWJv9UNtRUnh1ahcGAUUQdFKs6MaPU3gVAPPVnoaAEQeD2og0ydRpog4P
TqnkFRlK0hFlGYvFy/gZEcVDMiN3NO4bkYXR0qhqthf7FziH1lGHGc+QCPQ6rVP/mPDAjPtBO0Bw
1AtgykHPUlug0ronoU1A223nhUE8BDApYcVxbKOYRpB6MF+EDFaGGBscGCF0UO5CTOILlYuyIo8u
SrqGhJpgktTkMk9lPRAcEN5k/o8QHoZbFQ/LpBYJf6MF+nB0M7CPAhYwP2pxkLTd0bONnWQ7t8wD
+wTRoMqAWqeduu5VkKwA3CYucE1ROByjEMP8g3P5FbgocXup7mCjW1JT1CsDO74TMuO9WfQ+bXIi
ANk+VOvxqdn/n6188gPx+idxuEX8o7uXWvmjjB358BI0vbtnbDoE6RDqQzAWH/K+ukM+C89MlcpC
h+a3BZbr3q2MgTndSTrHZVeIMOFUL4wBadOYw/7QwkWpLmXR9oYS+IJGRw+9gdhDYkL4BG67smTk
RS1Gs/r/az/+eGdQKRnnyeKEvUHSgE8bZGmAGwLU3O8R5qVOJs/a3VDe67DllxVBVEphCEsZXu0P
m21196J/P34l9NRbJWVnAt3X1g1a9vYSMiDZ3fpdEAfCc5bvh8idbykqbO9SYqXm+5ld958NR+vJ
rPPEpsKdy1f3QaU1XBgrurbxkJHWUFz1nrjcLnGBCQpot9gTw0BhVefjV1kgAyIGxxZMX/qEi8DB
f0kIJ7ywjSB3KsO80/NsveElCaHzBoEXCAUzf8lghUVJ0E4ZJ7qxcP7Hn0NmosQI7NYQo9eT5d2c
YdUk2CmvpZFzwE3CCMTKhPwgbME/qnaBMdqO9o0mE8MrfSE5J3jw4IkJ0s67/DqmDEdnbZezj34x
YsLvnwiwQ8fUn/Omx5/1+UVuQHcGszlkhe/VU8y7+H20tytEeCRSxLESB+19O4b4RgIH65JaxhS5
ahUFRkV8CLsTiDq/SYg8gslZxGwPZVciZDtguODCi2g1fPPaL+9FLXbTtVuOgsoYvx289Z0L8Ghn
U8H61xad9t8hQhvvsQtIA2wSNsJtbg0elYs+/lEg9c6g1e66gmaLhhIHOP42CsWM6QgSqDBoP4/2
l64ii+l+rZylS0mhj7yCFdPgkBVEvoVdi0Qebp1syZ3lT0qcS2RLcD4ba/nMkwjIpu5FiO9J1BIN
m5irvE2jxAzLEaqlm7q1fO7W6PHLBnLUve5PTO+7CTP1+/tAzAiaAVwFI/yyrCwhDdbBE4WFmeVw
FDKx3CdYJ1C+EexTTrMzVWw3VfFZcaHsCqaCPLofJf/BZdtBlQxD8It3LcKAv3gFNbjMb1MtrT2c
DpNmnxX7MTkexVjIpQj/NeW4Ip3olrZGfCqud7m6wJMxuEYzfRd/u24sHlukGo3QtreYc22Y8dn0
THtkxdOkMkpvDC8S2Qn5hsWrLm/Mxp4ZzxFwi87Z4RFx72li6CPrxE+sMQ4GMvpekdjOutu95ogx
HSFi1OVdIARWvsoGEWXTXN4FnJoZCiq38l+oTGauF8pzJ2kvZe9CfYQj7GNCC72iZaMh8CRPeEiT
+VvBVemhGtjbC7qxrPWd/qIq5FAq/0EEzgN6BPe8dqEX+B7oPyrxS7nmWxR77icuIB8VHOfT+AyU
zm1Ul3Q/lZawLKFzhW88srkiRCyC137eYWFo5xi8HTRbMRUh6mlwaT6DSz1Ux2wzIXKI7BkZZXBg
bCD80t2I90DG8MdPfYbP3CmnDkB7tdGSh5d2QvqIqlFdP2Pzn923gvhhvOpHNOJC8R23bWS1mxrY
81+gcWYI/dRRis0FQCQkQV/cjPJ3CQdJD/wJCz9eIgAM006orsYYjobHdotyIyOK01u2/gSnFpUq
nzyaO0xWtRnKSukA22QFAvrFqFpdAxe77Esq+T41wGHlA6u57HZHJFy1MyZutEv9LYCKwks0fm18
OiR+yk6tWDgwEi/EQVIWmZBBhrs9oxu+3S052/xLsc+0I5ZaqNuTkWYB5A9uk2ZWtC6S5jE87BZc
0Zsao28gbIkw0mTDIAiYx835BkttvHtdCv/xAqfA9inx5Iybr2yhdP7HWoIIUqvtfY5xbsDNqTrP
hUs60JAJOqfPLSBVsZtPB9zggetzoxu7Jq0+1yL1Gz51PManiOXgNMMv7cdTPf7j6o09/ShbUk/w
GBC4h41JBjB+m8TKv+7vcq/U88dJsmYweizFkcF6CV9Zzae2AJuDIilh2hPY1G9aLUrJNpMUXvio
LObmBjiE6qcw1L2pP6ZCl8U8Q5XEFWX/zEFHVQQFHWbSKflUDfQ1rluYn8kwfGG9VRs78VhPOdba
FhkxIkaYwq3DEDTOKbwf1VveV3eOkBHibYV0liLIHvSi3qLPfo4DxTHfn6J1qJe7IHW//cwBRd2G
FUwzZohmKsHwy5Hw+tIbNE0Jzyn7DHV5pa829R0r3M6K0pr96yuDja1g0BbMuG6/g5DCajOJSzqL
GRI8b5Mn5Fs9ldBEVS0/L4dvrD+b38t05O80XXeMeMTmyB87MtkstnjkJoIGB9wqXyfL40pccXLt
DctyxGBt5zDA2nENUk49NPLGMK/GkSxy4hkJ1bPTl/wcgcS+UWBQ4lN+MH6kbb9wxD96clbBgeb9
4SB3WsJeH9rEXRfQDm6BAxo7YuIkPal28srR+0bsC05jxnhRZYytcnu1SCjKkSDkI1Agd1yYA9/j
SFm4HFxNACB5melCQJFoBQqZeL4qTfVKKFLOxkKRWeohRJXhOSuwGBsB8GKSy0OnhNIbiEF1tsyT
SrIq/fv7j9FYQxJlaZ1anm5nzqZHQpHoVVPlWlwAVtKGpOl8qfOvsBYMOFjjkdTE36VyJbdyOyoV
8U6768GGSCBs2HFY08SzfPaGXDUxOtrx8/egQJ6r6nEAkXG4QNjmoRM/F6D5UhSsENluMLK3IiD3
zLrTErQ7GNtKkcdjZ0UAUH/xzrAQS/aXHAyIAUmbNaJeLLS8Bb441EiXiUaUl+jjliJ02gqkoVUq
sbpKvEvMUQWWkZwR2D4Q1kj08+zMzK3KRUZZF5eqALGsBk8lt8aZ3c+5XrQP0/Cd76nyUDgJBTyJ
mxeof3AIaGEpiqtPnx1ZByn5B7D0vooFr4P8x6GcGK3Zh0Cd04nAM6iEFlgk97RqzBTgvFI5ZyxB
w2wZiHW99LCUANpY5fcaY6l0YVGezRCTCmyT53QYFWW6qtNurt1r23QpwDdOA08mDnPfeHNHR3mW
cGVmldPtQpYtA8aAOVOMxh/CkextCC7YWABowATKiBfgFap3QWx2g1f2FhoFS8Ok6g0bdf0vXuOF
1JSF3D8WVBLaZt/7PMTXjVn8gUbOXjMnKDfgWNLUsw9etcDcGX9OYp9o6pW/Q7T2wknoe2YTfXId
MmxHYvHxGP1x2DfqRQY8Mk+rrHkr0KkggMMPn/BIwvrVXR/gp4mqC8pr/cnv7i3LEHatClJvB/Np
u8gUjPXZ0i5XaMRxxgtYUGDjQN81WFXsqPLUoye8xuaqwAqsOASM5nvmaddesK6ZDfO0BWGNJ/M2
X9GKwKhpFfJiEVTOkCwsW0EfyDnSIkr0AfhtGFd6a9v/uwC1x+SHpQI1QuJi/i0ZoELfzyDX+TJE
2Qbt4C9TS38Flcn28Q2B7wo1J+D43fP4QZKHH8DNs2iNulvLlk76mKpEbX3IMT0fMWBk4E1I+2YP
Foc0eq+S+/Xdv/VQDhMTEl3+/awvKb/I8BC8xr8P4ZGY/bxvuznvze4N9y5CRr3BgI4jOJAT/wa8
9OYPb/bVECPshc7xl8StO22/VEESgXEqghnpLPJY5l4plrRUk37nPmsgTra6Nr5DSeP+T5vHnnJM
HzSl63lbIR8rq0RbG9wa3ivSOmxHIzn7WwBSxSmuC++xkP1pH2zlrca7eUzSEGCGSdgmN7c4jI4u
JnXVstsbNjmAQycUCgdU6rRcKrDpITvz6PEM9LeRUZ9HDJkHKNxqq0tpqW+hijyzbZ/ke2dZakxc
KtEHmnX2J9yduFcr0v0+fQU5NLEdLR1M+0M+K+YizypiUa0h1afKsUOKvWhpEtpopwxE/C1VcAzQ
56ACX89TdmtR4vYHOYlW6tNzRqS9jtIObbdCG6QF4jLWCf6PYv1Ivwk/CaJtfD2+HHBnSCx2En3R
pE9V4C0Uvb1MgNU15ivUFTCkYQO5UYSvETIKsGvZ274SvqZQcZTY0O0r9oEbTp3fDe1dxn5N4Qoz
jg6TqD/V22yLSyfyRgTR2pedyZr/7gRPhHlyEWf6ayINStWJ0lOqZcnc/+reqpo6JULTEVxBmyhk
3R8MccgGFlbnfbRTOsCK6+uM9NlKiTtr943cByQR6UiSN84Wh6vhaknQhGJ9H7gMy22UQfkm89UV
2bE9LuK2TPb0f8g0X3wGhIJt8UmaflB1qr98JRkDPeRheXldUrwO9HyS6n4oMYYMKMhHbUjw4GlE
ApUYgJjQBgjPrviot0y2ZszG8F0FhV02tIB+x9tgB1GVHwNUjaVUgaUik3fYd23S7eKsH6wfot+6
/iXV8zZO1+V1kGs8+EuoDY4PVh8ppC3qU0HqxhbdZzuU/aTfSh/b3RODqKZlnP6NXrWPX1XPE53O
xEi0jnSFKvlVpK+yNpPjz9d82GhhHZBaV2grmpSQ8Zp332JpSglPRRS4EPwaUo2efLAPYaGJhK2+
a5RLMDEFJ7oNOwACUnLjJTlA8rYevnhLtm1V9LZzYQISh/miiu3hs86PZinuSMrwo4Fo7R85skrA
hr3mWSWSsgNwyZgpLNqf44/KFnG/QeNFJNE5cJTVoWt9iVSQIEEB3FWafelHIxBGaYjBStZ0C63t
WERt1rx2aKa5swi7GSPE0v6DV77t2Uwmr1lSmj6100TlhzJbpGfXG9obdQI1P0c7//kYQCVGSARY
nyGMJdZ9ragwDtGRCf1/2igknuveOEe4eRp/SAnH7RP7N0VUyi1UHSWO9I/AG8Fto2lH4uLJ95ss
FlRPSklDN6JD8ahqD7PwetFEWDtnQ/g09cI1/EfDf1mff+Z4K23fz3/W5KVf9FQ6i+ON+uotii1s
rJJMqhNwc9n+4sdCUiPMbazfQYsFdy1GnWHf4LqYLjjanQ25xFKg4oF0mJhJiPQfPrmsfGruhOfC
3LwFTGoT9MNuLtte8ZvLTRaAPwQ+HNggFKrcDVaOm/N5qt+KfHWXMHfjl8/+aRQ1R3i7KHEWTZML
BPlSLNh+OQUeF7nFGedErEGhS0LKwkuu2TEy5sRNDrXdPMB8rzlP5KToTOV2x5iVf+GeZ4iNKQ+X
2GEpc8VeoWEfNzY3kSj1UKJaOX+mdqxk5+nl/D+UXHj+WmTsapb2/eIwGVa1qthyGRJ8fi+x8qRg
nPjLVFFFriRFNhFI/QkFNCcWnPyCEmoEvt5Ab6kGuhAhxL/I0tDo/2hfQkrAe07hK7BdK6t22Btb
E9JhPIAXlJyF2gtAOQYP39eznt0NW7dZosEjq1c+CKWG1lRxC8n5F6h9FzRmdKTegD/k1Z1Z/lHO
/xvWhhyYeBJgh+no/cAXfdHGgTxWbGe7zTLzVXZXZNA+tAVBwAyr6G23xOYrf/DTynHDvQEcxqHh
nPaR3dkFcHdvdZ4EZvTY/K1yJyoXr57uVwajl1k1q11ZBRqQYTYhL9c2UrztHY0Ig+vTT47H64Ai
6Gck33jH9M5L4XkzWmSEZnSapoz9frPhs1cNn+yRJP6mjjaB8hn1DsgQlAOrdwP3bw/JKmmKXD3A
jcu+MlxLz000BJVajft7vlLCqelLwg+dCGm8Uiypl+6owb6ZQmAOoN4eAYKD6ShOMGHitr3rGJWU
bfG9yP8rKpwtLwk4LBcDIw0qsV3BvpdKzhGaIUuOyHk0oJjcWrNOZZEYzrPaIa9yRCTZvUsciuPt
c+dJq1ZtoOK8Ap2HkAN3RsJiFD6dQp1KKkNpWo5ua3UFAPezkcoTLKblcaKww4LIfhuwcAfrIi7U
DBU8ntzj2R+qlRFzZHobWpJVeRQ66ymmL3NrU2GFtQFTp6OOCXImLoguIreULKjKmVmDlA4FLXlC
/7SfHeJc8qHJbm4QiISuh67/OTH7g+fZPYwfcse3TqqiA0lLG3rZic9QX0EL8voAl3hOTzhzt9Ay
txCCnyM9ul3CwMrZOAZzExlFlTpwUv6j2l/nNDpgbGEH3JgfM6Wnsz1luuH9v/273rn4OJXZJgGH
8PqryP9tam0dEvu98imIX7xIu6S2ekhnWSIFoObyX0CN/PcIQjj88Osf5ZhsFLKJ4Bhpzly14CkF
8thdDAWAeTfJhf/iB56ZswC5ulAz+a66+5VHyDHyc/QcqgzVwm+qRos0n4IClPoRnJvAtAwBSudZ
rXeGNT3ZOj0HH9dTZhAKELOdUZaWN5aeXS72jQHA4mf/pKOlL0DKgV+kiSjzkxllgp+75sJZahmw
OWIWd5kkqgmSqfZtw8iMItELvaFWHt2Ce81tx8B23/gsk0bAFT8tkn1IS73X6JFhjgSwE6j9j8+H
qCporCuoe4bdZ5TivSXiU4VoiI5d60OfUBC+nSu+92a+G+68gs9oHuusCmjHh/omzc7PxbuBq1CK
vqpuAnP1bVvBB/W1oMOjB6B237hJkqY04L0hcVNwrfrLOvvGwBjFC8sAld94xM9meR6LTUwiNpzv
HkFArCmam9GMCRqR4CXhftuA4oQk9MyZ40PsIbCSgZM+P6ZD3TapJqOnOQRAz6aFD+gKCnygFlOZ
E7Ys5HqD9rft+Oh5bMUQWMUD40z+MObCpJq7E5BiZdWVNrhw1fRTkBGwf8F19tqIArlT/oZODZ4+
/HX2VKzJoGz4G/L9E2Sct5KZTiYujA/mL6aO1DqU76QfqgYf9xJxjqQg6CPazPA73Si0ZtwNcYGR
SLHj8nzDBQ5nhQlvchp/46fELrjphAqwNQC099T/QgxtXlvoMdkWgkEne9ll4i8yABc7kgrE+aE6
U5KlDJbE43wDIitfXZowDXlHRxSBA1ljntKIJq9i4mIRyJ3pdX8U7jS5v4LHgEAGgsQ04Dtw+jIh
usMQqLVuHY9cm+AZ72qULsIo1NYaZpmgQ9+9NYkY9qZ2soodQWmW/uVEuSafckHfBGUQ+oGrs7uY
/9PMDZhBegHdlzXMqLViymM5n0X1jxktlmp2uzoGxTbd8hg6IM8ExCGUNpOfvJS3q5ap0zEsFcOw
GwNrxZFEL+isP49nVhGrAD0YL0PJl76/vi195Y54hKSWrhF9K3J9eajOw50VlSE6/FpiBpumNnXX
9XeLvbFtQVvH8d5qlR45463oSha0t6ttaww3TlCXKeaAWM6+GoHSPcU73P9WnhWFJaSQ0AeiRZgp
EoKN9ySrU4bsMy/vhRiKe848/gndJafu0DPLULx6BzRN4+qerSCownH6qKw/JN3HIRYlmHNEuoF0
v5FxnGaGX2iYuiTTbtpSyr1EbuhrxrxCcR5+g2qHZR1YMyh+Xskq94CmAc+jMuXV5amLKt/9nBZ0
6GvMaIKgQC8ilO31qQSKIfqwWe1EW2XXOJz4mib/oUhd3IGdaTkNJK9ZmFnjPi94Hkox3gvN1ujj
o9PnOCA833JAsDAkTH2BjuGhUWR+AwJ42pcasgTSZ3uYtnHrIlCqwEVYojAynEhzhrBf5kGn3rEE
5B70LRvuNR0rkCtgZ36jjN9jKbbyFsRFUjGuWx1Bh4R8cTIQZumRNHa2E0HLhN+AnUG/PHfYF3ic
/zTuJswrj+JS8yqFAmNRUbGUEiyYpyh3d1Gr6GRBHPQ6aOdqBtiwFhIp/Fxs4rrDPd248vatHkv/
E5YZWuliPTeHhO+xHD1wl569cZdebj6KaEMsjX+X/ISdoTajCZpCZ6GqKVH1srhmLoi23QmgF2YR
k6HHFLBoiX/E5cc5HbGtp18x80du+Vuea1jEZRAWfETV2X+EMg8i81Iy6Uxuhih11wXNQakMg3mK
wW4liWZj3gA77pUWNRw60GNiwvJMp6pZqseMF5yn+9w+O08mwxERTYq9DIMvLvFJHp4Szauy8FxK
PP377dnskYstCK5p0uEGqi8wZ0DdhQaSt2y2e7EXyuYedTogujSFDxY4SMfCl2TmgfBD1rCxCi8q
yHNBuvFM/yPVjctzodyIFNAa6BM11EsoomOsaOT74E3Rnmn5M2sVH31iyrGV8s1vWTswvbTk3TCA
XTpyf4AR5Im+8XGSr6EvXHDz1OklX9+aG9pJ7OJ+2nunT4UavlRfI+9jFYv+2BLtU8+us5dC/2De
7W07r9HskmeoxIlF7I/EfqfoW4kDJbExq/b9K2uL125JaBf/MbsHrc44M6ayXnAILmsi8RAO9YmP
B38gjQoeQ8HH36VFTjHXi0vP+Nl+DwbPyLnGo2t4xx8oV8uPQe0d/b5iD2KzfbQD1EFeQ2spCPix
bAR1f53wKJ9DKAaF6NHQ587FbBCu0BoNR783e6brr9D1p6xZ8SurtY5NYLfYplGMkar19o30Yo+J
e/BPnKdmsX4Yh+f1RAcE9iK/isWwBr1i7i5SILMvtF3IaPIOLFR//eLnC1LiuwJzGCnN0CsW4P6L
upxyMBAT6vRCMozFnx4BiCIz3xMmyPCIahqLPpkNQ1XK2DHyJIyc8PzyMQvoXd6G0bYHlpQr5dnm
Tv8A2Q5YCpl3MIO0TWmPV+sDpO8e4AjwYglH1tOdNR5Pm8GX/mkYNYaGeU8j8fw49os+CteVq67P
0T7awP9UeU0Ex/Q6NoybVReJMuZz8boinOD6xnSlEGcAr/Sr5nM54i99DxzW1emfbnQONm90pxgf
72BlWu8wcOFIZ5pEPkYARcITQUEx9bWYrHs3SFiNUgNC51UYtjvBbn0H+kiV5jJh7LL+Ck2nr1ZT
r5RVszQlAYLxz0rQUFiMk9hMrrG15pL7V5kBhnIeAl47gArM1GwLoQOpuHjvlHH3GNB5ELYY5/ei
QDpsrIpVQRucp1Wqmsa6ZIiYac0c3ylnsTrXKNzP9LYUqqlGc+Q9l/JnaaEd+3x3Bpk8LpNYIpIY
XyRISZLNGJ4UOV18W7LViKs8aWlTscX/Zx8lNIf9/w/DJecj8z5jRqYci58XbB1mKW7U0Y9Uzkvp
kIZNppfZBngve9T2n9cZkTb9bk+eTcX7LzRFKnGZwSRFKZv4GxzpCto1kDgUWITul6sWE3huOisY
yxp1qRxyukvEegXRm2Br81YP/+yXkwdSVMMaKXNxOS+qLPFeEB57Ks9kIV0FYRh4EsYowBvemPJu
Di+OL7hsSjGDyLxFDJMGhX7g2tscAomdAwMGoECX72078Scpv4+XS6YIye8bYCIdLAs3DUsAI7Tl
JitYitFN9aEwnaI9VvYo1nb8QrqU61ipP08qkRdjCq3m6TGUIANRuK0EAUdxBjTSjQpobBhAP+9f
8+ZDQM/WpX7XTKqgeqfgQZY+v3jd7cAeO+uHSQiFjG+IR0QxADupxv64VBK/yayQScFgUuMMY7sZ
pjGZHDWhQTDRaalUE75zfqQND6Eo2qiWou6QUB0s7wLxubRYoKofpU8mDswVKnPyRtHu8XXR6a80
A8YGY/AMfoF4vo77cAYGNI9Ml4MJqoVSIW7LNes/D52fa7YRB0DlDz4UqxG0+UPNE2KJRSGBAWMQ
M6DEsTeMQfjP4+FygBXTPUOkVRYrKJQu1qP10FI98cGPMnW/W8LyFXGb021wmi9wiFJEnHkri4Ct
M1ngUTYAlWpZpVyLOKx+X8uZdY2bCbzu4sKdtB/mEdbQ/xBezOZ8izTzxMuTsmFiZt1ZBZR+4yGG
vDushqLn5E73SXscZR8pEqESlJskwzzQMtLFuB+0M90EtZFEX5c7WtRa/fLtkzMe3mTgksHVzjdt
4z3o7WAwkrr7qqiZzer0Wfa/XmASx1sbZxFKuvw8u3U1VAgZp/I37JMl4d9XmscT4Fj4LdGII3w0
upMrPe3sw8hIlHDZIN/egKW1W2Ox0PkuU9bhSt8Qe0y4RB8VBX0qbqyqQ8LhcVfLHDhZAareBehj
B2L+OQVUENwvw1FxlO4J7JynsmBYytnJGKe41Yb5D2xWT0nLxE9NnJxLTQFXmfQVf9120fyad/1D
0TfFSyhZqMKf0DxszzKxE9XUhrsxdRq2TN1mC5icjyuszwTM+KP2bwqvLbymdXhpA88JfL//xbdv
uloNv+Fu/UMm0L1wgVRJOrN288Zpgo+6gpusZ04efv7V1YQnB35T0S62WA81CNDKrdHCZDr7BDA4
y+1pGgicJg+mEVq9PE4hHAeHtsSqErwZ00HFuK1iLvGmqh1EkiMjK/v9K7TnKp82sF8l/mP3Sy0r
/DxnsSXphkUHGUq158xmwDYtXaFP7+nVTuEEw0XE6p/BXrU5rwaFMe5JskIJa9N10l2+5oRoRn5O
B+G9Wb6+wMp+xYKW60uU3xXF0iLwr7D45z7wZTnILGoOmdwhKLcuaxtI0yVZmstnVfK5nr+i8PqQ
uzEyuIQO6eET73aNkku7VGw61O2fy3wz4yisNS1pZjyzyD5r57la0GaPHsahsp8iZyY87uT1QHQa
sh8oT4rM9KTa9KJSwuVOu+KIYPC8PpBTil2VHV6VcQJqiswoqU/McYXsE+oga/yY00NSV2G58ZR6
Ddyl+pvu3TSgrG7DM8Q5c2HpKWioIMQGDSp8Lkx9c8VWvtbHE5l5BlJKvE0VZZK4/GkikK4TfqQ1
y+8tksGqIgC4Ib+o82xRQh+knejrowGpRA3Lsj3OWaYzUqj+vFefPDnjRj3sifxFs1WiYC2tz90O
cRpUEoJs5vYLdPn1bdEFyu9MiEvU8nv69Bxkpxop201rzmADwS2/avypAF5LORb+hGdNoPLYTZ8r
xJmrvYHMtt+oZnoEyEOvaeenyWXDQTMKZKcY4t1eLK+Si+mM0Zlv1Xr6S39UuC2aLAWzHwd0boHK
kjrY01dCEjKnZfBfT+EGQguPz4bm1hddrZ8DKaiOO7nPyBvA6O/dlWqnRoSKLeENsFGhNc8CTWOR
GT3AtuDmuI8zrRWHAbqnYkKRKca9iiPsUT3rfOh28q1/waPQQkFpv7rr4Z+DcS+IsM4u8VA6zHcj
urtSjh2bQBT6nbMw027N69SkFXCa145AM6q5mwgl0rE74b730AD7GDO6eupHi6UeuHBvZfmd2Xfg
jkvMkEOlbIpjPe1ESVtoDxEvvN4GUoNecmPNpoMjfEsaJi7Ug7ugy5QSTAg3q1fPYbsm05blnpiQ
O3fdUe2a7qGdrTrGhdZG8eTSLmpVyvXUz1G95nHgoCo4bxfd3vMcOudZyFFFRZH8Fov1/E/5+cIA
3deC09h4kVBxftq/08aHsR1+Yr+ryImYMWYLtUaI5pnts0wswDuKV12AaQt+V3MzzVmuyioz6cdR
2Cc3vU3xqpVAwO9vJ7JVwnauezH2dPhd0jmlpm9T4RGm1Ji3czG7pAWpGXEhOWCuPAx/YTC1Ww+W
SNHVdaStkBprvCA04f7OtEZ6JL2NRRcDdnLy9QlhzWoUT5N1h3ByCgoLg6zj+75SpAVzV6H8tMYZ
TTe6UNiZCLK8vyVzMMAUneHp0t1HdzVqgAj/gu04x6g8Da2P3p61U+0eUOsyxnimZpUccylWZJ/m
FV83minP6QbFjBI4FWuYOyqxkQB/h0Rp6V4H0u374KfhDf1Y40lfaUy3s2i2isIh+XW+nllhfWVn
ZNcHtdQvS6YNuUO9qazLp2JRDXaw3JWCsWU9z4Kz+N6CyTMDhOglcueeZi0/5+BsrzHYtt6IUm5q
wtjs2SSs+ot1Oiy7byXEG3pP4gIZYQlt4my02vTL1qbvxiwiSTAC3cYy4xrU2mzK4XfWrRnM3Uq8
RP+n5gZkTQ3DQI5RyAFXomjX/Y5+DZaurh6fLnD+BRnpypv+AhlainKO6F8Z+6aawyI+xxv74aBf
BcBIds4JIhLbgQaw/sij8weSZehk3fuYikflRPauFcMorElGdaDI4uAaJ5QlREhkEYdsZEC7bAnX
zKjur1fPmlHbktnY2OnALI/ECFcvldD7nms6zH92xzdefPFFWTVtjRmPCcdu084TKNRgGr2GdQMX
GuhmrEcX4E6qbtnNSO17y07iZ5TeAieBOfR8aR4OZbn5BYX9Dc+oRuVqnF9cgjvmJCTJoERmbz87
iJgkvm8eTVt5MTiHLaOoukhEMZ+OuUO3MAmmGQRGY5jEXmrztXFyawA4cuJkT0uV4U/aACyv+OT0
GqCEO08NokKRiEIFUz1l+u5IJ8d5r4LD5yVJlDuP9MuK6nq0Vqjgr/0nbR1a6dvTIekAS+EzJi3n
+rHAZPm7xMn7b6q8txI8y2gJYxB09x4opx6xLk7fg67P5rOpKxq76unkd9qk8CI/6hisCGAKm675
/M+5P+H6HVvMzyUD3qZXn9jV5okiKhjGpyp5MC+Qnhkv1hwoWjyn5yAk3JL6migEv2vAdCvsT2kf
UpUjOmOwm9+ECoZn0/YD6uBV40rG/xd8aPDtsPWEJjrfrDKdzslBkST1klkPjPoHmMl0vJ7wK0Iz
ueMdk2B6HqwMybxDzudP9MjPukI/dVKpRrR+QlF5zB9zG2AI90hXKa0P6pI1x+888A4DEdJWCSIq
6Dy2IuQg20NJ71Zzys83kOFEsL4RUB063bMt1Lrt3+QkO3EVsmn81i06pi9DoXxGOX6z5oQnoSk1
XuFwoHLo35v+W7qaKAtA9YeX5Yx38AAMBCw1HAwbtOfM2oGFoocgQlNBG82U9uW2yRVUblEftSJA
8vpOGnYH4U/LesaYqI6bEuC/O1Cxo6Lx07MDXn8kw1Dsy8oRfHC+DhP/oUGaSbuluTV80EC9r38B
jfWGTOVbKyECbnTRO5ZG/Q0Bl+YMSmH2oVWSEEk94/++9ilNqxJVF53R0pTaljtxQgPSI4Pdz/ik
pPIE+wIjWr5Z32HL7kNgYE8o7/YmKRV72yC9KJNyI3ukPzq7l3lT710j3wWSmUYGwiYq7fLi7Jpz
nMMULTX58nSY7lHkpiMSQTQ29r+9DmhKyXU+MD1GWmiRu+NQaeKjwaDvJSpLW+8B9UZcqCw+wvy6
a/FS5d5bwyqoW4iaSPdug/9gS+LCS0JyOObZe8Mk70JfBcXzmkOSkDLvH1dKCaunC1rS4al2F1Ez
iC/OH7V1c6x7QjufknCLxNHlolfrCcbt239j0LnhxtnkbBaaljoSOuQDNWX+m8XjeCx9TcD9YXM+
U9h3QOakdFrNbodCQGoZ2wEdwMvypKp+t9Vo97k3Ge6ZhVPbmR+2B0ITXYfcla5ER6EktNDTSpT6
jFBHbhol7Ai65agTEebPEg+sJIzATARFZs98QrzfKs33FkwkI7TXHQ3wp93frCb46WRIfIkYAgHJ
SjvGLdHWezciBybrW2oUvk4EsQruiWrolNyRi2UcWh/2h9OhVbHgno4fFDcA23Ue313YUEao6Aiz
39zGV3zRmL3Im6DIsocjzVrrqUG8OCH1h1bIl/kYUaWEpv0SolnCdVtO0Tcuic6FOORNAljh0Rm0
tys9/bwSVdHTEJf3jB8YAAQARHE9tb6RfQE2baF3xNjxN/exB/c5R7kacOtm2NRnSaPZeMWbJDh1
+E1zCmp4t41EflAWpRmnwQ2SkBp8XtQN0c1ZqXfYgXfNq/OY11CyljEGFOqax6wOWzikPa0VpIkQ
LUxCyTt/3Bsc5qqhYAg0jOyUI3rSn8mio7GJpGJI7uMk/pn+M5d/gnLf1pNj0gPghc1Voi28XJZB
W9Igf9yh4BRV8Eb3DqzN7UmUOpQfarXk+mek/zLMn3j2KjM0GErMTjkNVbbCTkf+TAO8vIaOeRZo
XG/l47p0z/iaKq6N5b04Vz/eAllU8StEBKvVO+/YX0gK0pvROhmFdPr20ps6McHahDrFcF0zn9cN
D+/0hCq/bc/aprEmc6KP+OKsUctd7JyBEyHZXL2FSOgtTae/h7X+BosmC8Xzz6KNAwKKzyIDqRu1
ulEw8Ozx2g+I4owUj1Z1u5E/c1OCNYBCnPPFzJ4GA50yZp6Xz4KghmY7LWLaVTtBultUOl9Ipt8I
ljHAq755a3b8CAd+/ERIA7L5nusk3j2aL1tET67H0NaMbuWUH0smqHI2x2VE4/QmVZV9bqftVIQw
B51FcSwM63czN6fcvyR3EnGlm3aj2a5v4Zemz8ndg3RHaEUAGi4aw/ZkRPbUqI7J3o9QjJQgcXx1
AjMUR8+j/ctfgl7c8fwTxf1Z2AAEy9aRXbW4og6mHXm5pxJqlSiyVFsphRDWhtsETHr7RPmuuR7J
b/xH7ViBRwSGnjuwZeykxe/RnaRTxGScGhvMto9AAgmyg79lMP4XiUgtJooAG695iGBhw5lgXNCx
NVOKuzDBiilw71I/AaX+450vvdgW7zv5Yck7wjUpcCLECXfzJPDEDw73o10QUAp6GmT/MM/F+LQL
0JAK3XRhCOh0IgnssGbo7T0wBft8rkuV4jlafaZ+A3pK7ddo9gOxoT3AQD60/SJpKH03J7SB9cJ5
GdhM1kkvcxC136yRulBhlF0rfhX5hAjflDoBVOxWpmAjf3/dJkrEH3ioDCUOzMlaTZfuFfNwxE27
a9x7U1vRwlLxJsi9mzv+MrZX+JZh9FAd8N0g4wWEmxLWCmp1RjQWTTJVDnkSjNc9e/vAzXeLKmEe
5YbkxD1/kW57Gu+hQzmbRUVVPbH5NjAOKoPJSrjgAA0Jjm5DS+xDLSnodp2Ersnx8o0L0EuuxQUT
bVzU8jkrqRc5vFc8gxuV/DaVrtupqcmToackG3zEF82jKUwacadhCd1vCtuuyxJ9DvTzwa2A5I/e
r3K38ZessnITVVh/5X0Tv5O4ONP1WR6vKAtQF8XzWAkA73kPK6COCWBxmXHvOONe1HJ/j1ZCl3nt
+0lG5z7aEjCTNLYB3GQOsgyCUylZEhkgFZclNNSYD/iwcjKdDrRYhUvMfteBPpl0PumFVxAVOHH5
01oF3nfri+JLCc5kjxQkQe9m5A/q3zIURC0OfpKzUHW94lbCPF0PwI76MmyDVtKCqm19k+yFVQvs
Srlkso2DzSc0yvR3vHrLiCf6VIuN1Yzcmx0AaDQ6H5fa0Txu5Uz/gicjPemGpMp3hqCe9DqmhOGP
Z1wc8ZoJbLUUEnt5bQckYTZ1hJedPN/FN7dkiH7FuzPxPvctpABov4x3ZeU5XKAq+Ziz4c3wrZgW
6v9fk+6rVZSbrLBkcurRK1lhjeyCzX4cYGFeuj1Hy3UrDCGXnOT+X5ICTHvxN+GPEwH8VTuiFraz
hYtNSdAqxNIHE0SCy7LWCT6R7ZMc+hS+3wB2sda/2Cx8TBM00tQnSo/e2mzG+TWHIe+gj6BujoBb
6BTT/NsABn/mkYYMsWwDV3da7Ze8MKON8MNuGNWcMAb7eu9pHVMFioqfviB7iwG+36uSYsJHuCx8
Gzi8Am1EjWFQXpXd/wW+o2ZMNLgVz1AHBWCEb5M6A5b4iEpsBguKtQV68BNMj3WaOD5inKbw/46z
+nXMs4Zh4KQ4vVKtE5R787aeVvimpRZeloYAarshltcxuF/amHj2AYe5lvgItNQjp3P8HaGrQf4A
7jmJhShsHq+qURgX94eaPr1r/1pTbchKiuSp8cg4rl7PuZmT5RCc7/cXJyMQA5mika4brgIuCnkW
8EryY2Q6j66qHxkOhjeuO/3lTvJ6NrCXKm+GQ/m/I99ZaOvGMJbOzS3udLFAA4WUjsQ84A7zfiml
WuyD4k/dmapAAZiHXOVpIHx+DMyePTYukIhfHq3DUE/DlrBa/+4BPYzO2zeYH0030aFDZpDYca+H
7zXtgPOA4nosP7kYQdWadcdFSq7VRPiJnFgp+wxO7X8dqseg/pIkibi6OGOGL0sPOPBZivw/CSOi
ZkY/87h2YaKsOJ8JDF2/AJfvgAXcTzDRcPMkAi6n9f5quCuMEv5aKJIXmWWnKDwxYZTK3AaZL+a/
NvJQZ7FMWzSVIXomjgvOJLSi9nVHoYi51Cmp2v1tTii2uqGmNiUYU+U3N+vridlJbQFPd1GIZg72
JwBMjUuEHB63dp7uaiPmcgVUQqGw1F1M2IHWnVtOsXrAJsO4lNKcSQGnSM4kejTWaWaYzY2sw9bL
wP0p6L304GAo/LGbwJFivZ2GKbIAtymoWcCE4R+QiNLpvaWudVNrVdruh2hq5dacIeUSaZIjEETp
KsT+j/SER1kq3IZdk4eryFHOsPAwGd5Fs/llhtuCeIPAVXS/j+o+BjeUUP7X1vdd9I1HuLReHwrK
2tv4aYIILtHOot0nNVn22YnPzcdkMOtGyA2p3ElyUH3LqeNmfVsdQfsYeBHAiF0bIwR4XhaCvVhA
H+wJztzobBayIl10mAYX7rrq7gG2BElhWZ68Hx8BPhVg9J2kkiMEkr/7eb0+DlNJfjS0Fp8wPWrG
n3X2OWSNHp5jDVDgZSm58Dug7e0J2Byv08zGWQlZSObo49ia3KaGrYfMD9of1ywIj9gQeiN3Wj1y
Ty0QQnPndoA7QZUG6MpcQU5zggnGuT7tvDK3bu0kbBSCB/krp5IgZLcj22Ancq3zcU/Kd6IH5f9S
5k7pzZUycOoDn1bBzLHNtuWj6lzYBMv/wX+P8U0S3bCx0mYAAgmpguFk2rS66e7M0TPrwb31aZIv
G1JRFdIracXkMOiMa1pv9v8a0RdEOLShhx3jUqUQ908qR/SCxVyDaWUctBO3fzVAQb/I93l+yLME
C8f0c5+cuLf1V10Iss+KKMAfaCBlxr8ror0MD0POgWfNcUo49CxNt8MpDI70ZXF5lke5jP82gMrq
RyOtWtguVzyQ830HrLUGFnbxwPAR4sEtpoWJbEcG5Ax8fAPBhs4LhxiG3oPcC09vk2/BanAWxgfJ
wAz2yYzoKZY4+YZTA2Fm2HpIRdx7pjJFNj0yAAqsqU9SMxfq6OPIIercqE1QH8VRt2ETM+fAgqQy
nSyfLNl+UR72gdLg41jiHGde0EzQpef3W8EOEQvRw1B90JocUyFnsta9ToXQnsO4WI1cRSrrL/H8
f1N6v2SAJBpB0l7rkfjJJP8rsvptbyHz8T/xnfIJ9OSg8LfBlelxSbhusJheIJt5wG0q1K2pYv7Y
xVwdZymOunxKmngZ9tbcDSD6zhHpLNNyRkjOeT4cg+jctXSdDjWEQk87fgOnGia1mkfllxoCzlvj
xv8ta5/b9Cdxxy+4BblnfOc7JQki5puvMZDssFV7fPSYQzm6i1B8UrPw18LjQLQED1vb3yDCcjLY
wdQzUN89WHgi0oZzm00iB5jvc2+WE0SKj2bzUJg2DAdnoqdERyBKFZLEkpMDD3PnMb85zUTOb8J+
XuKlSXQAOTl4HecXLq+ASl3NiDIGz+8sILhlONZ1Eq51oDv5OvCCavY2Ww+GGmZCFUP79UaI9eT5
2MGBSaHKMTrkuIkd2+rSk4RnC/BYgHLpC/ELE+OQkyYhYU+zcJQ6+Nkd4hEqnKVEzaF/D79AhjX3
g2bwAVXCfLECSxtMkm/1LgrZe+L/RdqFxdDPjvIoriilDjkYEbqp4kmCbAIFdUw+Zbt37A0cY2k7
CvtFPtN2QO68UHryzqXkR/qQEeqzAoLe43KzxBOSbFpp4QZrLy25q7gZUZ+bSFGLC552v4c1/Zrj
0MEwRsW57jbik2pwlO/16PubEWJoo0vl6gjaQB4lVXuZ19E4/cYDtPAyix38QUtlF21QEmXtgTRI
RGq1QumqmFuD3QP5e7v5u+WqbmBqCuC1vpR4EWFtpMJpklnsLaTuo+J2mVuQF3pXrsNf3VsK0SUC
RPL3djxh8bqdpx5152qyugvwnEFx0trckQEk9s2W3k3wdzg6KUu1vJDWr0QSSKvTi9COl/o9mDur
5W1u/LPUACLDlX7m/tlQr/100321Bnag6cHpvmurtAy6WZxRE0AZsMHkRJz72Pg/6xhO51LbQHiS
b9sqispLNss86NFxxpkumXngwR1Cj2LR3ty+O2S6MWZdNvbH1QmGpqFlWd+2UsyJFFym6SM9XamP
BzjoOSl2c9PIZmTshFvmZzqke8iNLrDGBOt/oaod0T/GK7cuFMs/KOAT1lXwuuKlqWm+63EnF4jK
F4wML+ZWIcnJWq7XSMpHZcxImB9gSW+vqKcp1KX49mlpiqwROrSLeQTRAsNue5bJYXpjv4unoBut
/hBaIQm9/T9SIKCtCM7FqQp635FAzTyoBdRmWMo85uWbPhMtfTNm8wCJXBjDMr6213qA1rmTtcnE
kPu15Be6yWnuCaZhNZcKhkqrzTpoyP/Bu27TnOAqek5+8cWrbWC9xAwLKLvp3hlsiQQ+bPqvOoeZ
W4niOmEpTLw34ewstGs2Z64va+NqUDC7Fu/fXu2Fl+2FrDrRZxiJpTXZSK5JJbBkG62TFearrH8W
QXCeugH7A5llNxZBYQzieQHONnPYvc4sp3BXVe09GeLHshjwOERtM1dtTmE2k2QBZ6JABHJ6JBx0
DSDh/yvpJbl/taobH0uaFFThcg92MiFaEi9oJ9IOWAYH+yQn41XXfM5pU2DYvZJwMJpEmWG2MkWE
cEpDNSrHe+Kzs67w2FZwqhmNcQkJ29+lh3NbTXdoNM+qEdWZzb+2YqfU0M5Cvl5hqaohBA3L4WPh
UGCNVEQ9qafpZbr3l+oliHLRn4HgRvgoYhOvjUc2jSzyOi9+HZ0TLvr0ZJOp+aLkGd8l8qPNAAXQ
iPXLWLLIV7gy1bo2KQDTGuDnT8/O308FQ/gzJQ3zT9lLgEF9+YilPedTsj7WVLE2A0F3kaIHDHmX
L+pyJzHGP6C8hmwDPqQqd+4OFHAKEoFq6wlZ/iNc25WRuo5SBSEmZZDw8iorKrmd5EdYGe0ly+FU
Hr/ArlL+z3CtCojOcaiJSaWu40LCCcbUmJL1xMmkrjACGYImxln6FfLDzgI1ARxqlguzxqwV7vsb
Y2zJMmVOL9TZBMUSmaB4BMMcwiedEBNl5cUq+2EgWydp5hGBorHU8+iRWzfBUe/orsqeVWEH/Grv
gHWjeTGqbFGoMF2N6qAcjn6UbQXnSBqyMCN9xoPHC5C1pKbq2eDPT/pbdT9548p/RzCeEZQhukRa
StPxj9J9bt3dDVcohIHtVIiuIkxGkkoKAQj8mSvz+HOVcQGdfYvRNfyw01ktkJtAKKHqU+wQW0TX
FXYpMU3MbcL+TddpP0Tb4jZYbi9FDR92M4c5u1/unv5CdBRA0zRCeGYA09AoWI2UI7eAErlgvfyp
quwC8a5TCZNkN97EWpI4ROAgs+N3n6JddBVxnVQryR6YQpxMDMCZMCPSVk5KK88MrpCuP2qsQQHT
BDyIXxeO+1UPbN5OoRJK1MO7EwsVLY6foaryPgCFMXsm4s+dM4P7jbTuikcJNBWhSKQ7SOuqddcl
YT9Qy4+ENTUAvro92T3UHAHuZLawo9lsubZ+2azXV5ovujS2ToC/anMkfDLuKj5AbAuPg50FQQ7l
ZkhPUSMCX5M6HBZAM+QBzj0C0hvogDHgZtozq4sBL2nKx0UgJeLr/ePcv+ZGfxyyorq7oECxNURl
6ny5vC41GV12NNLmeslFRhf20kxKJvMnAlDUl4drXABfkJP3fzTlq7nXdghZRo2om/1uxBnHxCXg
CtdkSdlMTyQTRvi9rrjOMpRoIwjsQZhevfcsglYHGAxrFtfKTSippKJV4/dZFm9/7zNbCGHQKBSO
jtTwQVqY/WueMgzfdmK0MQn5CjRhwXy7hXxao42ACz87Ok/4t1isAyfBnE8VCE0nZKpvb8EiMYOc
ty5iRADCOSeZA8sGArGhUZOPATj78t4Rj67t6Ubc5VBw8Yw2LGQxhpi9yELwsPDWUuy0nXwLRtqb
MkUphlLUVKpVU2qV+ZIGleKDqSLfG6OgMR+lJea30jvoDjhY5Bfn/tcJQ4FpJhEYmDBeNWZu1pY9
uJnk+4fEHln0qV/Q49mAJftMegwlgTYt5ySQSj7qJfwP94igWSORzIf30O2m47Wz9AROVhKYwyeh
JMLD98sG4UusXREIGrMUGLUW9T4er0u5dYAL//5vBg+w+Ai7kMb3SnbC5PDFGiEEL+ier/dm/HRX
IpdZAQeheW2TK51xnFHlWnA17l5hlxv4NQg18DsgRa5hxgvevBUI6K+UHZ9KCeSqFmkWM0C0gdro
lwuVK8DMOac1LZMEC+rEx+Obvb7c/kyADWaBs75ouDt4k13nrU9/C/eAkT3USgr+mi4sPAXw2H5I
ieTBd48giGwQkSK+vhu9SbAWgUMWnXDiw/ZEAsu0gRLH7BghWdY9QACoDJCyXgi6ULR8LZYG58q5
N3kyDR54PmCukB7o9GSFlcxOse2RDdAiXA2IO8XBEy6qlAi5EBNUeWeYJa17gucqAjM40OCrsHVB
FUp4KTjaYmhL4LKfLSzJklgr5FCWb1w8bTCTK3EGcb0G7G/sGCyAff3+t+2aj6WRnRsCzmi+o9tv
LiCJyJmK84MdOafwSzWuDNUFPLNgcT9mlZYK6zroKDjE1RJul85RJvO3VklP1Ru2Tjtf7nHKY5R9
2Bz4ZAcIIMImuknvi20ZoUrz5XPbouLStYqmnnyrLNYJkd/YW164IZ/nddEU6t+ZeIu9/NtxO6eB
KRwuH3iskKbJbqX3OaNy4wS/Q+++1sPkwZQ3k9mxZ88xS+a8ZHfsh4y4L5Xzewth7PHhKvOvXn0C
uZagIZPNi8KuqEh38NNanckZVg4E8wvPApvkqNHYWqL958jQQLdM8+bat/wu/XPmmGpMvy+0NJIQ
OArFf+4Zxayy9w2nNc2K0/cKCEEdK1/bOCORmLhBq8Z5W+RXsGp0MTIqgXr7Aidbgkww02XfRVs5
m2Q5VwVQXFH+wpYU13ffR7r/5WKdiqecbtrpHTGVWq5Zsr7giZCo94sLKSRNM72lrpuFZy4RysiJ
rGhcdozTxnx+/ThmkOSpwmxjjW9Q6eSYGWbepOTFwDiWK2o2MfwJphl8m6s+AWWRl230FOi6kwo8
uVlHNzhdD6+YiURRhj8fzQibIHkc81uWNU/T/KEhSCCMXBbn/hw8d6wra7SzYArfMauSuR+NUp5D
JFG9LqtDmLoVsvTaVJVVg6zqXMVR+j29f6WYu9MU5ubWcyPJMIzzIjK5gyJ9byVM3Bf5ey7rkx25
9BNK6HcUEYvxZtgSPMSyV9Szh6W74sU7VdEGiMSW1bBXpuj6XrhwpZ5cynmDnyU1V+KSRAGDDuBK
BKAP7fdSLg+wM8CP40ivhbB8BXcJPt3ZP3KzuxMeH1NgBUS1eyRT/saCHMjmbnpTfjhw3Kq13T54
0VkQWVZux6tqPouDZOLDSfYhP8B23h8dCgDaKaQGIcz+zuw4B+jmpO9TFoyVmOsMPBFYr9WDffj8
u15pcF5gP1GnKb91hoCrC9La/ck9U8u23amiZLlTaSU3eq1qxHVb17AKi1JIih6fevMSK946fY2F
bLBv1SElcSMP0jtXpOPIk224SyrLk6yc8tZ+8eEfrkZB08gBnAqg1pv62vBaamOP0JcjmgqDXDYk
aIGh73gg1nLFMjX/+9c5g8KtftoGM1opFt5Ixfrz+ODjdsKwUjC19CKsQ4Fp0eAjhG2eoDh5ieR1
37voFDfEmVePaQpjGalQrzdQ5LkA/g/Rts7Oez9lLril5Hyd52gs9Rv4HBJZ/Zi0clSLI6kQVA+g
9/XtTWjjtDGkXy/pkyWlBLDrKfo0CQioNAuHJMICRiJ1tX9LZABa3LwPJS00rS8n5Zr+km/PQNm5
zKl6biGVCCawoBynI3nU87Xhj90C99woBxwxEaStmhHsjwbq7hK/VxFvK4LPbwQ7Yr0KoqwcyKzl
vmdJvTxom6HifJySaAg5/BhUxxY9FCEXf7soSjyaTiXBF+YKb32QfMa8VIpAUndgMBO+3A6qf2Tj
MZAprfv2nJqFJxpO3vN1Y6ZikuzUT710QSuDeVFsDWlZuSLTC3jNjPFYufm09s0LeG1VbOiIHt8/
HBiRFlm/oGGchgHCpHLG/Kdsu7ILcI+IOpwlnn1mGrozVDJofxWvcspuHtlttJl8sFpU/Sm6OOog
27TJ9wivFEw+7TOJ9UwxLrwQmhvkdHhKf3BjDFDKOV9CM2dLE06J9Wgo4VxqIOqEMY2orVUlGk12
TN8Yycqnh2tnetXyFyOLLEdAkZCz+VcwDs0CdVWY1BG3zD10brsNjO/Wago3NmJwgm8RcdU9ikhD
j949y3cgNDR+IWSVHEDtBoXfB1dK/1KFV51I0jpv7x3ndsCDTtj8cEE2AQptl2DHJoe6LZyDN5Ff
G9osjYJNS5b2kheXKn+nuOhISAWoTmYcY8Pd/YtyJ3Z+MBIiWEPtA0I+gS/C2gDzMmkKML4HuZ2v
G+E6DZdbIacdSFrFvhMBpGtWZQNncqC1LLsXluWEyr5RERekA8bFiYmXYUK49TklaZ8U06m33gNy
+tJNITWe3uF+b3dXbMOM/EQIyz9s9Ih819H07I4bfzScM/DvUR2MgVHD9d03/YCgpcfxJARMRPBN
QUR4+A9BjQYnW82KmHQKwuakX4ADnBG7NdiuauNwgXl2EWGyDJbGJ5ZJL54qbg/ic/i17/egVYaw
NU4boLoJCsc81L7eX3fmlWxLHoU/cfj/WfjyPCEZXWJFSc05tQCSrC8MJAzTlwUII26nD7cL04J5
J6rrUeEuO5PJdZnQtOFaPHTYPApVsyOBee66xNzDi8Sv9Z2YZSgHQ8bvdaJ+b3iKFYDuKS5+RLvW
lDApL1zGtW6+Qp6KhzDbtNxhrlI3Jh8z6ibSc9CAiF4cgCJxt/JQ85XZDRKnZ4jEUvWs8svaEtFt
zPwpsZTl2chHyvgttGAsZVNhjSGvBm+OEpcFAzhF7pw3MCi56MjmFGidxC9RcNkGxzkAxaH6/JtX
VgfsUsNQRWenk/FyWqSP1Jdv1vhVARj5QdivrwdgO9aUBKmbD48QpgsKoFD9NFawM1kf3PpILjoS
4AebyYVpad/e0HFwfsjjVDrHIXRAPkQYMFg76SNTHiVNuRF9++LXbV2F7AZ9TRcn+yqm/64zKNDQ
KbgiSCrjeYn4Mlmua/fIPmArthozwWPR3CJWbJPx3nNsThk+iQliD9kHOLJoa2mve6aVUoih9SaK
YC5XyWLXk1cuSSKknIX1Lc+yZ4Syyf/3Z/t6TAfQ9TMD6/QihcnL9GqgU7rgRuEno6N2PtIVKLSn
TUOdB7SFMQnKTbNKIQMNkr36HGAzsTY04vBBcqM6Gn5p2NVy7X6RXUgzRn7cTy2BExepmapmgmy6
CNGvds/P7iLL1ny1Kakatn0/E+G43vAx9GQ55voOuxU8XNsQovaRUwEY+NAnvAuxg3oBR46k1m8a
8jY5YeMaGkrb0oaV8gUqxm4m+0W2uPOFWIs5udmKxqi8e+AedIyvHHmBXZAykOwW7w6eLYcq05lp
+AXNkjkcbe9AdreYi4STApZvEazVHCiVgmU3leaCs/l8fchQ3F+pA93Q3fgbLLjUN/rFy9SDLMxN
txiDaYJJUFnlZASWoMHpZtvaPtiaD6eWSeyKhY3wJz0XtHcoTI8T1HX1SNdM4x956qRQFcG9kl/2
ypC2CI/IPjtgglspudRxy9V3y8gkw4mQZb24j4FsSaes+9hT7z+yOGC2hLShVPa8gpUE5TdKm5SN
naljjVQLV3J3+qDe06v1Ztr57bxoB+PYz4C/aZohPfV0/u0lYgCANwLqg2gmggEQ5zE61UCcf7GJ
OQ5LpZp74LBYZBO7KsXpKfqqYdFdwbTY7+vCi5YFhkM+Sy/ppABoC81y5ucg8zJ5KjQxH4dIrNGc
1DHQIS7g8/rc9gtt3ozP+Id6aqJCNj1e5SPgaLVWhpSTKrGUKLquZYxlVP5+lPWvdglnB31vJfGv
5Klzg+O420WqjMYRrwZamOhQ1/LFJUeIfT2zKsH7ABRVJMnem62omUup1Of5NlxpfVX9Voj3sWCR
WhCO7oipJfYZeVg87YJJXtzzELSSLJFMJuhRh/lIOUg6WeOVaaXSW9hMFIIoNfP4whIKL6bRTeM1
7LJNkxB82HfojoR3QoyA4cSAfW1i8hXU5DBL1Un3BMPDCcR/f+ydvtD6OC0LBwjitnNuJQXuu6sq
eXsakOYKl4KHzQheHoo62rmZ/uSIaOCO+oqcWjCV2EgPYLY2GRDLYlZoIBv/X/TBt5J/Kb90n1IQ
m0h/TV2fIGCIHG5pD0fYUo5BO7ctlw7H+yX7PWnYuhVYkdEqx5bDuF0tFDb9qYrkyObxH8AcguVQ
dr9J/iriTvTLJ5//1XFxUpeiY9bPyq1ehaDJ/sMrltcQIt71b2U5bdkEopSn+M/QYRN7n4M40Tzh
4MJZDC3+c7J/3bMTt66aCamqwtIeRLhzVqUU/mWzHif3OYMbL4S1+tzcQRq1Imb8z1EDDnFEji9r
8Mx12dcNaN+uRDi3jWSayI0i014IuN9kpGjPss1X0eWl5gqj35vlKKIE/6g5vJDS67qH0f0pgV1z
nHZYkagxuH6tsLKDgL5hJP+2LV64GOA/Yr8Cg9gn1WJExz65SlYZCnlgf8TlE1FUqpXc1iu8Tlv2
/KYH3/6HI0Ecj8Q2uPgtp6pF7Pm8fsqZ7rEO54f8/ea5ZGWXALxDF2grG1J/53apEXCIGtxmamUF
MDXcv5sssYZhshueL/cIxXeu/u4FtRzERvSYFNogsG4Yy9CJ+n1emyWqBW78V61SVGsRnvTjDQe/
iEECKbildXvMOWWeRL5bUOV6x+fxIYZHs2/Bh8IdcEWyA7G+rQDYOq3jykgMn7oc4R9fIRD5sgI7
LyVS3Wvt8NPy31GYHVDhHin87D/hyKaKPAkHNYIsiXPshlRHePjJfWwbJxp+ZLPAFWZI9yX21aBl
5Jncye2ZOvzeajbbDaFDZ6QKGYOnXLxEwnMtQHZhgUYheEQFCRHWMK70JHpWyLMB7ezou2iyUsXX
ze0peSPr90NeXVG3mD1vv7XcztUCy0ZlwHAOtow4c0azV4/rrLrCQpFuOKVijoxcF2/MN3+f+7q8
LEa8mbCsXucFgsdhWvQXMW6GaZcbxvoFe4RT4Yla6aJuPqBeMRCKUOfqpdhVaaQqdz9+sAl3lpEr
wIQBSN4P/kMCOoNRXxcgihgexNIe5IMIFdKdWim+wsi2HImcJE6jLtpXyOx8kjsdrpPLE2w97QWD
doe7YvGMmAUkNeaWH4mXRD/Ypel8HhO4aA5+4i/eGIZaF2FBtfQCLqmG0cbrTNhSCcR1zyOb0xKt
GmbqqQU/ryhL860th0My+OEqlqH/uGu60hNL7RtM0JzDUHi6JWyv4XAiD9EUhJCiGMqK24djV+Xi
mJcu9NZzGPL/ilPvX5f+gmhCdKawc4Ms+SwFgG67IJepvbnwRURU4Hl9tDEqkwpSC8i2sppr/MwW
fI1qyE9t+nCyUJdbo3e6QaLpjnIhAYj6lcnmPdfE2sIeoDM9E2b/84KZNynGIS/ao9BqlwKbpevT
f9VuPCixtwpn/I1zfPYj1J7t3MBFL88HpzxF0tsPrKyxqGM5hZvaE+zGizdFDH/6aGtScyy40VND
yvex/I7ZQrVd39svwT5m1cGv7O+0vdDvOI6Dnzt24k0GW4MS97kcA7CKACzqn6sh5vS6Ua3xIZ16
oyWQJ5A/pzaJ6YsSK3VdJk9kfrfM636fAsXat0qjcYF5vmQwCEHBxjrpKBc5jZ3uirjPEYABYPMn
TqMoZc6Vdhf200Dzzk0W20gAQA/QiT6Za2PO6ZJSSMMyMct4zkLGB768aVHvciYvASxa3YTi1iKm
Kb+IbiiHXb40776Q+pk0ut162nY/2tl0cJ+tYIF/V6n7QuRMCNEltw16gXN8SnXuWoMfWb5ReU1P
YI5Yjes4rQFsMXyQsm5XhhP2fubNse0suSl0wurIk0ztkTLMLB2LJjbYdqK7OnIC0JXD9FFnfjAN
qnvsCDMhev85E2eQXJEppr9U3DBoT5AHDOkOgam+x4L2UoS1UWnRyH+FWV/onxyog7WqBnwwVWbE
ZgjqLFemhHIAbhuVnHf6mSi3MsbDqqVLfeSAfJgsZdjPSMDMxlvb1h3QijJ2oF2ZxZEQXY/9uz9E
Wo6zyqZriBfFH3vO6WjNu2QPGWY71MEQ8AbqY2oJei1xSCn3Ka76hWxxCCWaiqfLm1b8j8qGzule
wLz3Gqz4Kguw5ngAP+IwQUj6UoLZGjuaVyqQoAxyVRWGHiqY9CjH82d8xQFQ0Uwzj4T/PP6W0oZS
gM6krmn4WyQxkhD88LJzUjWV3Ap9kkCkrOnYJojqG9QZqw6XDgiXchoQ1Or8WDjwB2nDIDhmFkhj
BIAFBbkgL/uRApf/IwHC/aPGafXf/vUErjjJMX7FiLDvpWyIfaq1yM9PQ+xGHzxKCl7Nx0G5Z7ah
4WKhYBASj/Vqjd4zx08z1fRwoaRJae+nHndsz5DEzAPOoEmkTSbs//xdDtnlxU19+f2kOoq6JZYo
n4Tc5rZ0TNJTpSYZk/sVfYtUMkJXlMkQE7nlbq+Yxd/eKfhrFFmafG5Qq0UCiKe0dAbop/qRte2g
DK+usfHsYJKfxOf5baCeA5KHHWffFeERbz2Bg21DX2AlD+e//kDf+LoazMzTHsYsddvKcxgOkNky
NQ+IDgNysWPYG5pyDySfljvIMZCRV5npntjYWiPPHPEFO1Zw2VDYwSvUUJlGxC+3CcwspZkt05LL
/tg38DnYcHWmA63oTQtSai9f4giNDO1bDNyvId1CRx7/ScHhtXDVMcJdXMdLlkyJdyacA1XYrDsF
TIsUOlwsEhVUvY/yb++8nMEIbAYOYa4e5zeW0e89WXPFie3iOcyeMFvGJ3IsNRulrxvEtWgSlT53
6HGrCuRkG00GbAwGdWKu5ygqnZDb1jxXTfFPxvllNTvIMxcx0NmdDCPDMKbY57G+whRGxiloGdQz
ZL4v5C2WkdOtenkflB5fzAyaIvICaEhAFsYjLrDFEcg7LLOGQ/ovqix1nba+IQ/iAMdk+94zdV0B
oTUHWqm6f9MLX2rA2ZPf42tBimfrUMQ5E+gVvhbLU4NOgA8y8u04KAdyyUqKHvOHrMjIu1fjwqxb
DvYUU0Ix8c2AckYSYMWEo0T0AmgpAdZOFdymSrLPI8ODlowbnm6Q5c6FrTrvi2gETHEMBs3KJGBc
fUPhoykaFTC9H/HXHbz4yc/QQvciv9ZDZEKppBo5v54TCeJ+wMLW90uTRrmheAcGQq/q7+ZjRZWG
0Q1Ry+P33It0KDJeDnJP+G+my7ctUEa7Qx3mOIbMHtgoO85cqGi0scOcxGf4ATR5pgpdYkqHZVMj
rVykr3+2thy9aU6AqREVgotYyX+IZCq1UhYsDKvIfMMiMcJT/wUXH6uAX08YRIdcA6aLhOfl6r31
wL2bdVoku0snBng/wEIfcynbRglcunqKBXJip6cNHfepRFGqd5MV8grnRTJYLY+L8knhFoD3sBwp
yuU4Th1F0lUxJz5eI4EjH9uLZKvqyLTV/JBuXBq5zCB8FroYHJRmuMAdQk5QNZn3hmJkLIrTGdLG
N+5rEv+QJMDvj4ZzVfVHyygASl3hWwN5qm3T+oevohVYn0tgO5MujDNyZtxpkL1v3fpz5re1ofrY
0WaoLEvBXzRESTTotB1X2QSFWqqZ7hx/jC9zAukgiXziDZ1g3+/X7wAmWVx9rOPDROtwJVNE2aDN
1GwO5IkbnX2KciqeTMfn0v5oKmiq8I72+BGxdXDpjjOWCXzMu36DObOx7iuB1iR+Au4yG7nWqyii
oWQfHIVDnjgJA6x/mAWc9bxgEBacNllcxcJ6r/p9sSmNBVhbX0W6loOupI39RZYSKrnOUJlSHm/C
hln2nM1DsE7rLJvftgr6oRxXgCrRCpOtxvy9s8zZxeMBL+XD2Q4j9aAhfLnbUCEeNCgxc5ub6JO0
Pbgb5wsHxdi/yiJqst4aIZZmQSticL7Hdby0UVOIDV1vv+OFK2qd2JQc3Cw2jj7FXHVqBhPQFimY
cTbRiYJtvNF9jwRMnTGjjMvO3Qxo4CU8xKPwGqDKukNY0SSytb58m8FZTqnwumSsEbGPwaAC1Tbm
CZbB7xGM85W2gntjyzZwXQljsj5u22YdXD6n6LnGvwcjuzL9yALG2xSVGniETeyWM4UMMjI7qycM
puE/XOmxuIOOg4b+FAd5hQFJ6n/z1TrfyCI6iaGyxMH+3adtXDjRuHckjmeWrb3tJCQ5XYX7xIzp
jm0zcoAvGVfWSpPl5zDY2fwU/qqq02PwMJqev7IJ7PtbCKTbhappbrs2EPiBu9JjCXpKy8TXNenb
yQ8UbG0mx1t545PgKsTYqgzH9jvr/2WUBpJe8cucfn1G/MdylduIZxQRhqKtQ8VAy/QxaWvOkXsx
3RU26xMGpa9bGQ+Vd9a+7TiHmEiRK0JAaHiGvECfVGc5CcwSNFVOLPzlYgc9ioulhfDfSKGJU8a0
o5s14tW4MoLLL/gA1rPSQ3kgzPX+ykkmJUayqR+DKg49X+CyFe4/1iFz3uEazMRAdFbumI+NeN2Q
Q10hfDCmBf+IbilSHkqIQb1geEaRKMC5KY0w6+g+Yy+6vKdFpMVuuf/OY7lOZCfp7Y1vWIwI+cKI
foqcXzHvSCCcg6WAB1rqLETw25yLo6emV2xAsewQDKUfMiNoZ7ek8KDjfqnIArOAQ5tQvzcSp+TE
UiNA7/19mabCG4Ty79kO0yHlzkaccbyojBm+k8fQtTJkYZ7FscpEA+wcViCGosPdbkoosneO0xKe
oevIfv7Oy+uomdxcqaU7ME5dkA9PslM5l6ul9JdJfyPj9UjbpgZUGoYU+rPiaoQg0t8Plp+ropgU
fhI84CKMUTExPpVUCEjGCGItro+uUlQvBZhR7zIhL69vcEyaz3L7tGyS1k3O7eoBQ4yCmr4X/HYS
+Eet7h6qefAv0BTp7bcFcohIBNm7EUcPv8+Q8+maZU7dHWwtzG+bjypwIPfWXEkx5YjU+B94KF0j
TZDAZFA/nNIwLQWujHYkdWF95ezjuYeyz7Mn/8jK5Gy5ak49gixWFK3E6AXzW6v3VY7ec7gJLl8R
WOSwhLMGkmc8rjR2f0ZOmx3ccNbxZ6uNmFgeBt5t95cavaM/9fFdD72tBw3vJqqz9Lj5erG1pH7r
CSsjvstlTBcA33Bu6y6O+9oTkV5bTodbTIt0Q5lZAfYyUZVUStTWoNqjiaUHoTXb1v/cKJJ2UNj5
T0dwYX0MjEUpggcWmP2rnXSLpD5Y5ClkjmW2iBfCaeUf1gV2tfp5l4uj7TI2oT0ZHSA8B+0/dzHR
lWsn1pzDZnNtBTJV/e15w1213Q/JhhuAEgDF2P9PYn8+7DKJjOo824xHqKryvIHHxz4lVDdsk6TS
DKIT8XzTb7+8hEBNnKdu2TeeYQJE6+WZDy3KMFQBAiiw6XCo0gl1EAnidgAYbJmNcjSPGDs8h/us
GKbJ2PZpSbvn6hvMMfNh6mbGOQmqWXIyH1Uco8sYOMgkYUJQpvtG3pe28htQcULU+X2PzVogZp9i
w6PCHQFenBao5sBgyg8FuY4RFWVk58VhgMA/7X4EB7rLAkWKP4Y2edFbCDW+r6Y6xUTd8zVYqO/g
hbaSNv07qkpccVt7VQIiyDjBVPTgUtlmdcL7kFFk2o7iYgwFG6Pvhzg73QJBZBzaWaXhapEg61SO
PzqaP0w/LfKYQKPYdhSENjfahNAzIT3U9yCbiroM48CXOtR3kRcAy9mAfKHewOkhrzq6BUzXejqj
3oM4ttGRDzNq/Di6J4+syPEUETBhXqybhxFyU+VPgHllm89/R1Pdn1C0Wbptz9TV6koIRXizcmWe
IbPUft31w0PXLyzbxleAXH7DYVt8gyrnZrVPmZ07RnOnea+4MGbalv5+W9ek7bpyhVNDnJ6fuqGE
WoTw+nWOz+v6nlwQek6yXyLKNWp/4j0X06kfuNWj6+rWX3/cdszaUkMSOvFtvclzqtWk+ITJowI7
iNdolef9zmPgZutfyewDHtVaGXTDJn2yz7YyXx0AdE6PQGfakYfk2YS7bBP3vQDHDEeLW3LzG10s
IlotazBJs5Ybbd1HGzr3+KguskSHJByScdJJQPlyTljFmCcyRpBrPjF/k6fi1KYw15J7zZd/EoDO
RWh1HSqkXSwORDSYW1jmPtNJDUwTzHLxFDZodjfNhgTmJ/irbhBmEhSJhrfjQ3i7hH7EbciPWZjC
sl+eiTLizIUz8V7tkPfAV5fjkI72Z/r4YVt139yc6ks5YlzIkcKxg2J1dTFzO9v1I0JE2Yl+Gzgy
vnTPvo74tY/Ff3e+eGF2GnJryNNRfckZc1MtvwWSlxGiplLUI7oXPQUJ2iUTu/aMyYBuHXvTtiol
2oon4c+k1cxfXpeqH8ckCT7wnGeXVfl6PXAGG/HCWHS2N7I8Cjf6vAwyF9vZUoopDCAqe+90Tjb1
9OIYEpm4ijkBe+zm+LPivppNjf8fBJxu0KGQSSScFtuzqavjrQxDJG6x/NRxe+xt3vKvJx+iv8mz
di8/EnQBub6fvttcbmxhSbnTcuaeUHD/vWxnf58o375C7ljKucH0QYhtdBTxx8id7ShUScbPDYPn
L/rhv+SneocN+HdSAmHzYlWYs21QU4+uG565r27t383KFZO5n3IzpNL5MBVlGSwT5lqKVqOJJrUQ
Oiwit5o3mq5Gh4jvVq809JICBpCt64OVWrN1m3FX3EyMlodYkNVrB5sKW8qghV4om9LJJ+KR/ay0
XK4+zLi1/lDk1V0qOWgIyICGwR9G3NTVGl20rdYIwhdCCVDHiYAseGqKwdl9b09qLVA8m1mkwigO
N85Ih8+Rja3+RoV+4fum4KcO9FcNqARX3OcXpWlm4nh35NT1wnDQ44Xi3UfXTXEAntuEOAk+OuiS
MPn0827cIuh7JpiRYiLpB83VrNXG3g+v1G+qcwp6Ml85UuZo/LT4GJuIzyVUDEk1NBaPPPpMpGvD
K40qRqXnRZ9gMBFYhGkqdvBAY7wgTUk81WBR0ZPDJD/yjOO8mSHGRdIEBrIUDk/GwQul0Ez0ywz+
jtwlzkSQaoDxKoe+oFkOA3I4QMT3myUyXYo7kLFIx+mlBm2LB+y1LR1N6RETCat6PtBZmtQTixL8
+sBOYeLTZvP/LMZDL2fOOrmpmcQMVNVFqnDWkd3J/R47RHP5lnSM6BnJPVDDOFZiLLQtXpoGIHjl
jZTCMwRmIoBuI09H7auy0PStbIAGjuK0YfwnzCVZNiiBYmqU6jTmIhspsDLxUIz97XjLClEofDwJ
kYTaITkDLCLN/rcTPqc2zTjWAa69ekySQ05Uc5wIQ19Dgvdf7Zh7ekwu8qPlZXjCxpUcZV6wHugU
96IbyNe1quKnENDGkR1umyobAEU/QYU7uozG4CGTCWU8H3eW3vA9AU98M2WpJWui5TAohFOaReug
UTIwTnBqtF41lRRyyqREY+OryL4Yb4OKc1CdH8esnOsKi337ggXQw/3Xovio+945T3H7SU6BGhfY
dWY1oqzKxlX8kOTwYfhPapXOBfOqYfBTel4666mLAxneRR0QFhcb+5V5kzNtWh5D4LYIEWnks5Qk
sPC4AWP6FGGnzWaSj20eKBJ0KEyjlkRUtZ9h8QsqpEUQY6js0dHL6jF0bYFKWHSomkWlzwTuw3vY
mNay1TnZfejKMIfapS6IBF2C2QQcuEuniJ4PkUHLwQ2UQ+j2gIWxIMv2xWaHOomUNfylhyHlwLvC
NwZmwL/UDic0vSPjMfxe82Efx/gC6qWN16l746jTPxjMfTIu08ve6tVYSUBN5geLdYnPD7PcpWJZ
UrAGSU7oR7byXZkhb0O6wVABKX65+V52L2xFGd4v40Qjb0vPVn5/AgAm3Qxr0agwQEKksC/tvHeX
YV6kbbdcpUxTGX1OfE95qAR8mAPdehWlmGdpvBwIKuC4xXaV2AE3uEntTSHPteVB65QPFmPli4hc
NiZVsUZ05MwmAVsOB1cieYb1rS/PoHyO/PdWqQwi+N1mm2GNbCef08G2KoRbNwKikoZGuU6Nwogo
byLhxGTF+mySudzHO9dFq0KO+xTaZifcy1flR6N8J9rviB4foqMvifyywGt8fzeB5jXrSted+wDd
3LL3RAUFymRWvTyvOKSLjvMj1fcpi9HljANZOrH3TcYlSiPxSYS2MyWqCf54tAEi6f9SRbK3aqMS
BFXjwY8voruDhCjqbomF+6cc69WS4EL58vpSRBeMKJ5L32C4Fus7HZ1WSMekhxqhpIBO0BcBdeLK
LBDAyHK2VmYiu8r681HofLwn2dl7F3zaZ8DPJtdOsAMjTpEQB3x+AemcxNYV7L+Xs0HKO6CPiznZ
iADB7qhDQVgZ2NSmHVS9Vw+mfhfPQH6vWH1SccsCMfdmQkqu1+RIui8znOAinQTYL+VfjVoAJlf/
SDBwaRylQhnekLkmNakZrxRPOg3xHmtjiTE5MVOij6be4prUbIbKlIxXO6lpj1qX1hwjGv2g6seX
d9lcrc1aFefW6ELGMabnXa+5TbHLYGp8bKb6CC0M/scAKQSS5Nxp9dS5M+9Dzz0RICPYmzbS5H7b
tmaR7m7eszR2VUPlbOaoh7EzVBJoJxiR/2xnjwiKjc0u1b7uFF6lH3tolX5JcXQLcFrluDpV60Nl
kARcAEZq4ZDaE+ad6RQGzFMDReRSCThXYVsDTct6hDz0DWP1GMyC02oXjuo4QV721DrWDmi2277+
Twg8zRMMtRUWvI3tQu2ImJFh40LgWfitwHZ4gltpgDxqguZePy+RMzBhqUIRLuyB9GU6E35Rg9i/
xdzGgP8ELMdd/GsTZ8+HQbSrQgQE8IrqRl1wjgPkkcr+EdEkEa6f79tgYK2Wc/hoCvDGZsmF5N3D
LDRFstTZXd2fLhPtxkloe8HcVTWiHo/tRJZ2UK5ZhwkvXxGLyXcnR6x8cL2DzkhN1Vx1DmthXmEG
YeNcNFxAd66KGTW6udGIyplO6qNT6Hpbde5rI8414UDizU5J6l32ozcVIX+pEUczr2wG91ynxr4L
Fzen68wrEWnGCGgEvRbex+k2R67EVOK0RRaC23NP//pglRdcdRMRpwQeu0jSJH/nE1iekXXDQuQP
CRCPbmtRmgamiI2SYh/h5c2f5rRLLPH/d7zgl+rYCZMvGZfOEI1xpougXsKKo6UQLE6G3cke72yu
Rwd2OV+1d3IPaqyWjeKVBbbDGHV1IJjm7rf/2KlgVml3VJW74QeKkPdd+pIN3eDKzQUJ/a7J+OR9
WDH+qDmwJBU4RxrY5nw3I+ikKxuwadY0koVb5O56BIMX9zb2Npy54YsuDgj9PFQhprIB1wlsTCOT
Uy0R4C9HdwST438IeQaIvPQXCgpQRYbv5lPezasJdbOt0EtaJwa1f3kkViUSH3a2OXdCUy/epxwL
VkyiSJ34vrCF5L6GRiyYBbp/+sR2Joo5DG4bmd0+tIS/L1ZetyLnKCuJJWIkLNtgA+RKqDkQgSqp
vJrUHfo0Q9jRLBAVe3nZEx5/Xg3k0rJEPve6vTwhn+3d6NUOLmzyGg83I6fTdcJLpu8iUGusEUM2
VGkyx1YF61Gqcej5i25pg2f9UlRgk0s37gh7fPz5/Ew82zJmx+PJjLH6cZ3CFjzUX0u9nEsxT8nI
pyipLLPjcDK8b91+pv0LdhBmlDKjTqmi0pYa66wyXB3nEFK6EY38BnKp3h8iS6dh9D4LPbAvVSs5
UCYxtq38sPvFFEoDNldhr8LRTCNEA/YoeimMXB61zOB9ASWQyLrVg+w9PMWSeESHrfVz4DOcy0W8
2ZAssfuP7X6YOCpCZBfdFiu1xu8oInQIZwgwKUavqZRA4WRo6ylv+G2wfYcVuthdxV0ZHOWwpY/w
ji1DXiiUnOvmIEa5q7eKiIC0ZRVBm8GQhosfVO3GaNo3BasoJRlHaOU1EY1lmgwuufPaszKQ7FSZ
+FPETNSQee3MZy8aAiMKX2ZK1/Fk7UpXJ/bGq924EDQdaaISXLJ/pvyu09+B9nAXtscuYfOS/aly
Hvc9zMJ+62raM4yU+ku7WmOirxPyv7ZUZyTfEePkR7GkuEs4ItO3NW8eyKccqHykKyNMuJ0oGb9e
oWU8MuebFl9vxhacbfySDrxlCgOaZjrqW9NtS5O1WfLNKZ33Q6jsjQwRirTzp453RhqMnIU/fUZO
Jx8heVc7bUkCWzKPWmXN+nPXGsPHrG9H0ks1clQmMX388K+z5D9gB0sF/EkbJEyLzajxyTfBUBps
3+Euq6Ooi/M0SAXu4nUwvW/kKYHNZQErkzq+Q1VOf/NT0wVI6DJThHRmjQ9xUqe4OhBDAtEvINwX
9z1yNCjjZZZ/80T9dyPbiMo8HXtdRB+q6EdDPiM6ASVgBtJm7FPQwkmCjy2RWr4A1J8TFIOdaqzq
nvpVFEQtZayc+VVWWC9+kffTZjDdDIjT58MbeDia6eXyhgWxn+lNSA5NVvHj0Xh8Sq3UbfxHhBRf
OgBfVGLTp4+TKH9dwV8SUvlvD6sOJg0ZPhnqMWT++LDS0Ai2fz00sT0PT/Nude6XAwn5y3FC6fCr
Q2mdS9lm7DH9JLKnQcCaExxW8RNDnN54z4twqVU6wzRDPa2hTFOM3Ivtijwj18jwfXCxFjstbP/r
5gQ9zglddawvN1y0vWNvUEDrAMTyTOfad7ywGveInexT1tAzw7jjGVkrWjgf+hTeMGJsyofXYVFk
IMi8A+3vegQSJAPaHfhdU4Bt9L+uw38Tm6+gx84XRX0X/LqhBaTw0sO1PS4VgkuDdoNa0oM3YGL9
QBgf3tpCunoqrKKCmjrju+E73zccNgdQMHUerXyk9ovH3jVPeIB14p1lV9gd9mJLeMiy4rVMr3Q5
Hyq8BzUT2CwljX+SGVJZeltlXfABh+kehYkzHdtpWKk1qOXRmw68V6EQz4idBAUt1BKo/C+epvmx
I3AZ9Bv5v+7JF4PWXgRKTMNhjN9dN2foatEGrVfx7/2f8jxTzJ8tB6FQlb0leCOSEkcqZohJfw8F
KJLRahpAJpInOuqhQYDhWmh2sg4gaSItacV3Q/ZRMZqBtAoIGfm/0bRbjP6KLukks7ENtU/ST9B/
xDZ6qWsrvfUaqc/TBCb4GcDo4TN95kWP9wYOUtjFxYa9IQ4oIwWCd8WKjgaOrG3OX/F7N/rVBnsb
WKDOW3Imoiq41HZ+zgCrb4Ks5Z3wEhotmxnqlkeTL5DuHuRF8NoNKj+KqFijLC/TuoHCZ3o+LWI4
H4H1Kn4sbnQtpJ1cxM0Er4IUlo2tfppfWf9UwhsE7wEPmHvimzHtBRjnw4cxl93a7VWzRC1DPT3O
yKEcrvkdTXP2LyRw693Gs+Fua+ZEGqIws0+0/Lh91Td+b58Uz+Qn0s3BYNO19fcRVZoZqIRAjZRd
xm6DaeB2CMcWnItpx5sQhxNrNlz1SLMSlPRcPlfRgAg9PFz+NK2qXONumHvUfgL0PaUcu1+xoj95
+0g+Jx8mbrnt45ASFlkYPWgih0glDWRIi8Uw/9YqeLWqjjKU6qQrLyWQ2s96gD6x+wAkHhffpsKd
PF4D4yoYoBM0ftWnG2CPBMwCrYkTscB4wamzW3JJl3hZDEMGfUmhwvqWKYbDRH62zzaSJT1oEHAr
E7yQ2uGqrq5CweStK/+CRmJqr6MhAV32ws7KgmkRDAMl6DXmrQoe3Ya7Z/Y1vO1m7M9s0+MD3xFe
U6qYyI6wY9gWykBqXgtG+DwXtyk1HwNpFLmpLAyLaAfZ4SVRB2sfvMOYZqEHsU4/JqeM2dOQy+Jb
LEmurdIHoc9fw17T0swutvp2SvcLvyruUoqsDu/QR1xAEpcge1sMDywBU0HSehg0xRzWOlAOb/70
Ux7A6jf/jc4fdlrWAZtgmMhhrG2GACSlpx62xwqx9SSBKvg6PxQknCYEpSKI/zYe0BnLeUYUWv3o
xyOxPWX4L1CpkhEjYus0DEzF2a9ul22f7GCXVGnz8CsjvU2MZ0S0Y6XTo4Sx9nKSEexEBePneybd
NW1+mLOqhe75mlBHmbPWLOr5udy+vb2zvELikEYCSzBqbiybmxK1dRsokjYNSH2ibinjIiJaJYVF
DXU2IuhDzySEC4V2YbA08GGrEVocgUHVIaZu1Cd+aDZai3TcmTKM4xpivBrLLJ71sPHIqKuKm518
bofY3ivZ/6qKKayOZjRhOgZAmkJT0iz7QzbWP2RhHNmYH030REu5+BN/8yWGwVeb+u0IxVBat7yV
aWwKeyVycqYuqhBg15xaIyIbtAWMdXarwRaFrX5cuFGVeJ+YTQcicttJ6mT+zLOuIN/E2OV65/sy
0iCQSqZHcAaTlmrmZw3qC5cnu4u3RfQhFPdhFUaXT7RFxfMUozWXd6UZjqSpyX1gKMR4ae1lh/KF
PgXDDQQt0jDV0PZ2ucBqhPZOxLzmdIPEkyvAVonMHJb6IDXOyVp5RoLDRep4H/S2ohtwIGXxLNEe
b/gD4DQh5IwI/LBxrKznm9yJYi/D6mt1L3h6g4iA0lbiI/Y/CDtj3HRf3yM2IvpW5tw7gki8tV5+
PFhW3fn6OF7KnvDhAYWLNYxeK9AzU+YrdhkDtPpk4UZSPYEKv8gBAbGgv8vjbzrrC7ZcZYvqPW//
FJOh/8P4aNDOHBxeaXCZQonfo1zWdjK4k9LJS6/dx57UxTmkyX5JFPP+5frX8/l2y0bc1ur8kqYA
FieQ4LP1E5wosgmTnbw3DxiuY6u8XM24q6JwqVq07AybUD1RN7msXlGyBJBfes4ke0DFj4Rea875
SdJL11VFLob5ssw8wwJGmBsmJFtbsXoPgi6JJDs+5J1EuDLG8iEbLCOfIbvhz2UU1MI1Gz/Vgrty
QbWkTjAmrMDemqCC85pB5zNOMs3jmFyRtwVe/ca0S4T9F3qiBRZp5d45ZbU8ZfJ53uJUCdDY0Q0s
yS8xdRjIyefrHaWiEUqkptGCOo3bx/zF1IpJYqGGFwT1PMvWCr8IoP3Jd9HcfIRkcUhABYq9JHf8
QvSpAVqgV2Vi/6DzQACuHH8QzYwl3jVba7u55hwleAvrLYGlBgm86l75IEJ7rHhDmDnGgT9atQDQ
vrf5uXBfZMqrYTbZr0keoL0R2AXaFQtWcOF1CwVa3UscV47xydw1uN0ul5yX8Ra5/LizCcBX2dDd
yJa122p2osf5Ay3MfPP2bwpr2p2xTvD/U5cxA6+lUbU7e0KA4P0R6DADONJoYgGZjgfHj9NL4uhT
lTWzCJt7pIte8gn/BfXM0r5eBrKbMog0saHN2oxID3TlRLANffwTzhsdN0FIje91Ty9ue1zajE6X
hn84ywlwnYcscxnlkVNmPweembbHpmBkMBhcKUpr/YbuAgOS5H1rro3XkCtxgN1GrYkFVidpCM/f
50b6YTdc8VmvJXjrePi+9tGkzu9F8oFva3jBmKsx9vuaIokATQ8p6QW3IvquiJ6/apWSRs3jqz1x
xyXs0dye31JrOM/s9qlyPIkJFuYOuUcsFf9aZsVLBK3ICvJY1tvWKO6aiQjMBGAGLZE07xEjASpJ
lDI5MxK6Fl5l9h4un7qftVgSX8uLByOY1r3VAHhkTnyKYtueDWzAnJ70TY0gDZhIRB+10slNeFG+
PTf3ydeOaUuUsdMbOa285Hgs1caopZj6CHEzdg7duxDfLyUxYzWBOf0TRzkIAqam8aEv7PeI8Ccn
0EUBHBGaEy1A8vqFhQydLGIQrkHJX4PeXrygdS/DLlNYkkCC6rZrpZjJue+a3wgMaWLGnjMuyD7m
xRY+F3bUL5jXqtYhbNd+WWIzBWnnWCeYSfqhMwDK7G16i2eQs2h9qKuC/cYiChvnX6JMLH+6Q08Y
a7R7daO4m8eTeQyz1ngZmz4HKLMT+OKl3Oa9bwnoznz9MlUop3c5FNCqbTVZ7o9jI2FWB3MJX6AE
KaGEo+S1wvsIcsbsoIDCVagVJN4gF+VRz7LtVfaVQhdSmLwhSZiZfdQV1ar+jSwOrVeds9QiYOWq
gfJGkrMhenad0FBBnwe0oM2+aOJIOzMhntgnJJpUgfxmNQUP4M98Y+0m1FtL2iYl3DRAzfTrg/Xt
BZVc+jjNDBl+YQT+pE7kOu/OvI/84JrBZWQ+cQZovSSde/rL2vP1z/319SHjhga9oJ0GWDUqvCX+
f3ekc+RPTn55RjOdU7q00B0OddXFFL/j8ZsIaWJW7XYbNJCc1xPqFkIZAeMVao5ElL2PknN4HRnF
mQVWZS6yxJn3OjrowSJvKq0HOxTdGaIYA4Ke01XJ7sknSBiZ0CyhMRhGD33TdtdzR5V97i7e3BXD
vEjP8ODT6/LzWRDfuwcmcksNq2jkMQGG8Pu/DahYureYmpapskU8DnxoXHf/qiHJDHrlsRyknb9i
RURoBmjk9mk0BX02s6vpgzRPHdo0lCNgro1FjthowYA6467rD6g5TD0YQR2VN/nUrh7TJAX34RGj
G1HpGFSQW7Dtve+NYIKp3WzNfrL5Xg5Ny6I1cYxdD3+7Q4kRpGIB/UHEtQiGyPsK8LbmjqPpDajb
eEgslmp8BCWfDFoQfR1DIFlW6gE7VxkoJ1V4je7KbZ7HKYssrXmzg3Vepe2PsO1hQOqt0Ax9JCrZ
EvqTa7/eK+IllC9y6XbO7f5c8R2il07zpTnifBLvtG96QV2FCtRXtDHPcYYivgWpYWnCG7XklM4j
d8l+1U+PN6DK0nBVYi9tZONOh8r2IQJAHYQHSR7LPZFTT/Cxugouoyk0cYgvg4NIVAQIvfEAHgiY
4ElG9UXWY9ZbxMdbO2NhN0zzRb3X9CFBUpafcYpD86bopcBp+o1wKnOmLPhXRQ8/6DogpnYhD68/
ErryWiz/sE2cFx9qTro8gxz0xSdogurf0uIkEHaXZGFZkR3lY8JOTzdKQA4RlZ2IjHjvCaKasSta
KAKdJ3OjCad10sj+h3rwtDbk1qBFUfp8Zh80yf0wkdy44tFUidtC8kEGeWb6WS6YO+/+/54R3JND
gq066+BqA5qhbY7uDt/RCNaZPEST7dLbAVVUsomdKhC4UZRkw76FieV22g+FjPry7E2/H9LwQ8Ox
l0HoNB2Id8mKGXeL5D5RnKi/KakYljlDqrZLHSFfMIYWG5kLiLkCmEX/QgZktelbfRW2ClHj8SpA
HXNfhsHnCap6e+QUO6C5sb5uWSkQcII3PfSbc1t95f+Dul6btf5lelC6qqFz41bX0fwtLNZ+9uAu
l8pdffo+lvqXXCH+QERROF2GtPQOBP5qHgobzOQKJcPEkHGSSTncHilYIIMKgqU21TuHOweGRzPY
SySDBAwsU8bGqhXoOgiF89Iu/dfYqLNwSdWvOGboFUHEajcpw4Fq0WE3qDCKAMhpTe0/9sN/WKSb
Xkubk3fLDzp+QWph2PojXgU8B7mbGBaf/FoBx8BaUkymA6H5tc8HrNif/usGAqXKmhYJibrZc4Dj
FazWzia39egOjNCx9/zjZ6lQ2nqLN1htdCTMHCVDci+AnmeFHeS/aBAPObLJSw2LF3V+RqdS9ZDe
ncD/08ZyC+rF41/Lh3Ge6q2QrWeMfEy4AnFY1VwLE7IvuRUeFHPnGh8EJ71/JY31bcFvjiPsPCRh
qPRJ+ST/TPN9U77vRDT0Uq6td1siGfmB8ofPW73ZC47TFFh37QOXMIuxn+AqXC/LXATQCfPJ/d7y
H+gZjHOn0hPtyMfV/tV1mXxlp6OpiclVViwkUhqHvjfDbm3KN1nSBdTkokepJNPAXAcRTbr+q2Fr
3VaS1zxT3nJ11056yp2hERrCSPw7J1tGYzjnrx2Pd3Sl35c+NyjrdGmwF4krxGM+99QNhW2H9rdb
j3LHc5ygFK61tPLM/KKVNCo6LXVuILC6AL9DlW5OchgLbM7vNfsH+9APqDMf+myKxmInc68QBVDp
jw/Bbw3zxC6pXOtqRVJ1ByLQ/KyNTnPlYLpjc24/PAknHx6BSWmyWmK8i+rKaVR8G+9jSgkOo9EC
EoKKY2IFxGSJi1XnQs+5E6wWPGoRC/OgiZmLg/D7z81IwbPXtOo/aN/lUy7esiIdMgN0dgrIykCI
eb9ruyTVjnFBTQunYmlvk3Pbka6NCcWBgTlw5mAQi8zy3thvzr11ljTOWlau6U3eOQG+yWQsEN5a
EjJOwwnDHmBSMxjH3o/jAV/QhgA8g99ndavJ6MHcQnDZPherlFJELjl7G8xoJ46WZwRwUM7Eb/Cg
qi/RueGatHUIMKTOlQuXTCLlUwJ1kv0kjsOMCq/xiVAWS4EQJOY6RKvQZWzK8rfVPTjfdXwvXUe0
c+qu+77aNEMpf8Ogdu6ssjt548z+zoTt+E9fnFJSjb29/DgEqMe7NkO9HOMvcvIWws1OloVon6vm
aHLo5TBpXgzfNnTHJPf3kBsAkuEZw7Dh4vQqs8M44vIs+bbM47moyg8IqcmpateOadIuFSjQBeKN
thIZWFynHyhnE27ACctwcc4RCPHY3prl4luWcU6Y4/59/jL5AB0h1xb9DlqzsilNRyv5snhaXSo3
rkhKnN0MI5nR1ewFCOAPdTr8kUyheE6I0OMwrByoXj5TXoSWws/jS8GIfJJf/cg4DOkDKlevpjzJ
IAo3Wd0p7B672PEQyV1fyv8tOTiAX91FYJ48a6jNl56nf59+sx1tuZyNleCnqmAYCtJFkDm1Rrel
dux9hUCIgY6NrwBpoIsUkSFeYBcU0epwEHuwLnxwJlwApignfchJrfrveSnanm8jjOMj8rf2xrVx
vs1JDROBvMg1/cWd7NgC6hF+t9AzqqVYYWR8/OSx7+KQTuGj2ztQPQNPIwjb5rBeNLDcK1DnT+e3
4II0lw0xPqCUW4cJasn3W1Pcb4dazDUc1oMbaLAHUQn9hAfugjFxAyTLI0jwZCsgv+m7/d3vvDem
bkc17d/eIychL4PmguQ85k4UH1RuAz1wErBRPKxHzxx5DNCOvZyekphom4LkotRhMqxniBwsGZDv
2YMASrjOhzxJAZWyYcKDPFFl3EutXbpTUv1TBf9UEfSK5RdlHWiRm9z6aoSHDZx7JY+YXcBb33Dg
gAX9eKThAu7tJZ/Rp3BFhrYECTm4fctP1/a08GUqhPvs4ujtujaYos7wBZ2K+nhOC1DxKgfN6Rn9
Qt7utI+F/IBzKbGF503jWflU3XNrYksyB63qz4oVtNYJgz4k91M8ZNT3O3lNthhuxcswuoZ5+sPG
0W5xBPkctqFntrn9HV+74kHAHXRby/aOLcy8NgRtiaCumPI8EKTHLDXlXmHj+clmyjxP6vryp23u
cNOL+z5dXs9o18FrfD0yNP4YZsc8+tx3r23b4ldOj3qTRs9QBEVpcpMI0C+tnyrKslbO8BnbGeRB
myyIGdFYML6tAl9xTwznD6CCBFlvRvC5gMszgaPiI2JIAYbrf9GiGx/rQ3F7Ac0qLiL1P6Qgcyxy
fz+MIew1uriQtpEBme/fO2Kw5UfRIllYM45avOd37ICVYZdqK0mPCzYnkpvb8gBUeyxPvFzbXXyA
BN+vxEXsOy2Q3TCN9SsB85OEZGu1nReFIdKJkC0CGUZxFWshp+4LHCC29CpuFESJzOKuEwDrMkgV
7AK8JIdRs7AyxfY8HYzLyJkfGRZ65WZ6s+uqQbMhDG7aHbvBaP3ZLO7kaQBGX1E+0TKlLRPq0JCN
IFxeK9D8KF9ymrrQ8+osyNpv5XQh4sECzi0AqUu3b8fuBC3aVDNUTjjMMKAxkH3VYrhfRQpbnevd
Tsz2GY8ZCwOUgTVQfXR9uep4mFUqMU/euKPWmNdyIshc9HIjb8JKaOVGguwjf/N8HoBjeg4wQ2ft
9Pxf7P19tNL8zSC4LPX2xfr+ZN4+QFv2ELqEb8wwWLs/sSKc4HyEDSpD5U6M/KjdIaag7/P0kJlh
YswCP/SONTCQAhdwwQNIYbWRHntzl7qXm5gu01fzZ7whs2PyUOcq5fz3KwOVM5exrmvhCjWLDWnI
9XmRq+EvKbiYs5oaKreF70h8kj3+cHHX0np961YRgpcaDTYowMaCsJBCgk+T5XyGVXmLJHp0d8Y2
UUp5j+LimfHAhhrHCzsVydHo7hmAL+i8TPhlfCxGvsq3PKXgrRDW57LPRgKulF26xuIQ0rBIZqMf
dSiVq53gcfR41nTbt6XBxvelItsCd7a8HZe7QAHPojCF0clCXSVK23OLYI9ZJNwOx8G6YgkB0zBM
sr6n7Vn3GF6ojtQ5lpkruWo+YfxjlM+py6dihAHVgFtuW/hZXFsFZIYwGfLTpo63mGjtbMWXeNi0
khW9bjhP3wbYz3P5E5t3q6XOQxNNroK0XEOA951beOdU7iuJk2DnxfPqudfFN1qyesPMURVFULvl
NiwumIQ47ghDCvUVDys1iB2j4Nh63THSbhalHaxJpzOXN4wfivjO+6mlntBG4DjRxkYgCoBlH00l
3OCBIlDS9ZrX04Gq6AQLrCYi96DqFSr87VzuNsL2CC4imqRyaxlf/PqOCZ5JLg15hLOuwmxW0gIx
NKbIOjguaZCOepAj2gymHiseDJC7Hblt0XeIsd/HtPZ4JJSIuRvAiAzWWXHobbpbtk6S8YmsqhYC
UN3pM/cZA20IfAETo/S/6OCFEPc4HTxyrOJ8vxhBnwT8Ugtq+wbJxNbXx2/k2LoWPdCUlPi1WULB
03gQYiddjtU0hBQ4Liz+14frE2G+hT4AB5zlSO/xkjl2862zwwS/ElmmeIh1UdPJgqL0590ChY34
Na3urAQt9U+3kLpTv9E081Iyrzuxvci53JTytsjJXrUBz2ZgLx1faY3hziVC5eyKomaeQkKbGbq8
sjK4/6Fj8pEPiR8LwwON7Pac38RXOm5IItupPgLe6qWZk8J6VSrr+CG1JSrlXPZSX6fLrQANDPIK
F/wFRNEFi8+RZcrSmBPlFtOs+wquSKC6Nz/P4xipJudt7BTsxbRDK2HeRYdBMoKXRlFHYGnHxf/Q
GmeBEOF4riMrcvv3r0D4kWVmL5bc/zixMBWHFHVoySpSrzn97c8pAIGvAeybiSzmokmREb37R5H8
Fip8nRFloFuRD8Hu9APDaDSo45rVh9I/r5C/rOU28KA+WA0fIMPm2N8Oixe39UBXq4lJr8nn2vy6
oHBojWmMXRS8Zlp6gEiQThGs89tLyKki3WxLuzvCKGQdB/YgsHfFLxKOiAecjhskgfXlND+QIDpW
OAGNv32pjwBwPty2ik2eHJKz5LGLPyo4kJd05FbiEbsOtNaiw9BY11Uw3raFOJpLhRsFvZzkyARH
wYbp5STb3qlmbadSvjl/zDWd9ytPCTTajjvzlwDvSjoL67W2KCdwXDIcDyrNvS3cvH66gLQ77IGk
+SCeEl8KgF0L0TQ0AwGYDx8MOiHiey/czYzhOllkgvQVBI1b32Hc1mRfvILQ03IJDj/EhX18JjtR
b+rwHc+/u0SeQDiEseCfveh9w0AWAu7rMJyi5p5pgsfb94CusRxq8fx/F5g2q8XgQsCxKAVC8pws
hC4VeVfXLY6F69oShRVwI/rPCyWyFh5Gnrye241duqG9SzxVxgXeLUrWwE0+fIVxSQCdZNbWtI5L
PZ8aMdUpUT0uuYfkJ1BCE7+Zz+/EPfj2HXgxhbs72INe8Pl7aZV1ukWktPscc9VKcpctPC0PiCuB
d4yLZObR3m//+QmxG5HvAENrdgq+xi2FhcoAoyFsJnlCDAPXNb5V7qTZuVhV/UhVWdL2AkOOQvad
7p5cLpm5JS/s/1anlmP0uIH3p78LSbkGkoS8JwZ4X/VPJhXplQaOy4ieGqCRtyhmH3X9ot1hJTi7
5MOgGiPOQa3V90B1vx3dbSDGgSd9G42QzSFnL/c8I6DmrFhjynIYTemDWDmez5NbQInK79ZkK/LK
dd9xLL8tTtxz0HYMca3QTD8wqroiJRebcoRbfrsDCR+inn3jEIqs4Z3QdDBUh3mOgRMXzrNF1q0W
7O//d/TQAwePicZ5rhU6sqVSKCsX+QLCJkgytMFEMhthcLqL8dTurRJwgOiFdg0gLlVBZuvFHbco
kwaXUHtE5hciaoACUcNr2GvXZbW0jKuuyMGxApFG/vBOheiOPhLWysRiKDnuQOg5Rb/u7zPykdHF
F06jXW1e6QMtW3QMBtgRFg3g0S3IFbyma8VUg+x/GuCxj3cGjbrxaifJEzaGAG2uTEH76g4AkFZ8
sS02EJJ6zwb0abMQeXND9kqIil9sPRM86zCixeLCTNl5GMnP1whRmsN4Rl0JEDN5gphrrT6nLgpf
L61opLu7KvUV2puzUhVBJ6WhMDeBg10xuF4OxeNj/A3U7YmF4dcrjhQfmBE19axMLzXsuRj35skA
0WGfAbZLdQKCClWu+pS9dXwzJIS9XlEs6g7v3DU2iVf6WqeULmhgIBtDS2ocdm5rRKaTuiHgP+gR
gEXz+tcjI5J0D0qv3BWoZXjNPG5CEiWuYAImA0tSMYDzQWUUhbHBRFceveQJ6jEzdq+oOGIK6fZi
UT0L8s9J34ioWFHdaBuheLjiLPTpHrzsTu90lvdpEz/vZQhilIZJyC+LkXCwEBinn9saMLrYY1OP
buRYIdhbdXe5LkioBbLNwr/HlzdQfWx8i+gDRFvpPQO8OcpvJvGYRQqiWeP+yKIsCUYnHEwEJ/Xz
PFAcjCLMAOcxm+4WGYRXUy7Ti5P5XHtVC85LHTD3iUIa+gF7J83gXTzf83vWlpZSnsmRmSAMp8vw
5SFgEAFqrLCBdu+RzQmyhZKRVRYFlm/GMh5x6yLEZasMyAfCRLaNSIa/4Jpr5rLbUSOw2n9QkTBz
Sqb/ZEtDqk1DwTHMJ2cTqoSCytCFFhKi/fhYHINo9zJTNg9bhuwg4/KMvF8ckzs9Nx82Rf8FOhZE
lqYWdOtruFp1f6ECFYPPiJPRftkJJio7u+yCPV5qxDfdbzgDM3hA8Wf02a1kSw45Ah8mPi/T4kpa
aDVElOazjVOK4hDBbH7+opqKvZ5al1e+z0B1gBgf04jRTsaupamVg+rempCWIJ+2eTTxbhcRb8j7
emBv/ulGWFx5jjTKG1GDyRl4gMy7lZG3K4BJHg5vmGp6j9kaEEltNQP3bGD7WLKNuPT5VU+lrCVg
No/6ZvR9JcNJ9nm5iPYq4mg978NzpVoXXeBAMzaUcxV9MKGeyxcvcg1ouwM+D9KJE6cNG8w/gdEw
SF52QlZmPW51KYrF5v83wIs2BW090qG6+oBknNFE2JSn6Fn1vQJJ1NtqGUGSupp3OJraJSWdi7au
rJpC3YIANeAvs6SQCIznzOAv+OaTmgAOlVP29xn8akSxXT2LLVOsseW/PcOYpKefHW7lCty+zp8h
Lg3xeTT8oYpyF2niICFgNfvCYVTiJxOGkxUm3YyUCTntiOE7rlKrItIclt+9Dbt5o7sHhKNhFgqc
ddZKzj2S+nv0pTceJIfsAfeG305AL086CTA+zcH7/CHxpQcAGotH5nc2mpbXWroccc6rIqBEqhXT
sr/85mrC93rE9Frmj4UWPcIUEC3OxbkLeo3tZfmKMxPColyrrjMgCYC+06qQxF//eUxG0sWa6ju/
l6ZcGUfYUUmo0E/lRrf92iZP1j3kZeAlwpIPq2Wqca06YQH04auIzp0+ynGgZ0qSNSGYc/M8vPS4
Or0p7HYrLW9/8PtABbXgH6XHYQLrnUBOwD8DAVUMaFvW+ZAuZwxax4/etVvH0Z3cyLubR+I29L27
nWrN06IUBB+JCgXmXSSBUpvvSO2Tw3Nuv8k99+OJ7o0kA1dVWXaUHtRhyj3uvx733V2mvRioZvFX
XRh/32qq9rxFI8aggDEWJs0QeOn6NSn8C3nfMmRNdebGiCFfNgPpsvZm6q7p7xTCpflczdPNSbhM
iS9+TH9N5jNPL2gphz8jxUz+XkdVJK7Wb0tE6I1KNHvynmrN9oetfWAEGoj5rD23E7bL3l+iPu11
AslyTjx0+z+8U0OvsNE/E3wz09hHn0JXNzDewgdz/FBJGiCbzmcY6caMb6YX1A6jn37ixnwL4lXN
YJPHfg8xjCfrtBTpIqRAiJN8Ld01OwoXWtYIBynoDALo+7+0xyfxdF6mAQK1lgSLIW+SratieWOb
SQpzANeDOrteaN+37wZhcJNnpnJBssvi4YfLxzotUx0WoJRlZXEg+nwDwmfl/w/cv4hR2eLhDo2I
XWsVaLasv/sFA7u3YuWNg5xM8bBhiKcjQm61eTG2lMUAdKK4mWzJhCzh4GL7fnOHgYX7E1Pb3zGc
GjiHdWVO+t9KnGgycpXTxjPrXeHdod5P/ioX5krfuYB/JG5HMqhYVzh7uFdTR19K6aEYKuO8vdPM
RoxvcZbqCTVP40XAWg0T04YU4jW37SXLGq+Bg68Ho3pOXD4IcHBEKVSiewNlFwQZhD45E8f5h1SJ
3n4A70Ef56Djf76dT3tAon7SfbXyccXcMliUDQrvBbpEE3nYF6nftQy/RFouyeprKpj1qyjwRsp2
pYoJHGkR83zSf1rGVwdIoS9fhAReLqokpB9yTs67q+Jj3FwZRq8/CzU/v48FO4Vx9CtLaaYE0+xw
Mq5EzFzZN2loOl0gn45/NQ1KpMQ33zhie4CSPzILT9MRCYZBA9MpCazLnWj8CasnAw+lppgtP2d9
YzwjkiUZmmGmPiz7HyWxh3q6CTAwDt0khBocljlapYUgDsixhey3g6xDKAVCj/+SPv7KKm+X2mOY
w2+UU2Zs2XIW523MUVTqcqeBe1qrPtnoac+Dd6M/oNnb+lEO0g/mLmyKaBZ8HM9opQuKXQFkMwgI
NV1v8pYx/FYpeI+BTfOpRXvaTQqUffGFoKN8muoUQ+4kd0fDXxK88tjNJz1btVQW2w1jXXdeDxSy
a24PE9T8HtEYP1WxQTh24Q2zEZHkmmySeHoylv+mwNlFspcNCaqihW8qqtNDcJnlmDWWtNrA2tw0
4nPlvjEI3K5GN7KI92FGfDVZBIorNQgaLG70l/yptng8KbljV2+kettxKGnuke2dJ2FWg9xnxoBG
SJq4AqDvvtnyugb7YyHDr+VZQHVleC+2tgG0Rjf/RHoIrRAKNp23YPWFA6j2oCpHHmjWApLvX8LK
iCKknrtI8/nmIrIpY18AGQ1Usv9at0o2qdtEAv6/nKQCZgEa0riSyg+v5zxDGPhFBUc+56CCJopM
zXuoZLWjrjzXPB0R47sHmkBlSJlY75xWjp2Cw5YH9QVEzoy+/h+nGEtUinFGs9YB9fVQdFMnVg//
6u9+fFkshqDZd0f+mtakPCKhJxvD/ELs0Qi2ld1Keb338YlaNzi/t5lHKETiq9/bf7X3ZzPNXMW9
UYy9fBgjCiuu6kwfowy+kOCKAckvUJ9DKr9fEGppZpClJtgWC3qmbjWBmn5JZifi2m2V8r60+1+w
I2uXMziYmH0m0fg1a3Fk1E1KeThh7/qLM2Yehipn/3q4+pYeUVktepsdEFNKSkDDw3IWDJyp7ePO
L2wLAOSoXWRJLRIz/BH5chGdanC3Et29Gnk+TVdq1cdPtZRFmwKyGq1fxclO+p4/Rfn5gRFcCPvB
NLLjBHMWers7LSWywsoH/PC1iO6aqISAYihlFqh0xP6+yorMGgYUq7/EW1nA/MJ140QUE0HVkG3n
kSgwH1EirUjO+ZiWV5ch+kKSxixL6skBAxiK/aipCbfZe0aHvVbXhy3kjTKh/0PV/uLGDcQK4LVh
uDPnTRMrYj8QaaiQVH2pVCFpiY9q8wEyIfezkp9220V/TSbWDX12oOnMOVUVqR4EpVUUewLwAv2C
KJ7sna6ohbcImtABk48VccJOsB/ZbTTemHDEcaX2ZnWFejxeTTr1GIdScqkwZmDohvrdTgczaRtz
uf8lYGIfWfYmk95YtTxPodsBHfIYezrp1ZabCGnM2HE+zrNl0HBk8WIRdE87T6YVIg9/LJbgERd2
kEBY37KVrFR4MI85uocHj4GFzRUNuGzOktyIOUx79eI4SVUOIxqxkEkycSPLcFCqfQr6Op+xPwBg
LlTKSSqCodJ0z6vHxP0SmV7Pl/UXZe5k8fIv83PKCpYuKSSCUld9YsVVMlO5txFtmZLPZfo9qcIq
6n9kCGBHbyvIkMHwvF1sN8sD4J9+J/i8G12AtJINu61vPtzzaGYIykx6Jn3iOdpyazwNL1FJQQPz
t29RhF+5dxIsI4ck4EKblDXnse937DfBTzTn4FmnkEwKUU8xMedQbuRUVLaEjooIak7BAwFsawO3
Y/kr2jSI2BhEy19RjVcV34N1fKq0zTFYSwackkJYSIgrceb3HYcWOpc1OgDbmjpg5XN+sm+JD8pw
I3C5OQNKMwrmoQtp8ciNDm486/AI2tidbsUGOtdu6JG0qjTPEGZOsGRAetazKQC+rWSqsaOR5l0h
ZJHFBOtnKSMVPo6w+jMg9VE2gywA5WmJ5XAP3fWw0rlvO3ZqeIqXFiHfzG4dg/gTBqwp95voQeLA
c6n28+IYnDqHBE6E2dmJqSc5ler+NI00Aieenhavsh09Qk0/DG56PNQAMoVYT0+yPwlmgw+KAnOu
0A7RczbP7h+DYOpJjCDcuiVuon2+U0ursvlHl7WT4l6kctyMKZx3dEGl/fM1Djn4XdTEgqZgSAQt
jTYqgI972luravVBdCOYfgbDn8r0ci3FuAavq16yM1uIPwodRnZt3JYi2ZTOxycI+EOUmkqYF1fh
68NBwh5EC+ybM8/1M/hDsw6HJt5zTGITLi80gCQkF7c+3zzszpyOc8DpCwyhIQ7Zjh0AfFrd2Nfa
NcjPAOwHNQ31S1rNeKQBrvzbkrpS8GUfQtUjU24Fs6gSKOGxkjc8oWw7PN/+BfTq4/epJEDKPMJC
/unkASxI6ltTuO+r5tB3WJxdaAZJhHyaLuulJCsWwe4QOJrHdz4gXlTWh6zWavXM1Zw2DItUd1OV
PsfeqCRMxehR7dwHsDE2CdZHxQ+08esvDWvucFKQUELJqqLYi6UhDAaZE6GTcyQrw5RrFngma5Pq
CQudjA8HC1f2+Ns5usBBSM4JSLxruWUJE5vV35ngdD/o/in/KoMtXGqgLiv9o4ftp6TDY/t9mt6D
GwYWasfbZr6DyK+WSzvKftmlOP+NjCTtftTSLLXUajHuFEora61j0eWDpdEdArQI/qcWzTDaNCS2
Lao3v9kzzjmYbSZQiz+utvIiEIUPA0BiUCmCCDr8Lnoewn+4vYpVXphZtSh7GuY/ymepW9IkjKb+
cVg3CH3BJHMRIwwYurxGDHtvkHNl+01U6yD1cH2oYpth0vPVldyDDWADHoUljLuYKGnsCDesBEcU
6MXkPwssoE0yhqBTKycmBcaO/FdKiIJY6VpiVuh+1SXGrWSYx3RUwMeAQZr0uAodf+Aa639QlrHu
8yjBYotC43l98EXGZbnRnnRbYsLAQey/ejwBKt+no1DM6GhZZVTqYtXGDvuYvsX7EuHrKtLF4MNa
JwpHzePz3CWNa9ChLhWdLOWLPMYXOAgEHDZWNqZolcGVF3wscTbLJDN+ClWqb6kyPfc8+9UghBBK
au5dy5C6fxKszN897Y29bOW7YgbfYjjXrKc13IxGJtQxfuedZyYJL7T/NCG+YdyhOVul0N2A3IR9
rhiiZ7fnn3NDkQp0VjI7T/x7wa+pVOS6cdX/0zSB5qrt1jBS3BVqk6NUgGsxYzXdZ7RRBEEY4QKs
fa7aSFsDgqPNub+xqqfh7RcX2Ik8S8XNZ1XbDRmk4zjEfeD3r3Qo8AdKU3tpsXfFS0Kf3NP5CTMz
gOR6b3IKhqVrI9WL4ykVwT8eOeq+J3EVXF7A1TQ5ZHDuIbbrenIwgjC1yEfKdgb4EOkxk9qJQfQZ
BM/JnCZYOWqoyFHEs+LYuOdRueauD5Aj3wmRj0Omgacxb/qMZx23K404OqTNKRh+XLfumVjB27Qz
1htT0x1eu7m3gV/NsvLMn6IKkevU/27bwaAlh+TbsyD0sTSZGUWmEMm7o8Od37Al8b2LT+wqeeaM
734czKAPw7tyO6vSMOoY3XkQV6V0E+IogjfzJNdUxc1q+A+oI4GN8RFbzlG7F5gxECPYbB9jRIkW
86E78RJPrc8DqSPkqbdtE0lIvCTcoq44bWb+iAMH8oQ365n8IxdeIlHJ8rBnBa/wHvaOyJb9lhtb
3x6srYT1nTx08SL/g6NqdnwLaURyHNqhHOQ+0q8oTXerJ6pqp3aavug+7uRJ9vQMnBsgfN830Oum
TVVwLci8EoSumTkeECLNwOOgaqQn33f+J5FTL5a5QxcyA/Oc3H6+PbPSzzlznt/DW59vJyEcdrCC
vXsTcL9hlxH7h2I3wkNfjrxqBEPGjlOldroraph73rx/h4gUwHoUstJLTd3O58enhEM/DzYfKxbY
OU2sE62nolu7FsU6l+BP+QQGWHEXJipjbl87+DikEWfjiaCUKHAaSBnNke4X6ZIdY6sHULFHrdJz
OcdCceobFhdm9uBBQ8Ru21ntlOuxogKJQYgLM7YuopHa1BQZ7hjzsoltL76U8T8XrxAsGvH/XDc9
f3DLF4tU0hp8H+Rybpoci0rIHaZSAGYjzyC1dUVtD13XwBOnT4yK4sGMnI+JLKW0Scvt5xm3oBCH
XJTEWgiN3d8S8gdEC0nGDIal8NHId5kiykYm9qwAHrRPMwF6xj1CSqCT5RQnIxjzhV7omgpuQAjA
9B23lHg2sNVgBbWYLxyHDVpBhXZ3mm+tw1iOJoG+9/5r1lJTkQegQqE12R0NWwuxaGHaclDPK+5O
us6yznkmYIFoNn0VTns73jADz12PNFX4zUqLa01e/S1IArhUDT/6aD2hi36A/BlFZdl1w99dI6YG
NMHe8Z1O3Asuw5FOBInG226uzUcWUKSLtm5uce52zdRwS3KXEGNEOtEBr2ok3Qab05RMUyXo/f/k
BWD5Py9iWdv3q5s+2wdLVarY1tzHQ2oqbwfmmmgOlG3lQMuF68V9k2V9zXbHQawvLE1VN+ubrKGm
S60ll84ypvZCmZR0snqriJ2qqv5ZgtezNG8v7vOjcGGQcBhwB/iYNbRTSKl4iczmUm/5eDf5GDVV
qqzj0TMNS/t5SBAYhfi4QdtMx+Avh2nTNHs6vQKfyBNGJjg62U1mX8K7/YABW2E9hdg7lzBLz1se
4UYC31VyW9Qfv85nHXliuVlsuybbcFpmaOJGjnTR3R7pfm4hgYoIUX0M41838za4Jot957DPQLkV
c8bZ3/J2A2EUWr/pzN/r1FbIaJ53h+R/hD5ytpiQ1KGMB79c3b4KctIUD7td/LAzqU4wnnSL5TZE
vapJnovekmTOoYzgqUxYSpXe2VycBGJ5Waq5vFEqSVtf9Fb50C4WP722qWagW1Udj8vkDgtNVujU
2278CGnmcEZ84O2cnWPzGe8EewkqmN4Q4FkV2rpN+XGc/lfpoRpGmLBfsU2vLvWLh3wpfJP4NAl9
NGw/Zgafu20sP0T8SFV8Dgh7MZ9ObXa8T8ZaiTafsgo7U2M+JV1+QqL/B23doV+KaTwYuylNL30Z
louOtI/nctccIE3DI8GuiT/XOSZw2/ToYqKBBlEslelqaarynTfydnK+EKBSJNdMG0xhzrVaiivU
FpZBvK6rgjtnsVdrbkRs6Ptq2FYQ7Kot4Jwfv4+e5fAsu1n1FMIzowc1hNDXRaYP1T5fzOwWS3w8
XVP2UwjRLrC0tvs7YgsXPlRzwJJ5csPbgbAkwTq/Da39BNfJiZgoA1ZvgthVYHvo+NYgwpv10+RT
H4quo+XplB1t7z9Wdlj4LXJv12AAiL3OOSrtAJp0ufu0tlf+Bdbg8gUZwk3mYrl6XnrFCYR3wsjM
bCMqiiNekBrJq4ok552v5EmuRLZ9FmY6D92+pmAnwOL6PhWoWFVHh6Ovx84D9T5Z2zuagrCgCX/P
KXvUqmrgv4uU7eCXe23OQvpWr/vKYZJRxliHNm95o7+RULcEm5ib83tJK3BbOqhn1cZWyQIOJrv6
zLYk/AmAwDBYFxx+QbSWqG5yrdr9FCsxJXhgZPjDt0u4Hyn0Ie3DEbeJpH3hymtLFc/eQXv9kAH2
6zWANsDs1eb5AkZJEpjFTrkjfk2WAmfEe3C33FgxnPmW81LyBTFBtI4uFUc5h/rzRMKKMXGLynoe
kA6DaotvQqLKIWcuKQSvNiaR7Gz+BHJLW+OI42Ii2D9KnXP2NGXA0qzcrG2/4uyzskl48zu+RMiU
J3TqyhMiWoRzQNJgWD/qKbBAARi5r+44xZI3zqkbAcq9ZtwIdZHGBpkN7SURGhJzV6CIqcIdc84o
lB2Lvdo1fX9/hqqOzXeI1ncS6AvM9twArZOY711GiC288+guDkgsqh5yw5NW0E4BFLfjV4erU2HH
EvBrvcwnwajhqz80tkCMhOYuRk06dyWdBNx/F2KNOqD2xE31AtbNDJyDy1te6+G3aqAdMhrMK4wb
vG/D56im3lRmoYQ5+XVZjJeptAjAbcixcMmOM3W2+YHnpQE8+//ciY/Q0pC08D0e+IV9psz3BjFb
qPt+eQith2BnrUo/uU+54C3H3rAA1sw7TOxJyITcQuGE54XG8Cizr/BWQGPhkuOn9Aadxa17kKau
dlVJA94tFh8dbu9WnOEuac4UsquYa21Nep2MOiXPyI6yjDFLSNOEWgHbXtgP8iYfVj9RVzRt/P2X
taKeu5j9hP4k5BoihHpAc3xndQIayTNuZeV2GloS21hw0PSPKw7ztlQmSbX9fvqJbPIzYrZww11Z
KhCIt2hN+7tgXtE1tc/AeUV1uvRkirbmoXF7x4qOmhALRFRxum/hs575EU6QEdTaymD4f4n4LEqR
zhF2tbkFpMcpBM8aBm9a1YksTNf1tpGzEixUzLLwl/SvBaO6qmt0ynmRwEH/Y9UIahdb3BXIqEbB
TsrMpwZpqERC0hkumDO7xkb7hf6atAxLT0tKJEGkF7rHO3IYfjc87nmTFfe95rmZ2JfEoYzK32s7
SlQE1Q6PkFAScQlY+V+2sTKciDM37ogQz3tCPWQot/5/HTvp4QndWVmZkLDOyawtFL+SpwOhEkJG
ywneOKfVdj+617rJV5Vja6rNfcCaAHra1gDwHtpV2cuyhrPt3mzperwBaG9aBxG8I5AKo+2YC9wD
MnUlqXi6RIMNzuswTB4dSALA6r48XWtjDmMjKAqVcA4PUHNtHjB6o2x09AJM8r4hgDn784ZwLZN+
Gz2l0UG9qpudGVZJwlGB1TmYR5RcJQWGOKVZqdMcPQIqJyi+8RpH2ByXTpV3kFECPA+aE84o2CQ6
CXvNwYiL5cqg/FW6ybMPnlGEXU7+PaNaryKioM6/0YrxO0c0ys8NOTKa/vRoPSVZJFoy7PeOYFeP
Wz4sKiNRDo7EwjBmpQjjyUOJbpLvN6Dd3pQp2TDFC2pXqp9p1lDK8Crnd+OuovELPUv9Xgz4FAit
lDrAboJvDRz2UMVG8ixJuIf+5LYqOeOjrxEnWb8syOSr4Nit41yS3mPhl5Br0UmIdK4EWoCWImcF
1prHAb6l6TIowgMA4HYt14w4iyKycEQGiilGaai1mcXPWCQPZEIgck+12b/LY4TUIHx7qSZ71vkX
laPVevVgFPXZPJy3jn4Zc6MMwNZiuwx/zyxcbxg+uljDc2E2ZYaFwVKx42t7K0K3nkexuRwh4AG2
siAhkh+bkFoxmvVBlmCnsv3btIufML8+Poe5PHG2i+ZbP4p0Uifpi3MccFrEKp7oWIBPKSA68Nm8
HUVxjraldYK7jJ1ngubSEfl5bWrnl4vyBbb8t7SU/aOWDm+andJWUUViryAsluavwfiXe4Y/SNHn
V2dGqm+WE6M4S3ZRM+nVZwiRUPEW5/1XmzARIaWD+YlAZZADh0kdb9hQklif0goz/1CNJ9YtPmHL
lJrAK0Zval4X8iLtUH3PDZJr65Avh05pJH8Yjw4m4CqhO8IvvQDWO+ii+xQow/h0qkiSpt4+ywia
lReeCNcq0sok4T6yZZJkx5FcJP9Q+MiKOCcwaLNEG78YQP9eJIUBB76J334PSuUVAZynAtVVexOm
wJ/XZ5YST8/0YmI0wRtTPaOpmAw2TBzuLOuWhAx3CKIsTrsQi6/+3A7wJPzXBMNsImY6LQcZB7w0
iv9uO6YI6mnEwv+l+PtBlbEfdBIwHxJ7KqEZp+0A0s+P+vJiBQmOpXY84XFI8iPNLQiZ8X/dg4fQ
+c885173B6ZGUSuzTpoNUrvexx27uGnQ+ur3NTmWbO0jAZRd7GjAEdmZ6ml2F9jaCLRSCwIR8Voh
ksKoiCE4ufk1+AOQQizKd3vs46gjT7mYXmjhW5gEsxdHVT99F8B3psytPouucRr8EAac1LEYhSWd
7ormRhfvUUd+xKhE3W8x33Xarf4nGYMcl/1HtvoriRRvihWiwTj9Y0/BDZ6/PPYehtt0Xg3olFJG
N1Y57WYfbq0WIfEHtYxBRNH5FXxLvIGmjX1VfbS7g0/1ZBaRSHWECb1kE5Bx30V2XdyXm7s4BOgf
EQM5M2PPXm5a7Kz126+pEckJPYQ4OB6ONK77yDpeuF0DDKMg2/CUjN7yHe7GDz6as+aiKxrXZdOn
FMTGRbkYmkkrGTcDEAMfUx1Af+o2xyPBaMEc/1j5OZszXxBySL7chG4sv+1+YB+EOXEJYjnNK32t
CCOMsBtWotGw4D+Yu23pSyXMR7weQalOdX9Mj/tdiqJZQSSx2D9R+ASZ8ZVVlZ5/iZq9XtsPngF4
zvLinIZrF376MYHbmXnF/KAx8rnUfFY5zFG+LRdyIuPmUOhu01PwUMXicpAgCDT28j119E9v4Nw7
gdCaltJKPyxD7AmtcDbYR4OUMk6hoOKtnfve7/wPX5BOXRfP9TaciBl2xBdl1DiBc21iBIOrFkjc
o0wD0FD38OTqSXHXu2RtW97grNDUN2oieXJTIKDm1Q1QOBYvOE99rzY9D5J4mvvSmBONA83KufjK
yECwUnMPXxE/hHrzQNLJm6e+qxSonBBys1vPbQrzmsaBToYqrhP8CgEZssTFsSNeZnRrn14T9gYF
kvmxHnbUaz3JGj+GE1MTV1YWO9KoawRidA0XZohZ1l3tTKpuBN/aTVca+YLwwx0SOZv5Eb6/g4zH
SXzQujXMB4cQj+ncy4KAbKGJi4feZAnK92kldHglywJgdpU6F31Rpk5rxYvXAOVjEmWfX10oyEF0
gHz/9aWQCWHqdJuV0ztTPM19HPw1LWMVdfmDQXzmkFHDdBwNBTa+Mul7WNPW2wOhBTtgwWQHXhHZ
eLjBQl9TOs46+6/TTcRwbhoXFK7geKilluSEk3a+R+b2Ntw2F9hd0zynjHRFNmbhjxCUxixjE56Z
+wn1IziQWRTUa2fA5NyhRkuhS0DIIUF8ONeXZyY2diZzBiqt1hRO6b0FGAnGuTwll5lRfZ5mLNZt
1M4Naoq23+VT/T/OD+TIlMPBUiMuzKPWdu1/uSiuCu9eoFYJjEKa51XiF38omTEtb61g9+zyQQT/
caktCdRBKMNTCWS+ssrv7bKjtwmQKM0ojhf6p4sDd2huI3daBHNzErtbpwmRGneHlsWcY2k2mwxT
W4VLa4GbmywZW6TfNgNCD9Zckswz7xtDPWE9suCNhoAT14wj+Mcme6uqGM1mDyTyOW10r91T+Wy8
uQIUe4r706Ih2iCzO2vnAtopG2+orM0cpwAbO01ajfDld98ErMjwmTj3iMXF6Z8cOaNJB6L+0NoJ
+B+iOKiOv6VfAkpPoLqTkxfYoxCS10uFYnSn2CZOMZlZn9EZ5mwtkvoU12EVi4lUZhm/Jz7u+52C
Ad9jpt7KNSBQPuoansXRmOvX+3tqatlJjLxyBFUCDP++GyOBLiAEGMAvb6l4lfXpq1yTeJzu53Xg
qMi9aS0WqVrakiKFrHxEjda8kxkgbLRcErqKcBdIupyXxnY+ZG0WS76yRcYKx20jG/Ru2XimyP5H
uStqEnzm0AoLNN7qmfCXzVGoWHU5K/Q0k3injmypYl6GPr9F9I1GGnwAZBYKLcolMt2zvq1baIL8
wqgFpyJb14pOvTid+QzsbJ8PTzHtjARU8/ieLoEObPZDoZnW805Z27pfmJHsLm7P6j+sAiZP2loW
DZyP3I3VwCGQwMW88N4LaXcB6QW4UZblXnWH0O+LyRpxmbPpXRTlFdcszCM2zT7eAQqqD+dBZwxD
qsjCVuxY+NA2nGU7IwGr/hCsG8eoNoDvkIsyifGG5NmCdDH6rSzNmxLU8JSCkWziuSvKhOoCro59
LuGK9at5gzvWAS7BS2eeIXPCd/ByF9Axml3loV9w+YsmY85NQodA8vVe5aw6PbuBGFrIWMeguTZ3
H52oBpkv7NlldwavybGrui9zjLJWagQQudx9DU+H3QOmqP+xpDiuPt36z5qtFhBWzryo2Xo2jIJU
gKOqx7upUuAxCaAkvLnGrW7PIhNDD0Cm5Nh5pukAAYwsiJmN8zw5Y83FkOPNZ3qlW5/4c7RuLpyZ
3Siu9BlF5hbCH/+lqLvmcfa6av4ik/m5hVoafU9bRqLnsJoqzeyyLIoXbNJmD1z1+nzkgSLV97sJ
h455dbj+1V5HtceClzGQP3ftrQn+g3vDb+5plTMXPNN1TwQsjSluiyeIWP0JbXqAbcUGQ54GuHTB
nTMAG0YqxMsUYYygPke0M1ubuFKq5zZnMPduLpC+KRqAvc3/H3kcq2u9IkkHqLSYMh8iGPwQ6Yle
8+Ok9jOtYrfpuRGRRVHRiDxcpXHdZqNJYXcPWKaoLquA6F/dK6aAlnZeEKUEhv2zdPhg3n1T5EeT
u75ovlaAzh9RYH3Ss3wIyjcwbXJ+EpcBeCu0o1KIR+WBD3RFTGl2s3iumGmFDFY0fwRnA3m740zY
OlGO/ALVa60oFbXV44pz2AZ0aGI4FSvhIqu/vxQAC7mLH7LX6yrcvkO6cRK+VdSA8kLBfw+R/8Wm
PL4o2qJ6UX4ZPo5/vOPXjwAkgI7hSZ/HXMztALeSsMabM7fgnGLe1l0y1hTE5JosPZCthiHqHtsa
EGvHyOUwawElaR4q0Cz/s/w0UNEnTfMeFsTCfvJgM7Bs2UQJQuQTr7sJSsC9iO6Lxs72zNk4PxS7
7H4nELnG8YUxE2P+KAjpYh0xfk5SZe0SSakQcGUxVm4osjBhSvOenV4t/E+9Kl8vhGSfqVb87HZh
bUGzTiBNpXDiJBR+mpyxGQZq+I48kzigw/22ihAXSD84HFjv8ljfhmMJscpfvcntK95EQkWrlqy0
hJvxqIXM142/skPiQxNp6sQQh7fkOhsDL7+wgNzPpoYYP0Z040QXJjGhv4Lq/XNyoKoKI8I0ULZd
EL3QfqXEb1sCaCJZfKIbJipmVWDwDtIhof0ApU/xBvsj3oLKdduxO9qqbuSFIwpIlZFc60+2q+Lp
+2c1lMufKDKS0EP42a+4WVWtq+F8cRHhzC5mUJ37xyRptxpY1SZpcOvbt36YbimQbcGGfUHl6akC
r1DSN/75ZEMme1TerneOPNZNAvfNkiqmqx0VTbXKeTVxu8XAgBCJdvdIrJOi2P9pJUTA3DFE/Ebn
8haCeBEFjctmXLdeUooveUbJ6ytFtcjR9VcH8EOTBZqTe0U595RqAR3HD7dvW7D1g1DZVNVCIQwK
INIPZmzQMgZ1siWjWr2Dr8XPTpCA2BfWPT9pHtzFbbW0VNFL1/ExM6MqFTXEsxFG9FBLAd80J/ig
GRYGXE2EpOrKsralysoJNIa/D7X1MttRL2huMNWbpv5eYbtj5KKDs7LAUHygdpkqYitDbim/AFWt
D/SGBh9v5HByTIoNSIN5U3Ao/LAtYUI21BH2/t1hDRPdu6QqzrBYvKDLujwlC0x43yWwX8RhghUe
FailxB4BpKfHxdInEYOHKML+KJsKxM2BNyCq3HglWm1qLyFp7Hza3r00qSP8tzMinNCCYqsUJ62T
CqZZCRvcoctLLC3wtVsKRKE6rO3sKVtGhkBtdxAdBWpNPzxeABbiSNqYmmL1MglFc77Z68NznoBx
jOseUOFc40runAlVaQchJO2cR+W/+0IDZoA8+n6lHAAQf/0c5Oo+3cSXKFlmeUprwhB6zSZ3/7rh
w2XaD2uIt0jWc8NfcfWghxvyu5uEVl6D6CELHL5X4u61vWkCKHtEhpIzVVHT3gUrRfdNSMr2uD83
sXMBWZklrkTR02rupd+g6pLKXSp8K7lwGwJ04xkNITrjf1n8f6AWzB+TJdB1zRtg0z2Omxti3ZzB
UDbvNCQeExKH2vIcugQPN1aBrHRSGLlA3oJAHtSyXhq0jd3xSHR3F6SpGO9nVoH+cigxmUTVIV9S
/hifbLezwUACJ5jV0x3IpPheThTAkCILaK8d6WRraLhYhKrpWQVZzk3HtOez3bXqqkWP+OHiyT5E
V57L57DXrbpA5qGrKtq+taMN4yoSxJklkh9aBvN2Sb8WPmpoJNr6ExKvzGLn+Ouib2veIYCotoOi
osNyYQPK7FCFaufBsSyyaL9eG7s6tVVmavf+eT7e+LN+0TiviT6JwA11uGiMK7erv4SZp5sqoO8o
CNeS+uBGEmLMsNijsSWYWOesiUYbdblr/VpLP56LslNOZTLsV6coyea0lr+jhcudUAMtTOYLoJhs
suc5jcPWeU+lodQXHsAWvznSvnuArKQkUIpWent44El+LF9fLzxqStrEBic4lkWVOuC3n3LkB0f/
rBqPqVUzNOiZ/l17TAlML8pqdirmOBOoO7kp961UJMh23H7mGREqZIRNPImpxabj3tOytS6/GLYP
hjrA1eAZqrLfZPcYYWtqUY9z5rk5G1PUN2+Ou1pWCTN0EhwS6BWrWczwa/Ri4EER2HqxOm/lEuE7
DnkthBreVjzQvPthy/3JCgJya93wXEiw7t+jD5Y41g/KbfzQ4UuSpT8LDTjILlwisGH38nrLfqHM
hFkTQ3Ot8garBJyGyMH6CIsPZWHs7LAs1HMWOZWEvmkhoQ+WijGMhAv46Bpk6l9K8D2Cy7XW/9Wo
VrFAy8bdjI/j/66Vnz7KzwTYc4+iulKp2UlOk/TieufpTaHQfzHRY23x6ubbQkgn4laoax/Wf8wy
abmevuQH4sLhCvOu3CGcNLV1Sj61bUkOnBW2zYHQSNR9kCa1OD0J2SRsvMX3iYpE9mSIzVlxLYu0
hQT1VOPfNiSCBCoj06BTsoaxs7unwe+4aYUKSTHKKIFx2zcQwhNuXGbww2PBzUQfAu237pDI5+zn
otSpQfN+Dkyug+pcV/rZrdi++GhNUILMpjgbSomcS3b9w1UtsSCVbO2zrOZdAtybjU+SHlfmQj6S
Ejbrof3D/2uiYzGBsJCGohpI962/D8EmVjpf9fIQpeGOACyTnMlGIfwq+gTbXkbpLvqZf7xbG7Pu
MPVn8J7nuSGGDvETvnW6ttpMr5CT9anPyeuIryksEly4I51KOdOLCU3jb16CmmcM5ZIdgDPA5PG3
O9aijfgBGn9GhQZvJgXgteOFzLrip82BWLosUpCAYaNo1RW/lfMjiQyzDDFzZnaE+IQG/NPfIlwn
zR4l0dBZJPlgGf9qSf8tdLFK5ow57VX6UDw8moLEQ5b53WeF5A6KOum5eROhJyx/dImixUIVFI22
GN6sckKv7sDYQ8K3eK7d/91zXhJMB/XD7VeabheaWwVkw6YVaCuBQ+C7CgBi6qKwHGanZCpDcL06
kCK8Orgj2xYeP8UM2oA1mW8ARr9G3xeprSp/4AJ9VCryhZzKzBZ2Uz2JEUh+77d2RXUTA0NA3lQW
COzzJ5OAZVazsXJ7V4QRtO00oS6ppY7endbEssK7JVhGZrU83J+ccWuUtnY1a3ejZGT5EJTEY4+3
bLb25fzCfLjYX8IUmcOK0Bxu4zQYIBxj9DdUvu2ZU9i+SRwC5PZmZ+cyqj7ARtGMGD49zSbsXytl
IyyF0TUQ1ENaBssT6RI725zMJYOigW/L3HnJTOV7K8m+QlbNp/ojI3yjqF6m4v4lUELNOUOQmuUt
YqSeFCYhtRQC8ONngvLBhY7SWtuCgH3esu3TxDNB/sBvMFKHxifY8666GErfIQsJbpSH3agkTiR6
SZVcaTbvLhRvN57RhGeguUKG/QeG9bwE+97kJ2poGqmcfnPbwzU1p8a2FQY7wV10xFdTFuEchigX
l3VsuiwmzHLGGH2bwJ++qHzyML7uS3cEuxOi2sAu9cZJm6t7CJE6+3Q07ziPCMgsi9z6nOkQy+50
IzKWK7JOeIYeKi4El4OtxVLEDx1q6q0QqA0MWFgS/WUaobWF6L4esuHHrvCBalLyNeAl/rk7VwQ5
HHu3ycPV+U+ylDWdbnVZbw+Zm0dHN8qKqC9UBm1dcN0X7VRvwb4Zw5sYreWbIniyzufmhYga2aZd
qQB+b9XM27p5dWuNuvkdnN0bJTQktwXGtggDUtD00vY7cYKomK5gq1ygMLGnP3maZy/WaT0WThZO
rAs1SJodNExzgOUhJ6imOTXW+owod2UQ8/11hiTxbOziWHI5LTMWYCEPNQyIsrJMUpYYYwTm85Up
aXl4+FeYclaKXDZbDBoChosf1aCTZr/9xgA8gK6lse6JE3KFI4RvBsq0ZpD1l8Mku0lFihC5soIb
h2JZThmU4BhQJcir1Gz1H2NdccVcjZVN7f03cSiMuqxew9IBxu4ZGnDASAmDlL1yNqRs0ba92Ec0
7SWI57vsChoTq0nqd+63jtUiTBAd45PmlYU5k8Mty4dCKN65Jhbi4GBbwRKiBgM6TSSS2V16jgOb
PZZ6ciqdz1YT6drFDrtuqJTYl2lZ0SbdV6NVFtscakw+FFQAmW/FrSUphaVDDJFzmHVBLOeYys93
bnUd8yhtCJZUSW5bTwUCKxpbJy79r+K806YmY2NOe8ZXyGk1bmYk2qyVoM77Ng0P21y+z4Pjxsaw
e1VSZtFlXHyjuGDueRRiGh76MgEHh/Qq5vOP//3dfzR5FglCZf8jDFWZc7+qy7NMPGp2XZjT5Klp
WJsbbzFow7VbLOWdKxf+wSYhdiOtYt7WK0Di32b6kvOTDfWTk5idaLMnluuD09h2NED5cC7LItc3
EtcpYlWkPqICjqrpLr4/FX6t/jyOWZJGJZ5kEjBNh1olFgCv65WWy7dLX7NneQMvZER4Gxf9QouB
4/i7H28j60CxJDK6oLxapIu3Cl2l+ddW8iMg2+rmcd6Q0ZspINJnru4MkZ2SUMTc4BQb7+Y6z/RW
+dzwtwEQWwSx9Q9mPK7+5IezP2CU/U5fO79jyL4ThDvW6K7NV/reFhI8InM8zFTVPueGCjUaf0CG
pZpXgbtnBsTC91hzjO39axhat6bR7+ZPHgEDci6wRalRBgX1CmCzw+ruK6+MFi9SuV/25/tjVgdt
7KEvtbraaGotOOrnM6MwrnltLdnlok8G8s+gHG+31q7qJif+eo637jKrXYQibOnYia5ZTvJ5qZ8d
BQrIIDJ2rTfEEuoJT6iznhuxyw2bCLs7LZUIf7+2UQCiSgGvBoZtXFBjvX4rJWLjMgsB8DxstMSW
XlfGkX4kXfv+Lh1gzmGg+lRmCQceQP9o+Y1vn6fRO/QGt1OF0HUBzQ/0kpHjaXydRpoX1lkplTHo
zct8B44KvV4MblsszpLtGkeHkgNzwOszCO32H9r5wr9s4LcKN3KIXYin8YB+S+0nSMWLblRExKGQ
g7b8oY0LMXugfP/uGwfbyoSid38tJA+2kWHRPP70QQoReKamEnp65tYI5q35SXvw3Mc+5W982Doh
wLOO2uMKCv5YQbzYvwZWb3vxzSefcT7uaymH4Eg2jWBWj4/sJLEc7kt++AYe/rEHhHz4dc2DUDwe
IxMJ20UJt8uJAopKrv2EU+5ph618Y2FqhgoasWDuCAS+iKDzHqeXXVqbyRknMBmo+z4VvyPRRoGB
fnj/RZPxr6eOvoFN3bS8+hbRUJBvYpeRPzqxwDuWepOINrt/FF4KI0XmQnYdBPbMInHzhrjRutqH
jteVCSBXtJBVCuWN2mDbL08d50PQ9jXjz4WmMxCCkL9ZGtB0gBhAmBz9/08w7QIKrBkMUfoeSODB
jaUjhYoayAVJrFgRE4XBYNMeUjy5m907hxQFO8WEqBXMVr8wt/BdtAOmWSTJp+BGL91hg7g2fxa3
kMbZKdOHLA9sdJRxgusXPdYuwk7eNKRZ0+xQe/waxkf4R7RF/ZtNZs2e2j7AQ8LOKhILZH3b3Lhu
rUQ2nHtPtPRu2sL5uk4eqVyBImdBGXKxxP1jbLMeRijyerr285GLEeURV0EYjF7Jlw87HqGzCRLB
Pkqm9wabM61dvS5u4bXOKCVbQxAt7mSOk9dTjVM88/Zsf+dukgEPRZ8wqfJJU0qvhiNCnOTE9BO8
arsff8NPUkvo6nHm5CD9q3Xrqad2aZE1ecmxfIVbiy26Zr5/gPLM3BM8cq82RLpJnlGcCqlIUHkX
xJIXSpnPirTThC5eRiB1SlSNxrRKbe74yKAxOJFKK23Dj2HRVdtfNOW4hkzCIQybHOxExNN/hZGt
jJKrX8SpMicEo8/PMd2jQ6uHZC/a9DEkKnH7BslcedLPc9Io+EcLb0W1A/ZqIbvVtHtwY3xOXR6R
K47wLLkbdkwJQvtKjAx7y5c5w/AxLFdZkimuulOLsSfyXKE0MG5Bz7QiD2ahdG+bdx/Ma/RXlLNj
imh8QOcZDgHfZbt1OUvH9mkvYE3VNkqMthudfMyj7FMX7FhrGjEyoEGGxrXAsDSOLGp1DFNf9b4L
z5+xXBfbqYl88izrpV0EDICvwaW0FVAmnd2HKn2pDPue8phhrE3HmVh8ZLOfYrTPrudCf373obMP
zLZ/5a0YVkwsjnpUqCWWO3DBpAIxnIF492Bd8yxpx+EPgiAAmjx0U9eNxO7/5NhzLavwtt9vQTZh
n0q+dHAlYao0tCGZ2xOkAl5aib5oGdNGZ6AEuhPsbTPMAVoaK1KU3UGHZyxtCYYYdKiGd0rd86lt
DlJjUejmCn3mt6k2C1i97S+9jPcg89a+j2UXLx/WUGSm6t6Ajhiu+RLFAP6sTSqzSBZwiomEtTv4
E5Z1CoM0MhhPLEeyyeOA2agK8bpWn8EOCJYMyr4Ctm/hct3H/f4O+XWz9UStUyW900wTKSH5ZSGD
abKFktrLLxZWYXKGiE3p5qMV95W5zPhpnHlh5k5M05D9G/EsX/wXJnxRB40ULOpE/aX/2urUHciN
Qaj8ohXAqcgK/xBZH+rjTjKCLQmsawsUiiH/cLWjBUkRmlOvnVW7SjJ/5x26Z/F+4F67IBIjsn4W
T1T9xAFidvOb8fjZeQq6dKunF5PXjPCpOw7SgFOu2XftFdTtko8KyX/IqPLMvLzpDvIp3fu1rCCp
NkkTL5C8tHi83x02MTS1GHzu9gDzVShqjANfYsTFbFDWO2Bm+lW/WRcEC2D0ub2PAtr/+CO+ZhZV
BcuRVX4hXPzBUxYuHCyuq44YRQPGtox5a0USc5teRNc9FqsN2YrW8iTrEXkhdFbgJvScaMEzkIgy
DznBtEacWMOSzSYaJVz4Y5iWFIhmgRUIMFi7wILPolVpkxqHtU0uwcEHMhTKYfyr85bwyUE9zB9G
aW5Z6PmVilPNaOVNF/1CEeXyClLG4b3sINlHRB/WftYJfctY4WMK0k2A/Tio6zaCqjcPP7ode29T
q49PFNa2oUOtHUumwZZWi6SGtPH8nx085mChWuhWMLYWrCilvczAekejIFHyM++HBB49fiF5zQoU
7alfiFHbpGLek3aXizCsnZAOZZoRRwVwJgUwjkV61ay8y/u4bcmNPdtOJof4wv06n0eOzoLsyyMP
85ytc//uzBXWhvx9ounMs+DAzjTRpKr4qg6vkMg40dZP1kjZDiv3BD7Jwrkb429phtNf/RQpSe7V
uY/bVIeU1ShqRFN+gDIsZBz52zHP+TYlgV/+gNBGr7r0TlQG1jcaunKAoy/dupXX+NgKNJ5OYSfg
Kv0VUzMDC5m/ieMDP3x1oVSVHi7fhpHCeB/Ok4FfBGqeyBrfbP1MmpD6NdOPImYleDFORhiqLc2M
tVCtlObJo4WT+OnbzSqrK0YLZ/BjLBsVX61bvAUYVFiLtbKvL0E+DL1WIAmJHDQRd9e4aRw4qjDI
yV3kM3XJ4cHotqZYbOiPtr0cwAITd82ZVzDhwEYKJuS4IRudujcq4pwdVR3VH1bRHOVIYTH60BLq
gsij3Of2P5sNfhplbbzQxXwcnCKYxAvH5GlGsU1+eiJHtoLjjsa3bF22so8TOsrZhG4Lt/MbsJ/T
qasSs4lVCWZ+1x2tl7zKKtwkxTsxzXtVJ8lTBj+kxAU0AKAgKIXGceNANsC/Rvmilvj910TH5k5T
nQnurWwwFi4t4Txvl6PX5IainaKHJFDH0LCIFYZF7ISUZLR7PMyWCa7Ny2Oi6zeW58JwD7ZkjiOC
byhIX1AL7IBas/0lyxRn6D9vwTsTEF1kydTqU94qKv3apmouoMu1vEWlqEOM0/GTHJpYfodwBvWn
PLyUC7tHnaRoY8/+8wulH5D8aVwbSuHP7KE3xswkPeI723W3PPKg9PScc9YQz0fp0syheGJNDYjX
1x7RhHwYIsz2SzFGHPXu20+tmVRE/eWgxInSUJFf/wPp3K4IiR3h0y84+viajsKwHHzVasD5mKO9
tGlYdlp1S/b2IZbE/2SgG8B6QkM+mRl6lxF0DhPn1Il7c7vUyeYx/NtBC8yuok1BOKgDOsjtbxzd
C8/LC8pNhZZGOGnlGg+Ir2zXHmG932aBnPOjuURbCWR5XQUK2XTkC+VXYjRbrji+zPt/Hv2Lm0zk
oft4HWBOc8SIr+O4gtdaJzGNPY8+gP4HJ6BxeBKzSNgQJAZbWYKv9eYUj6hWjws8oBAn8TmMd2C0
WLsMkldJNpRUTViM/yOLtWX5Pe9aSXocjluE5DwwIdh8hHv1YeviWBYRZkrfXyhJ9/elHsG98zBU
61qfc0UncgdQl1BOCykFdw/gud7sYHFnuvUAahi0HRO/pa+tOcmQqiytwnxs2V69bi4f+QEWJHr6
fDCtk2IaMKR0cdJoTq2eOS1NJ1ENnk+EfbbCkR2vJhi3H0W55iOXOnK3h0KwM4V0tmrzfRDQ+t5A
Ojfj/I3S3WnUzerAZTHKve//W/rAYTRG984nsPhpJ/08T0pF3QqZGIfD5lpaH5SeweISd8oIO72r
WhZN5jEqdrWhh9RlvAjIF+b/b4uP9Nt47tDI3DXdfxsMsIOp2ilJuUW3hzuHU38Ehm+8U32lUBYb
XXCbB/a5ELPOc4kdWEOgXizVDD06WFlj867Zo24tEYd3ml7MWL2jQow/ctjEDiu16A/X1VUQMpz3
ZyzHhuBW1oQLJMUn5Z2K4kOlPdH+KwuTBaFowPOIR5l5PH0J0GIFwd9GbBLfHC1cIyL2K1eEAhyi
z7usABDLcjbRTFAtAfF7jcoLo00B50zovdmwDA5N1wl8cmsqZ8Aemh5RaJTc4IlAOwKKwnbCz+df
qndlGFl5fg4jxm18Ft8dIwA+F8xzAhSzOBQN1Pdk5opmvxzcF/gRzF3aNNP+Nd6PRKtLQz5pwmeT
UfX6VL6GKHw3QCJfFq2hK2HuzuNfF57WWkBup11FxbmKmmBZ3gEMyuzKXq0oEp04VHnneDhqF4VH
/nhz7iEWZxyZRFOCz2nrTI8rt8OaKrPIwntPqOOui3/cp9l/IgMaXbUKZ6MghQpe5bltCiyypsmB
yBc8q9LrVoKgY6Fxg2CaTOH/1WWd//5eDrs+SgCtwQ3LEzAXsHLNrLyonzLjDYSxZjwXtYe0NNJA
IfR5DvLT+l0mCl5Pp2aRGA/mFiUZAQrVE43DwTpMLUnQQXD2xr09r4Nt5GbXMr4+IO8X5mbl84Zc
6g7RVtG4ULLz44BiasrpJ0s9Fpl6AApwidiENJ9wkfmLyfmm0oklX/w/UgautQZWIO+wTaT6pUjM
Y+HXugmu/dRctPotU02oREGqQVzl1fi3ASQTV5HrkP6BMD44IEXyh06E8oLeqFmYAKJlWSllnHyL
lBb3S3a41dUP4Llxw7VIbziFUq9Ru8nufrxUTz0TqxNLABC6UJZUfLMcZHWXdKxsBr7WWaMCqRwF
iabISnfbVkRx95+waD37cm01ugRouFEpWEBzE8pFwFoKkNy+jK+Civ8O22TSLVFrnV3A0jszq8kB
bSAASTsHa/CHdpJarKlT+SGJIZhqqlHiLGNdpOwQ5zZzThuSyzOW5Q+Vl5wgamsNGbExBbdiUNH0
LpiHA2ZEPs6FIw7jgqXQ4M6+qkLbXLiFOPaZpp16vnCwcjne/0I3pfJpvZYuFGXYUCW5J7MsqF7p
EgAmE0IbgS0RKIQfTDFg2XFnYkdnU6V/o4nSY5dXBQSmK1ZDYCb22tuERIe0srrDlaj76onFq/cX
5vY28ZxOzlCS1n1phrIfGUHsky8lTqvIqTnJASfWFAS2AunxceR0ZiNvNyXEsIscZ0AY7Ej9OFCY
F7DQeTiO93/moqPz6sOOYD5g+ZcHBIORCsctB95rMMCnNtZHoeVP/dywIz8J1DEDz6n9asayhMbQ
SAHUdmBJ4FEHnfLPHs9xJzngimc+S0oCqF7lpgTtKVfyKRXeiYK2g7RyflaceSC1SEtYo/2AgGP2
5JXSd8IDUE17hdQvbDGz3WWxBs5HTtnLUeISIOKtK8kxdGdNi9gr43Mz4R4vNsBlRgLoO48q2go7
GIt62YeJhLO310uVpExzsZQtC0cx65H36U70dJag7a2UfXsoEz3HPvVoc5aPsRLArmYvA9lmsOSz
s0mTBDqk4EfjLClJP+lZ+j/e/wLyZdZNl9c2rZic6Pde8S2lf1ehxdaTKHpHpyvzABdcEI7D//MR
iPpq5EPI1k7pemSfVwZ/TQ/e9DTYjxhrtkgaIEzrXwVRV5XRHfrxcBs7VHBXlc6CYGQOElmF2vZP
0pZ7a2yXvKGjAPjv1bbQkUuXztp4S5B/zykLjZ2XwZURS+sG7VCZSbxg3v1DWFt9p3og1giLCvGp
09+uHXRfxtT+ktBYiBHQKggiBbl0eZTyDZN5KfSPwD+Vi/9GoszblyXHWHPLsyjtDN1qNv7ocFff
683OQ6RyFXnRwlL8RHs0///csdcucZ+06ngEABTYd7nlFuI3/oEMATAmD4GtgjDs4uBeh3KqkMFa
vZ8u9n3/mLbDsXCjX/UsT388x1tBdG+LWQR++4/sTgiOLDkJT0fJ1U2Oq5J14Wpivs9cpMfm7agg
FTzPIaPUnnN59+aAPWeJqoOXaM+DSwa/bQqYkLn8X/N9xHsnbAPOLOkXInUEZv7ApF1kTkpA0uP7
JmbOgXAyTKHfwtiJ929PXbUo8wGPW8EPMMdiN7UUA8+CYYY6J3MqdL3S8V2o+XtW4jhlAcYaqDeF
a/Idh6mt/4usvkUBoTT9jHiIiyZMOumvTKQJXKqgcbYrT95Hb4Sd/bAJK8asDTng/S+hLyJn/mNM
YNEcRGr3/4YwnrkHF8FCennOzKi0qvxLM/93McgHHjDLKSgyL8S74sgrrgnZ+mmvTuW+Pe4iL8fu
+dRfOeK9bk4amZA3qXoPPRlp63xHs4H3dg93zfoKLXSEaIWdwKVqSLzSkM7Q56lUKB5W31xYlsWc
O/w5MSl1Ec15LfT5TZQYntYnKARXN7eSVCO5BkiPHE/nhgRGCFgJ2y5vtEHNEOJxSgVzG55Mt0g3
AtsPiZsEiKtAix0cuxnfJyAy4U3RbAGFEj92o6dZldzZh1fPTFaji1RT6cfrRgzlGMCc+Nx8nDe/
5B3Xnatww9XOMPEpHBO36vq8sx+nsbdo09zSXIjGyl+23LuKcYm9xSGAmronscG3jfH5BtRRPxvq
XNH7HUsU39KdlrmHDwFumYyiyIWZ7v0rYqho0iTpASLAgJjU9g5oQhWvS0tDMShpAyECE1kdBkkm
CNxTGSQ9n4JZsOdultvybZmU6mkOk2QqLudk/Z4ru63jChRS8raivhMMCSRtjikipVXrGjp5WI3Q
/lHCUrOCMTxeb4xun1iTMJJObMO7DMti9lAe8uWJkoSzcd+MAHoIrmp3bX9WXPvRvjHKLHIiS7HQ
kYsUZ+xFC1Rv61UtEeNSYiwHH6Asap5FoAJ3nxeUcB5FjraYInVKqVCobaTIdAQZ7XmKz/MZaG4r
lhLZ74/9Bqg8I/sR8gNerGC7MJhG1+/TwgL0G9Iqpg+uNNUyEFpxBBRfzkgurUaFuP2fxgBAVxzF
xG+C4Dka9x/nUYzDHzKOzYcFclDRlrTryYG43EmQoinc01jiJyy/2Dr5Wqu6uPFE3bkfmCKJ59jE
KrRh3Lqpg0kl0rr2kCvjxkuiURdR1ZFrLwnSJWzPrEZD6be/607I0fQJU/dJqphuz1ZUY/A6R6r0
siEOfjC6NpYGLLk4x0+7zjMviRJ7SLPcreMJ+/TSFmh5XMHYqY4HWnG0mjSVLlLJPEfEtLgLyGiv
VVwBaDF3Nz0lUEzm9gEZ34t2WR+Ew3YNygtc2J1mcNwamyB4X8YIIpO8van1S8EQB3nmRQqM23GZ
aPgsqhZ4FwD5LCK6IVkfCmFgIniDFQU4Qge5avKITGL2L8yZCpq/eB6hXSXHrbi48tSxeEkU4hHp
onmhGyIHV149TTkIlsGjK4dPRZuKrjDvHfrhqvgKCFn9MG5RM0ntK7StPqFQg8fAFnW7CCPYuiAb
DT8Qr4vq/AYKU07chzMjmaydfMYKxJCoT5hHPxLcfiICIBBIncPyx6bOehzlWhxRt5JBxRTZTNdX
8885SHYId5YzOzsAkkZVaGkXKcItrL5P+2TNM1OOU459g5vDLL4WzDugzeGcM6p/AD/HTYUub21K
PYd+qKJ+PxYh4fQKPSniNhZX+ofDLjZfYQA6wUUt5rpMV2hjzqqejco7SpiQpNxMPjS5ZfLY0svB
+WFfJYOVoZ0Zn28VQX3i6mGuRU1/9okuzPiue3nce9XRcFeKW6PLPZdtypSp0fpS6xa+h8GUAgqF
Y+47IVn0On6h1pd4+PD7djFKkDuG/nfs2w9M3g3aLGJo2uYq9maouyIvvpp8mYrY4jp+sXrWON/0
G8N+PIP9DlAez1PNG+5Ct4Mr1tT0VZko6OBqfpZmMA83GJNMaL+ZpjLq6Cg/YG0mtvYTYiBC8q6d
+DG1GfkQk/DOHZ8Ag1EFXJTJO0v/znIhDzsEzfS3WQRx4D/kWVoBA3ZabOR2OQVzB276KyBDu1yr
TgTuRWv6OkXLnlFTfJL//54Pi8t/sMVqwIYXVv+035QdVlGezXPxVf4EKWjVLrrj0R9LxFcjx8mN
+0bg0lCPKk0kdsdy5d/OcupBvuuBvk6rnNnQ9ybj2wUCe4t+fXySv6EWVI73CJCXnpjyuvmKzmnF
f3oL9KPq4rAAFKyg9qpeZfJ0mVu8AFxYVz7laQsfKegiEBT9jFyRcorufAKs8xuujd8/KDM9dxg4
MJ6x4fNMByB44WV+WmzRj7QbJwxsEuPPXvLg9SOBZTbDKk0F5cLvS1/FJ60meI87/dfUtlXDggBg
dbSv0pvFsU7FyNMiSWdIjF06vd8OEs9d+GRXwbaQyLvA6PGyH5jvd6RqrhW6tZL5TizSzMleosT2
eHQ3sMfhvcYc54ts7STHol4FpI9iAjodJkmcixzfDCR8Yh9ZqiuwA440BdaXioVeALlhxOVCmATA
E74eCJmxWXSLjiiv4wxr+8hgP2YV9a2JN1jgP2mW7pqKC3cwbYIqfmFl32rOEIfBhjgMPmwHfiCo
laoRxSOMs4thU78lIcbS101KNgVtKU0zFLKReZZQQIszboJ/QGm36VCyIkiDatGz+KebJF0Efb15
aX4FiYh+aeyqo5jSfFFTDm2uHx3imS/Arqbruif9nhU5D7O14SKi2uACCHcgga5tq4cMKJm4nkDz
mY9jAuf7Va7pk45ZWcvz1E4plfUhFVquWhUMAPZ33FjrU9M2aWfNY/JBYVMa8w+NOmcDeiLfzqHL
pRDMuGMSpBh06DXOIinztjfXihaeo+fdfArq1cymXASbusAgeNNOO+2K48aT6XyK/BdtbwogOq0Y
mXtVxphGQYIsNDDlYI6FlBEVOxSnNaFZbHIeQGBFz0dmblKcLRaJEN/faIIub+iaJVouQ167kZHr
ByuDD47kPEROfdY/s8xQR2/b+hDCJZlKU98OvyrKOSOKE436FvkcuGFj6UTcvi5lM8MCGi78/wh7
CcVpmiNz+FVUkW6eybbq1SJkIr3zKENaN0L0ivPX6WtXBrCg65Ec4R7e+Ni/BxJ8GO/9eAg00wet
O8tCXMl/5KoNScz7ukKqKNhR0nV6uxl87Mn5uhfSdJMeBr8sUwmM3zgkwiESez3tW2erzooTHJxT
niGmaNfDIN+W1r8hI1vAOC/+1KHenwuvrivJbxNtN+D1+GXNiP4c/y0BWanZsF9TLBY8jfDZig1v
jwG3M1u0POlVAhB6gymrHvGxgUn25oVWU+w6DOclVZUWAa4Fwk+nEwBr2bcp2nV1Vd6xk+NT+The
6eY/DSgu+fAS7jSGHq+PmymePKEQuabIqJfYbMtZaQUNAVqoIcCr0b9jrGmSN5Tl+WduyvxPFnOe
yeo9LxOtCoKjXjpIzmIwUGUNxdIv1JvgWJymgUW9inZZn2eCHuuBGke/Ooh3m0l+F6XT0LUg8WKr
qMy0V4UKCBd1EIm5jUR64Sr+hnqLqCmpZp4SYDVY9UE5auJ20xEIz5bJ3Utlr9mj4B10QZVuZ02m
/2fMYkY0fhY893vTdTlXuuv81PbDIjrX+0867E0Bpo4coHDXNatSNjVDvDpj3dL6+OqPZPNW4usc
lGm+0xEbhXgJAdAHzhU77UR9TYJ0KzQkKZqJ+WQa76cy1HGXAvRWkLnmYcjA8qQ6B8k5PGAn1MDJ
dOzrym6MJPVXmBXMsT2RbiKDtbT6G/978U9jZeZj7CEqdYlsO8lHEm1RwsruRCJjaefReeDci55T
SQkueYopI/wm8AtspolATn0P1kyALL6TP7Fzj8cnLOcNUA9nCx1F8Fp4qC7tJMYpgmjoMJyq9B6S
uLeNNJkIFVgdlqCFCb5ebZHSLIQzfAE6AM1vwVmj1pyYIPu7besZnl6uQx4q5KUmjiAOGOvehwVk
EThYZ987cXQuj3eY4TSkqG31LjnT1aLn+mpMd4qByKglOwfTJGercfdE5s5z6efH/jXXbhTkyPPS
C07eYbOR6fIhnnHEjIasvxpaAsiDqertt6aY+mRrp4Tahf2g30snnOSu/QYL3xTPMTUgcUuYIUaJ
pR9LUK22f7ud3l2f9o0zpOEB57koPvm3Cj5jqYKRTYX6Jw2cdQViJ8J3iMrtntZUuRXxEaKYQME0
0s4QV+kPENyT0pOKS4XBtmzCxn4okrOgs/TwITBwJM1vU5caZTk817uorHLEu3/yFCwv7O8H7qfq
RK542G/QbVLryFXhjzLresnI4Jhqvi7rKvKmdzcJAnsjJPnq6stw7okRv34MGRbNRiTu3uVI0Nfr
89M4RXn+70EjomT4vTrCBetNK6UVrXuzlLUlS6f897ocZhMZzUcqyewUVa+YeB12O7l6Fwvyutns
j9O3rJ7TG3/2iwYHrxffXC1ZkQYCCUFevvOIPQDOTwGNR2RQDbuqbEapLf9jMeAv6a3WVANyvqAz
y1ER0TCwPBZNTO8PZOW/IBLem3QgoTjyRl8HAg3nlxLmihzy53VC4kX8/APyKfzq9rwKRdflfGS8
Df06NL1hr1vN3e4YnZXVMDMWn89wUmmJ5shaASBscN3z2P64kKasujea25ceYzmE5+NlwviQMy8u
f36Rtrpb8P0Ckfh8JOV2s3yNqhlILE5C2b/Tr8/ocOeZ8ykoEEcvtLtuJkyWGa6xLV25zEa0ErnS
pL3nUNWvIYsscK3pi9mlcwgT0tZdZvbepp7lmNsM3YA4fz2Kue2cZ6HcnL/Q7fH9rOyhMBmcdhCv
zLgdzMFRxJHjXpG4y2iY92Fgr3hjeSrPMZpeDiJ1074tPnavA6P7uyrIqM8DXyDc2kB0fw2O0E/S
12LxFd17J3QwcYUg0Y3cHwe6CwwySCgsfp77AIlx5LTFJ5UkuUwPcAqIAca8WeYouHIq3oAl4UOy
AE/DYzWChnzGEdiDvMi3maLECqs0xiXfE+nS1/e0XTJOj3GkD5FnFfQ2TRoW+e7+eT12oxsmFx9R
Ds6A8QxRo4u/QB2H4NDqtWZaMzfkcmjWPNggCB/lfh9PPCMJsQ0BouLY6cQ6EhOKYTrQ5mkJshqE
O4hpMyVA+AiioJvUYeWTiJo7BU3BlyFO17mhZokfWRoiBchS3X8i77GL2rlnKeCIebBzmeb3f2rw
DOUX1S5zCMeKHQLHKHZK9FMymXxICW3bzJe0viacB3KzyIdFJpXUjKAIrdmAF3rRf0ILM3v2rr+D
Yh/dwxmlj7EAeSqXis4qEctNLBu3yJ/1E3l3L/mkXCUDrKo78S/Xxh4/2o1O7xfjpBZxLKccoM1x
WYiJ1NByAtbsIRMazxyEskBb6wiUAg1LVcYxH4wWi16z6mATXb0BTH02mKrCcXhlNAP25V17aHRs
RuApn2zlM+j/SCf+h/1u/g+3nBmpPQVRYtz02nMgJh6E1vI6t0ry+BBoPL4qau8oun/U527zXGUB
rSzKbeJQ5eCfEw3/aXzB0OUiwmj5xhNUcsbvTWWohxEPrsPKf8SFXfnSmV3+jD1OG54sGgDv3/2H
V3uwzLQRMqQVEl1Z3690Ssh8O0SBibt4X10GTrTHlrTPFxYqXP7ow4nTWwz5hj7o6U39Ft7PXsG0
NUF0M4uzkaDpXN/acQSNyVKBUX12kl7w/ETnkqbJh76M+G9QpuozJnE2Hik9w7XOhC8JKbPeNTJn
ga0Jpf5/GcTf0zSsgi3CWsybPkEfCHBFcKVYMpwA16OXf7oPvu/t6baP2QZBJT9YhDEg5od+jl9s
dD9QPtMNtmxb8MXI8+fSrixingxW5lQADjwI8qZTe8MmHhlZDKJDxcDYN2VcjHkZiU+13PB6tjCX
iecmPKCTjMNFKEzaCpmgXM7irHx41b0mwZsLbIb7x4fWmTwcbXIz/ujKOo9knF0vads7B7iNueyh
qHFDzKrnQfNp2MBpjZWRkYRoIDr+MM77gxyoq2k8Tk16JpvGIbUW+qeY8eVUVmzJH2ON431ZIymQ
g610h5MrblNvi/XqhzBUgJVDYIQx6dLlaMswgswZU4Pt1wdhisPQl79Ocf+vUMcD17StdlGCAGL+
3QBgJXZxbxrZybzVyudYOJTjZFjn6AimPAINZBObkIYZYxRo2GZ4HXR2x/nuJMjWlds2wWVUZ7Dp
7f2LK/Gym7b3b/CtRhDQZTHeedbewgy0p6QNkcaXepiBDTsSbOQFUb2Sm59KcuhI9YiwutwP7zIk
7r74FrQMySC2z56ihUQvCiO6kDHWtW+/cUwt4G5eKPTwFhrVPZ/lYYrRxvMkidVLZ4ByZxbdhXh1
Fm02TliHJtloZNBxs/97T56k+EiYJzofXFdrbypIIvDawYWNBOUuCG4BJRPJH8qfq9W7Mj8MsKoh
IOTVCcz6zPKpLfFXfCq0eQ7jv894QgPW20QIfMYE4j0TaipVKlB6No6e0F6a9sCc+kvLkUay1VfK
nIMZGLsSwVOMvXLCuoAJZKxPS5yctiReZaQw3eNRURVU8gnCgtAosDu6N7JNDxJAKIIK3Ur4B4pP
+oVw2FrJrXSovwpN68JxVPetliEC/1RHarcZKYThlsABpIEtlPNN5iJSI5ms1Zm3ugPkPxL8QW+T
ZMKu5pylJXBwWH5kzoZXPT8p5+BEfFXXowlc0Bw7tXSeP5EmhW1FgbxGkADE+hRJxlM5+5n+5p1+
r0Q2KHHVjsmQRKZIdjIHSvwH46OlBKmrtRhfYXqOUgL1WuttEr0zTT0m9O4Ancf0amOZ8Djk4Bys
fBIvfNRseJNDmTFcPW9BYDLbK5Lt+NFXr95VwjDdFMsSj2iz80Db+V7aUYWYPCE56Az2J4erIaZG
8J+fHun7iLiAbh0MNdqQKB8l87uQNAntyGjx1qraEwplS/eSsTo2DzIWXMVZ+jfstH9hBu/10FZp
Im4d920+5zZ76Gz4iFNohyScKjw8DJ8EgF76O10VpFQ87RL4KPmCaP9DBP/WMUF+JO2HcqHMnL4q
xyRalwqlVXgsAV1w92/GABabx20zorz4vmJQAr6lvb+5gzSBiJndOX8XI/Y6A0J+w8cnzgF+WQGh
DjdBj5nWveWb3kAb8esJV/EkZ/jJyeiGBSDml5BdMQW0+sLHgc+SvlDMwPUc9vEFPtJ4E6D8hwlP
YMj/Cnv5B7iMaIhD3mvFQ6UbbeGt1/vmK0ysVsMbrFtXXhk2xKZIg/STObqFXSLn2ypQhVEtrkFY
qrVZbULXWS89w9EmCODfUIdXyx+XzunbD4J8QX/FQlAPdyeDiHP/lme5QPtw4hJWagD+VDKZm7w6
SiuzyLim+t5CpNG6HBJQHA0P2BxOxN4H2XhrrWBoMx8eGw15Vs0jq3jtovJe8IoUW7JHw3eypK3r
m1+CKuKQwqBfMj1tUyO/st8h76U9m5S7zpU18lqyK2phfqqkV6D9Z2uLU7A37vwdQ2vvKV6ykq1K
QZ1QDPylgz52VgZHTcZG6krGL75CtCg+rd+eqiZt/F+WHgcise+RlcLQomVj0bPJIUDtaF//IVYg
Ya5TNAY0Pu86tImItkJbFuHE2b4Ku5t3MFsq4uGIgSgi3q1GCoga+RofUlWf1zIzdrbR09+iA6QM
Imcib6Xg3GtnFwpXXsfU2uCOZTsukO+kLAMnIRx2fU3l8pfiMSalvtpYDMNhJ0AnZ1nBF00oBEzH
0pNEpQdPKImwwfo9XTyyY3xA1J6Cn7q9vaOjkQ+3e0xpq4K6mH2gU2iHtJgq6U4WZqPFJGfGLDbj
qBMtSM+51V+dmvBXMpzgOnVe1siESWvJ/XBmDMs0TrK82xz10Z8f6cFGD1lDL/JvRS2yHMdHryvD
ByRvHszTcCnMcVUbvw0hNNzJNs6q/zLWU1RWAhTbPjCOfmKr3246VbgiBzFJCFqtNuN9BBvfuibM
9Ux/2AgzLsZBqf6ezdBmFwy7FDIwSMSIaWVZUbSs7+AsoyTdGU2uIgWT9KlD6XPtQsjnmvZIKpb5
cisH5osuFHyd8NqKYv3G0wPNPVjkPXohir8Dm7fU6unZgaKTo4k+HH0IEisK+NkejALEV/yrEnhT
mgH4syVyV+HLrh4egxY34UUKFBxJwnd21Wym5NuDpRAegvtd9WWBuvcwdlb/hOI+aKWs0WPpjBdJ
+8E7118kjL66Ex9MWXfM1NsE1Fzmif2NspYDw2IGN4wIZPF+uALxycDJ53TdG9FFXE6DksGJ/qZn
rnaY5998PZieWfcKAGrbuRH7Dh8GTTI53w/UCWnXY5boJBFVEhv6pCwz/6B9abZWz6VxN0n7M+i/
obolhoTAUfaTqOaU+BxbrvcMX64aqrD09sFdph1fNPH68dxvbtsRcjPAJfIOE1i62TNeiPrYi9nr
fbtrOrnSkOCTwT22EtpTQXEbiHTnTcREUeOZZBuGrIRIKAi9VgiCzgV4WroxXsMLDPWwLC6MJOmo
fSWvru25L6o5kejW5u++NiLx9R64GZzUM2rnWpNd61+O919z8/PpL4xBxdtHfhsDPdXsjSuYXWH0
kTwNtkub1dWaheEA6RdrzAvOL/TI9aUZfJv1sOrmSeIHcHYc+ZS2n9+Wwzw4lGqhOyMbDE7qIe3L
I6cwVrA8vqL4hh/Ois7RaqKXPodzDWLVdXjgREHVeni3qVtIGG3mjj9Sa2Qhxj6UlGZ0iNe0mQx/
BfQmhm13GMoiH1em0Nkx9aiGHdwVyac8AtX+2rT0lT5E12lkJQ0jn24pQcxnlFv5/VAc0m3hPQiV
kLBWmExCV6hT4DAMJrYxG1o39aS3y4vxMfwiBIPM+pmwwZVYWeEmYQvN6MEgsU9ptJ8rSAqyZF/q
qwQILUFTX33bPPp2L1N/S1i4l309W6LGGkvevacDAB1M76vVKPlOj6Eumfi0mlig6oIjEHtJE03m
SwiiBvNM4WaCc+BSh7NbvyZXc1+2p1+2cbs798VgJuH23gXGVxzf8kRrUsNS/Z7vsiAKPozwoIQX
GsFRUcxJY+xmt5jIgg3oslurWA40V3UO/ruluG0Iz4RYz2+iALqOXiYFkq4kKUy16sWt967dDvi4
kyeabyc3AaNAqHomU4kj9mgk4h+Ag5JLVJkbUcNhhaSCLwo6pBKSWrp5TUaF4RkyfLlQSMSmumVj
/QFykO5oH1u00niaqJ0Om8uvNyPPBv749Ky5Zk14SLtloODdT65EtVcN1qce5sN9OoURrsamKmwA
cseczPc+a45Zy1VSqct5MTrKluOoH9BUMBsSl4s5TOrOoZeE9ovXeXlATzgNlrRyFUwn7gakBcyj
RgFjVCL2pIEjoHX7/A5nl97ritOE/0jB2hcbc37ordDjIArV3JikQcL3nRwSv6k/2U0itbUEXdjE
rNjAbORGvUDshxJ0SMcrRgCZ/fwwLXG+YCRXA825qhNIlMwQ0k9Unvk6Ne/MDk04zJiQKjyXmEsu
A+D6lHQO+Cy5d646EUAcThUANWVPnBNY3d+SBBWPQ8Cy7GD523XzeGnd4QDS2kBoOVB//t3pDECt
3ogMIR3+1Jseyta9lSMnPsvg2WhxGzy4LTMx89jVWdbXweLBLsx7zkgnCCW8sqCCMIjhljlc+Ps+
H5cdkR85NcJpjPtP/MHgddxKe8ok7KXAYmP/Go2vnIDQ1FB1pGVvgf/CpyNmR462P4WmJeyEkPqn
u2WGa1zRchgbMttCpj0kRpRdxJTtjurr8qNW5EJaWPfe0n1m/UqUxJsovU3rjLMpyqQIDk3vxLS/
kRpRYaYFV5eJXIY2tgiDMP1DOy477GMG9yxDx/Wabpu2geQ4XzMuwt5KDSESfHam/TjczY6xmXA6
azrty9Sp7xB7qe/kgCmzQ4DEXP21tEq/IUI2eVm+LK4szAxlX64e6NVrRF8aOX8KGHgTEh54jnZM
oAN95uaIhYqGi63C9VN97OZ0a6PPsLPwaZYbHMy2jKV7c6UYtWReHmg1vqgPhSYdAST0R7rbLez6
XCrWAILRsMGiA+dkBLEG00JfpYLfNMTRIn8u7B5Zm8WDnQwrqtGpFHc/eH7+tXE/Y0w7lk9jxyiB
cs+KpiL9TAwwqIelJgZlVm+d29OY+XsefsPtROSd7fh2OJRidfUpcmBrrqGLQZLiAJixSuCHNvw/
+hpLHTrFpFRESsvJCf2o+ZDUlCRSsWJuj4Ai7oE6RlZkVJhGOkxF8KZBZXwf4DCNYopJFLKAgCUI
nnOFZGKMsTcZYQcMj9o7ydlV/7OeSLyBqR6JhI0r2EkmnsgYQV5LZjH6F8Tuk8TqehnHKR5zvV8d
DRfJwpuny/hEsz0kIDGeKjD7p9SL2N7SPoPbk0sQpUEWCpXCy9JAFyn+bSlwCeYVoDG1bHON6YN7
rf4nVE9JcArJ16yCJWJ01QxpKJoCXQXgRxGha/IKS82pwQ0cogEntmvDnT9WNUA4RpvLGn5somhH
pi37ordIxo+meOciGlfv6tYpCNO34kJ5FsxbzGB3JFtz8CqeYL7jLbSLMv2Mlvba2rxoZbQvBzPx
RF/6y0z+FPi10c3KtcRvlHQieZRT1/lfgP9uId4ln+PmNCS6FEhIO8MWZVseuJ/4rjTanU+mfIK7
P8q/wcyfIPHMhJo+pkYQjCzLmfK8qL6uW8TCfkpRfduHgizmurq63g404t4cZxA8jWM410RDarFh
MOgF1EA/qZ6gHwkK8Mr4pW6SPLBa4H19wmJUcAre/OoKQd1xV3UbTz4X+kCF1t30Cr37l5hfKJ2P
7GiULA08fzgj5CDBw59vG7KvymGypgssH8rqMH1OjSCVSp61yZliRmAs5ck8lGMrSmjN6hCNLguE
BOvkX+5qsZJKytviSEC4tsHRN8V8d/57gSTdxXcBlEGYsGqeTLy8BFmxBx/UnIu2SdSFp7pkeXv9
n7shYPHxaaxHREo2koE3fQEdpuDFTAs9JA2Z3sEAESPuS6it72PTrTudUdMjS1Tu0ocKWDk5SOAm
oMB6PbklRRrkRaRABKI3O05rBdKlQvUFpGnYVWjdgwkCISBLZMf2PkBdAmgpF35se7DbsYGxrWA4
NR5VrMGqzDxY0+ig1oZffmk053QGXtuYM/EI9Tfw/vJCXMPTYtgS/m/JwzasXJCS2/9T0NG1LYA/
hMPROtZ0bRyizEFammjN5oFjrXKs2YZlXKxoNvu+qHhpbAi5W1XtT94YA9x0DncBZZebuqvzJzwV
NQGuwaJu6v8nRgkfePSThrpNEbLA4sVQxlpl8SwC29RQ6sL9fC+0G77ipc4UD2BvddArSFm1f2+i
A0XuuFbsZjC2gTsq1NJv8YJxqPIylmkyIOLXHcf7elJzxgOG2rynUN36sPeBurOUq4zvXbSgEl+m
BKGFTbJyoNCAqdznynav1FAehlWrCDjswLqeSHK7juYsy75xc7tEmVDinZ4zHQpJ03zXBOMlRza5
kci++rrok71Ie61dYJOq6i0iaQHT1xxj5AzXdIZ7/F2aY7kfkS3J5m4kfI99OSvnH1wJTJKSvmEZ
PlYBJyl1OHwH/5QMOr0kcXQ7EwwxqspM5LsQOSzl2FD6EsJ7ahRfkUwnDGbriTpw7fCIAr+EpHYN
tn7WpWrjmmvnNjdIJb+9fdBVT863yQExySnFrfVWZGcUGZdTraV84lKxt+i/eVWfxqzerYwTJhmB
D679a/bXbtrmaNEQJYZ3Rjgy4GiQESFuGPpGnwdHS4TEV1pLCmf9i4pMa7QHP9xppX6EeLpdzVnt
ogDKh/U3K5g6nik2T9GAVM2W8ZyoCWiDsJQxH3WN+4R5kd9JuXgL4dgnkN1J8PTV6kf0zxXmdipr
mTe6Tei/q/no2IUkoFuc8p7M4ey7+7a9ItWQZXVqu0vA1hhXNt2AL+qXtDWH4gPFWuvdzPlX1YB4
4+AG1mdumMPoj8CArWQl2bK/WQss7IosmOBXba0hDyI9YH1Jwwf6JRkr2aBPwW3RCiDuDnzrlYzP
0lUjcpHqGso7to5rE/O1eX6T56a1YWWoria3V2bU+MRK8O6fFFngMxVLo2A4kCi1HG7yUVGaKQB7
4w6+mTpxdyP3Vsk5SoQno+VJCem9hoL6rEghIsgr/FicGpGCwo+Y7YZdEMtUm2R2DpCnf4HY9YBy
I0/Xqm7kQ0zb0tSi+S8VVpfbPbUsDYroeayC5TTrjfWOzHXLxTjcizseqc1ujFvVs0PZZAadlNTO
UG/ZITS2U3Ua9vJicwhiT2uMnw+Gohy6OraQF2YPr4t0vNeD+tGBMKAvZV4osM2rj9FY/hCmaBAx
NrdEWJCc1PE/+EkL178y1lcB9XwYdnSfBDa9rWp8L/xruNFW3okhwGhcT9fRW5rL3XlYUD4h8V3j
ocq5odm0NjeET4G55SjC2FyenXbnvvqRtcdCUCDj6jTZ7ZlO5Y8q/dD54Oc9nEJp+b1AbEv1OCse
NEdNe3ZUUCeue4nQs3lrdwh+ZoqZ7jn5XTJ8GbNTedVTqIFfFrhx+d3+keeUiYIiNysAntumGo0b
themZ8moroC8zszVK/jkaqrmBVjQiHEhiH1jP9m+KOoLaK6iFVmD9ilPGuNYiPgTCSZSkYxLP0ZB
0rIZNed/EAnXzaVLnHIEoKFM5pHblFBN3RZKIxHzdrxIBO6rjm0nHmUkSkmkNsleuv6uQ68eXW+J
0KfpPGmFO+3oFY8C1LmvpkdYEzcKL+LL7gpUVl43b8SLeproQn8X126Zbvufef6OYkLkkxUwFJxE
Sb0mvAZIOJmkC7+V1n3WWLyFCTfIV2GewaE3FAIxZ+OI1Zf8WHet3AotXWXBBMSAyNNs/aNG54lS
oDapSvuObnEF91GMyPxm6tRfzbR2YVuacar+7CGUhGJsKQqkcZUG9F2BOkIPAF8W1fCLE690s50J
t6MgC1M03Q0hKmKSlGowNq6QXJFYRXFGT2//Z2VwLsk+TzBO2WGjnRIa04NxSKwwQCiztlGLMVzo
6g1DM4b5ege5DkuC8YFDyy+bKJnOmy7bxJeJ22KncVYDY3f0M/L+5ygdIY0rIK5wNzy0jv1LkQXd
Wz3EMe7csTusEuO2x6cSD/e1v+gEN5Zf/NEf79USoTbnJkDk7jWI0XXw8T3DpWz3iAoKm2mLnSLb
s5/ZaLxFDTgtJck+MeAqGOKX5cRlj0cpHjlElDRIKq8lcscU8RAlsMhjmb2J3AdwIP/Rkm7vf4Az
bDRmaGl3DhHBye0fOQpsa5sSLFE//lOjBXEwtxsTlFrbqatR2D9pEWhmg3GsTqibefe6Q6TBteY1
+claVNok+YmLZfAAStDAnRcpvLR5XaGX7My9Jy6l21kgzTBVGsCgJcThGhlRX5AMysGOqWH6k6I+
zgUym1RYWN18OOCtRRef1vwVSJVJJhd8eu3zJYuZYVZ6Trx9ie7yWCDHrkb0b/3MjWxgJlfrOYHi
lOsLJJk+GynzZbmnnxAaANtrzNGi9Ep4E4KcAlS07k65IrHOjGRWj27ZeW0Doxc3CKZO2EbI/7hK
3nL8/do4v5K4pZ6zjEYE7QdyEWDPTGWeHWQJyhtqFHBvDhD4UR3F9aAJjWqTucntHxI4t8bt6JNb
T2fn1dqq+z6Y0v5q4SNUrKUdS3sHHwhaXNKx+47t/oHK/caqeejM3MCRf16oaNFEftbiL4ZDp7Uq
lEXOpc3nA1MPAcm5W6rHtluwh+Il0EfAD1eI2n8j0Rn3JLz2jL6jEZkQlA/oV9p8zijNe0BkWHZz
5slgxsZfL9tIpSoD6AXzGEKVcyMxPh7a7WF2OXE2m4YhvPe5MIHcG1mW319kDYZS1E2zp5xaCYmT
WTtKwB53jfEPyLeVcCO+b9j0VGjB78a4FLGgRqqI6dAVoNrhX7wvQ4wo/l1GKkjxUFK6TFKG1s6X
zC//jo9bcXOGJA45Fd3Aulxi7TEUGhc1/5mB/3eymg37/kJy2a30ZLmoRSpIy/ROqwmB6Zj+ZRC5
sbUwiqK4Y4R6kZofRDUEX5gnzgd141mXJqX5NQ4UJLJ8jttBJJYEDI+xJ8+0lwAZHbaW2vqIppFl
CEdLLGkliauwHie+aXorlwbecWdQbjK0PDnxBiWAUVf6+yC6dCplyagSYpOC8gpGNSIBpo9hb4MB
QTUFe4HH5Y5hmTbzc9Osa8IgYF0WKROPP3Q5/krK/wKwZfMNo5Qvnw499jIQVY2L9tt0/ANvikYv
BD04kulyoN4XhmLEfL57Def+F5lNLqOhwO5oZ45Vqs8FD+awCopb/2Y7APvvNAwKjuaFUG3pNUaS
ZBS1t1jqSJxA4jguXP5WuQY2touicZwsBy6Rg8FhWlZWYBrZiQomAYJ5JbFjCOcwsyJ0KT1Itlgc
ZfUMJMFo+IrvT11E53E9+vt87EBGXObKlOBmKPboKvu6JAm4MgWWWW364LC9yRqyuaQ38lo9wQLb
DBO/gsa3WuSos0e6bZQcvdWoDwHibnhe7PsVVhDY4qjTd3dNeQ4kTR22kr6+ycg4+I+SzUkmgG7R
/4Ku2q+J25DFr7PjQBuafkonXv0a6TwJW8msb5SdhQY5uugPBsO4OS89DcNvC2Bn7FJKt0BhUZV9
nmQZ2f53yBTEfNY2iRl6C++Xm+x5U/5P5MW3BP2QkqcXhLfjq9+qv/obpseaiXEJ/0cUoVC5mM6n
O5ySYHymccboccJ0kSWbui8pnkk7U+cSE30CWg/RWIu9WNma5kVcJz6vuUBvUNFwHWrqtpZ1zgqe
7Mkq46DYUkXm+NncfIpcOusTcpxuzVJfydC12kc9YhTWbKYDtxMt41pZsm2TjekP28aqf4InUTII
ShPhc2vB/YiyBRlwa8kEqHQj9mSWwj0GiP40Sxnu9SSffaijKA+Ik4/pENBTJNGXG6dnEH1P2HWq
Lnw1CZ4G/0XtrzUn5TZWjM+gs+ICF7yBZjr25kYGF0U7e67/ke+Hx3ytZB/lk35Kr7jXDRE0/zxq
mdUs+L3A2jNt7i8ygkukcBNsPs9CJuuA7slTsoxtzB6qgFq1GT9dBEuEqQC6pkrkz4141G+7Rk9p
Pub1aJpmXaBpmvNcGgwkGGCFlFsJM0QbOLA/t/bwlaiDCXKF19dgbbfQ5d4G6rI3l0Cz86QCxVcw
Qby9Elx4rid7/6uULTrFv07vdRSz8HFpMFgR4VC2aybCOhW1XimkynYb29tSPCrdT+pmQccaTXlZ
sjKJ3HOoIR06U3DPfcmkytKlpdX67pfjyZH7U98oN/G+Ie8OBufdZTkjS8JUH/KHa/CUUDh7s6Xp
CpyO/Dv5MWACKDdJpGZkjieF0xNYa4FGPZjtUW63z7Rdm0KX76fRam8hIgZvOBb3vSdLc32tLo5X
Jdo0HRCZy3wWmNGabSYNVDnsXDlmGDUHkH+bl5JD277MGI24byCVHuj7EvO5FGrAqItilFbDdg0I
Wy/RrVG2hUDBXZMpr/DES1YfyYBQpzeai79hFXTpJBdp6Mq3lwpgYiutnEkGwz+sgvpbvqvKGLE2
IHY1+Jp0zNMUDRL5CjPFbB5B7P6omPqw7VKkkGoRwsO30CPrufExIWsxRtjxpRrSGSCcu2mLVVUM
GyHhiHM3C7G5FoUiVkbjjgXBQ8EfiqRPM0zQcqgzS1slFQ7VkNMx9PjY3RhwZ1KhWSimHAfKHAut
xo2h8rJTULlVQP6Jxj6R/kixELIVwwSJ0EDsGJQa6UzuXy93mB/xffZjLbEFn2FMPBn50y+dk+Y9
WL43tVL7MfbGayIIVvh03q5g/FIRZsYW5UAjgEy8zcNC7vY8hxHR8RO/emzkLBcCz78u46hixuvO
3X2LCycN+vLUMIScsF8rdHytypO03LA13jaTM1dwLFAlsPH7+YwwWK/sAjWCBon1rpPSx3yILqXi
KUO4iuQzWJBzborIqosS56oyHzrJ+TtEvs3CpQwPN4i2Bt+UuD2xiAKuEGQ9NU9F3eQ7hM8PzIPN
eReBybcrLOuGabFPRbFxSZSkUkG7YWU+OiUV3AwBsi1ZRm4LIJ21aFPKvshcD3PzZFeUHchMq/yc
Zq7dZJ8tvg10K1vZgch4up2NQKavM3kU4TRTieo5bIpx60f14XL4jrvlSiY/B931wKdNNXz9Q3fN
rNZQrsGTCz8AXOyQiCXyNLoFcadSHNZxcXabjpjSJQfPfSL4CtH1GHnOor2exPK3Q/e8lFtZKl5d
LCd9JMHOor6R+Ie9Cr8bl4jf5H4ejYBSbbnKG5stttpDvHRQk9xCWEB7FoqiVE+JYgqqfvHx7IKw
VVMOUIedTpAqmP9mUSLMJOJ6m4nIePzvc8VxpFZ9FY9pSkNf1LhQFNWFeJEINpmWwhIbPz0km5bZ
3R38nhLpoIe8xBT1I9622eDo82YcUlGatwt5oXijEuKPAslO5KWfM5sF9/tuOdDXR4s1EqPECvHs
vQxkM2XL52CxyqiECPBJz928xVPygZXuBm1ki0h5g8iw82oLSyReatAOG5FSU7HabAyZkSSFf8eD
/lXTcGCmBJ+3ehVzxOoY+8hlzC+nIVA01u+n/iGpeYtCFgSHFYYRZM67G6RmtA5/tCgO5y9UGPHz
qbVJ5SQ8ktqimaMiGBsgAA6H9apmji1Y/bi1XewxwtCtfBjRWLSonc2pg2k0JchgQOwumzw9joXE
AvNdMbj3NO+mkpILkhTioA9qVEW9GyWBN9QXjFSgcPoTGsY9mfUFda39I4GPyJUjkwAayFk8ihYx
RR1u5+48OkpZ3j9UNnUK2oyRoBGFhAvDo3JtC5XQzb4i2rhIRoFoZvCiL0boGcvmxh9KhKaY9pmZ
fFhmiljwGP6sMeftSI96uzTqkxHfa+18CreKGibupQJYgNxNjJlda2LP0JpcFRXHDrIfdLR5MnD+
8WuK0y8inrveOEXRe4bz3Oiva+GVvQuqtZ4dP5Xn01/dbi2msVYLm2/mEN5b4YEV5b16FDrt48Fc
jYunxXt2fQVG46JGhcBsxw4RdA4OM+5bTwJ5YbLfrqn6vPVfJ8eYwPTipDtBWVugJOHuUEz0JDUT
tpoF3zb2YACtMqj381nVpupiVZfoBip42Jpi9XqAHYFTIKT/Fao6W7MBKdgl3EY2DgCCHu8uVqeY
anVOQvcIQ3rmvoCCKw3RkSV0MYz295wnpxQje9UL/+RTQI32qqXrlLgFov8QnttRYDdSt3hyXR05
v4fpcut0u1bQqyvu6lwFIxQixybnC1kHwvSuC/K+cNAfxhHRoFW2YY9fjUSX0cbqQJCxV+DsOCZX
URbGLQ6M8/4IpSiu9AmXLqSwsbZDNDGy44fu1fVwliyRDWsJCnLNiVd5WZ37NwtMA3r06xhLssGV
NWl1TlP8pPTpim5c+GLtSMeUTJOzit0Bfa8tDS0PO35aaNmRqAFAUKntgvVwYwhsJuU/A1uTFBJu
yoz6cNvfatApPTLKAXRVSAA2ZUW7FgFZ7toh+RQg4Z0eVT+abW4QmrLSXmVVEX900okyHZAx+je0
NowM+tJOLDB2gBRnkiwz18V7tW7RxNH/Dsf3yYG/qEPOXxL/p8IrLrSjnwm91fcteEErL6hq45gp
VWJX6mbMMcyThK+GWZKtXVu3vLSA+pnvpqkKLVftS99OXabgKWVt2J6VXhxa0AU2rHUqWJa4WPtO
AOp4ACgwhj5rDAhhniSw5y4/A9j09KhUjAt7XeJT0k0ry137hfUeIw09xhcDKCA1+bTtSTIOYGK8
CHVDctBipsfc5VvmiIR0rNSGq1lNPrRYqJyj82lbIP078Mphc7XeD9a1YaRqc0ZzvqlQAqm2gwl4
bdfkGWk9rU/481d2dIhEzs8m3snVb/eXEyMN2F5Nocq5fDG+kKDYR95nn6nMQiAeAn8fiqIEVPDB
7qvFt7Maw65feIr+w5scEiJFSL7P760OViTHVuXTRdyRgPo9t5PrUIYY5kc/LbO+LHXOGDdYPuX2
46TkbS2AtCuxjXEYn8R3XX7L1avwHbJbiTC4bGe5M27G1JzBRTq8krZ3OFHbAazToxAso7Qap5AO
+8V1IFxZYTohv1WdrmTm3HLQDHMYs9ALNm43iEqpoF2POLuep69KeStT4iVZcLuHzFOaHaOfFINY
wdWgSpldv7bGkBusvR6qHdR+5bb6WVFJ2I3MNK6IG5Eb96/kdAln5pzijKz+sdHTAnQ8kRiUajnF
Jl5IcSwBtpOs0jL1xO4zm4ahuj0rP3OsOa8XuZ2RSPhfoznNq+K0zC1ssEusDD6upvJhSPamoCPc
JsihUnWQSVcyHTiyGOYAxbghegO/8A4h16AAoho6ctaRj8N7QdCfI80XPUDC2cWDLXV6pSdGvEIP
jdp7W8zBB4XPphXpZVsCfZi8/P1qRaovIWuSS+PV7TUAuLvDgheQjSGvjdVy4xWyl+FBHA59aDQT
V+5qfxqJm2rAb8xDh5sB9htcEZIilB+1f8AWBlvU9Okap2xtMucLhyDOE1SwpMMdm/dAG1puFahc
himBFejSM/Jkp+hMmQlDpBFINqfdC8DXuiVkTDB1CtGK42P8PwmfeeObuyzspm3ex/yhzEfbi4CR
R+Dv1mLAdZ04fQ0hl+x5bYcpqdubmeQFpwGavrk0m71Ik/Iq8DhczL7mmSjZTEVeDz6Q7g/gllzN
eI0tRjx+nzSMggw45pE/x4kZOIstdB3a4lfeXaL/hvuQeDwNSdoazYQyGA4fGhYLZN/qRZkYy2rO
eD/QeVoF0d6wn1avRgWQ7mtrqx6K1qqC+BDAjyJCFOqVdvZRjyHLofU74cHwbWzqcdwanpZ6/i7t
1WTCZCmHsHhknzdGT6EM5IUUeGj3BN012M5EnUQgpa+/pqUqePkEo3ukue91Bu3/xUZAeiC2ZauT
hvxSWde5Ll6MkDHkx16ljY9+Khfg2KyIg3VmIfW0hDpWakFAPkqP97SHSD1p50JMdwRX3KegHbM1
q2kAwE5C3ihihzuT2os4+l7EoQflWcS6mQi7h1/dJaJGyYCJL955u3Jmt49eV/COlgiKplbatkWG
pgk7Z4HwT40+w99h2vPgdubrZCLhjAPcJXXIdy8EVMsETXVMA29pNwVi0Z2xt0WE0zG3Oms1a2SF
pnPDFNcHckQ7pD4yk/sBxTJTlF1XH4M3ZDazZwlGCZPvRs7NQ9YZMS85s/rmoj1mXrSoP5xK8kFj
ccZ5XdpOImGvmlyf5AZlpgGQtfj3aN6Bp542UBGunOcZTlYempH33kl0w1jMLb9vzmkIIOtXyIfX
D0XJJ+kg7rxh/g194maaao2V1+VB03jrtsT1QpyMRsSQiiczyx1Q8itd6rnuIkqD7ozP24VCuCsh
F6JFta6ytEEfeEAEEn+MiPiQ33ZV4orI5E5hr0Xx1tsSKRVMdn2+XS7ZvoRcBV13Y3P91B+tWdP9
gkOoymnY8g3t+rMUHYnbLZpBsvWwB37DMFgzWkcBoAY48J9o4RudWQeWem/a22SoaksrWP7t8ozO
r1HvugP13JFhLA0EPunI31VgtUzi/17Vqwcowcowmh9Rokr1Cqrc5qS6Na851wQIrx91rbBskQyY
s4Kqi8JYfqEAVIGiTMSsryXtzSD7G+kXgQtGL/LM7BRiuRkL5U7O6lpaOW6KZfptS0AZ4mXKXTwU
KPL/r0Toio1rnjNogr1EzTGOG1OE8bwJe+QwT+h6a7G+wB6if9aysdIQ0xsK95+gEQAa+cKWP7qW
aF2ymgNWaQzfUkYCWF5+F3M2KspUXrqX0qgD3TQHzbiZItwU4oGmNBwisKM8BX8TS8nO/b7mMFye
qio0gmNzaZ99hWO/to5A4l2ZYXSMvirzeLN+omeqJslX4sDntMdxGGM+Kfo5fPuA2bSIcX6OBmCk
0QDe7BYOpeR4aRjMxNmSzkC8u9lc9gFGAyxAW4h9aI51KZ4ed4pVvcZWI7RMWr4tSFpPHksCt11N
k1KF1y4C4EqOysf4MvDh0CMCYq9yxJzLo8/h4VPO/eF13Eggj7+Jo5CsO+xOdJMVxNUHeFSgYx/T
HAe/K8OL107kid6lcL4ypgORDaNviAlbQfdSp30Edpsom5cFIMi6wi7t/N+TpAopwS25UymyL+mU
D6P2GfvvbQT/oo3F6R8HtpW70ELWDj5X/OcLoXl3huI2x6k4lLo3RLSWJ9XANCHmOenTeTxsE/AV
4C1/bxj6VHC+nLpLp3PgnNL0GMksxG+zhpnb4s08cRUTfR8Z5hulc7U3xwpgewsV3hxCOOdfZJ1X
U5pmtrrXdkzKwKMxJAqisiH7A4HhO9Pl5dTa36dqdyfBxldfROCkQbyiYu3OeSAXx54TUSqTxrgg
UETDIMpsX3at0TBoxM4JyN5a/vWUPrTMiGtOQDgt9bXXPzhobvfbpBUm+9EDpSDRa1iYMpy5QVND
U6Necw2H4lJPFGU3D9wQPzWCpRdppTIYl08xQlRR1ZdFAc2PAj3UpxOmBH0U8rpFFk7mcHpnXN8z
h3bZd8pkHDQh7PqjdB4YWl6mV+C4mf+fwb87xDQPvM0NMOvxzM93qC6p9yhqkNWQASGNBG7+XXEr
pKWC8IVQW1em72NPPszp3Fpgf1LfIFvgVLLciOy5iZK9deK7PyZMxF9OQVurxldgrciAe2BCKpqx
bExbolwwuq8BKASSLppRneyjAaVDiBAdFhAInjJ1o8fzKghhGe0og213+kyPk8DnZTrco8uI+1EH
kK880luhXoeZxb/3+DZFYz7WwEPy5St7NZ7sRNNwudR00fgl1gcPmnEHPqdhX1WE80/7ELpAomyl
+3P49tnvQMPkxxyjbH2IKQg+Nk4eml/iW5riTqcN/MWumn9y/Mf/5MVGjU6TnAYbQ3+2NZzJIITE
fVmyS+daWKoX/pfjlJ5ha2NthMRPnSZO1P8+hE/LYJuvdrr386vjVUKXGF0lch1NTTLpU+RvAMus
c6PIQQ3BTOGCXtwW2igvOnbVL5tHxPib88IhWcns3zmQ3Q6OV1Dao44QVxH15elQUgGOJguj/fRN
/28dg1VzgiR5vhFxjxJ4sSV7BEcCxWmfcJ7RgTtvfyl5cxeqI8NGKfNZK6CiB3pzlF82vViiJIdh
LJKVzkiB8AE+z4KE8JMssp/DmTL9G4C7eP9WQhNFlB8hQBZcuyIK95YIwQhV9qYm5Q7J9MKcK5+o
Y2JZZcfeXjOPxlogALOFEfYYZ4aG6EbGVt7/cLtEGllZoInM2VfEMsHRdLgx8rMe+wb0Us79WYyg
WQqfu471pd26Yvfl09UUCM0tCHLVNYRNgK2srjB+liCtfZiMxi0/CHuHZtpAA7iiORlyj90/ssaj
kHOalUHpKVEvZUtzmTtTF2tLhI3im7IXpmiX0hFiOVo9yrCQYp6XypxNvPo2J94+S92NPW8dnDmb
vcrhP82kbIQaXYpOlI40P979rr7n34q4wmKkyPoJpQCvEPb33o16mpUM2uT1ASCBuS0pkSmpJp+v
bGodD7GXbSPm3mTq1BkAOUub07N9ti7rRYdV6o24SqVYRHBe5IeAYg0kiBFvlddSlYYK5vZmI64U
QRixwMUW0VMfqX4zf8NrauqAvBJJrLGAjVVJTfh2YKjAGzpcqi6F9Uzmh9qWxnLmiDaYVeS1Q/Gz
C357hQYqpynkVTjRQkjn06IS7mf+wOgBk7G8oz6EZI+0nGiec03I2HGHyGGRmWEy/QgU+GPNKWhe
7hf3JSPByXgDYH+4fbDWX9mhZyBJUJ3TGMIFojiRRbijgTghilRQxkkhfSZc/+eU8wH94meaBbQT
mlIHNBMchvkTLaeUjA54TJ9TvH9mp9oIEqbaWulFv29aAkeryp92fTdY+t7LdakGxoSw3aOEBJwh
MMabEwWucxG23JlfB5ceM1+87Cq1aV20RQcLHpRpYjXxQciU0V9pCTWsaixQsqcT6hcoCnchmA6J
2k1fg/5SBMqndM1dL9MwkekyXVRX5wb6YDIyVnWjff+oPKxnL7oAFit2bpOU0etwe0EIFGvDXfGo
k51QuwAYxRh/9kW4dHIU7tOmYmRWxeXXJd4jG4Z4vk1uF0okAy5OAzEgZOnzW6srKvlqKGbRe5sf
/sq1/DYJucwqIrnH7bFj6zMgrexHwykNDXaK0JWd9h+AYE6SUhQtGPyb4aImiXkV0CAOHicOxMS5
g9P4PsKPUm2g7a684s0qSW1PKIDLXyY4tSqjMgri+NJ3pZKS/CKGY59i24O4DsaDtqNFD+TVZsdF
AQYjAya3m6VFeYwjgWaXIzy6mcUtVYJYwb1ogr6yvZ65slZp+EMgb4XVuVagyRdLdmsGP5Ts1pb9
9bBx3J+WFyninOujMJbPCkYubKwObhJCkW/7WGG6OabL4eiRDQoPwocJHIMSlwkckC0/UQGElsxs
rs+WEzkNiNKuM7kLZ/0479UiyGliurn0DQN551lEzuPDfFrb3KM7Gi9wuur2wimzdM7mD5p6Cqx9
Ud7rAT+GsGnbdl/P//oNWK6/Tl3ibZOU83yFgiMV7MjIkKTbjCr9Bb36gJV6Hy574Nqg+Dx2V4m5
ei/U52My2mvTZIDW1Y0lyUCCu1XaR9gKO6zAq2yIX/sBMQl41n/cS3z8c0wKNpX1W08T0daTNySR
TBCFH78uvOSWWSQ9DuTrWZYVA15zwH7pjsHRAOEVsiiVxYs8B0Su1Ma6oBxVXg6vcT5ZxTywaMA1
qM318X/Q1AemHxpSVSs+L7bPasm5SC+UU6Bwn0VKgAaNmJEIIQT5kzhff9I0WL/utYSJAQSH/Y4a
EoG4ruZAcDsWIEqJC8ed5/P2MDYS1UZeH9R3u23zq9uZPlnoBuKDBoiO6S3rjthbXOgeAy2LyV4r
Ho0dIZDK8tTZimYuQ3q4h4ybtVf3e7GhlIcNR+zapWxBVFEWGoouNdwKZfP1r5KaDFM7ItVwbH4m
/JknSyG9Oyo50gXXIQN4O/nAx2vYsSLLs/922cRlvVpmsBmmIlU/CIIyD9nKkgnxdxN1IDmVhLBU
WjyKe4iAKA5OfUPvfrhxnh9ydoNQo3oEaoHxzQPNZOfEpz4T8ZQ91pWWxGm5dZvS7j1ItxLQ9nUF
YrN0bPcTVBRadrTL3E625XA1tj4Pltpl0IdsNfQkMS6WcKO4FNdOTjRmTlWIKhhp32tIXWNx5HIo
TyCdQehUivw3ywhgXA0Ky3DmaXkw5yvH209nALcGcKWh6zCmuo+uyauYtABbeBzj981/LG9JJuuv
G/O1JEbX8641D2TOhU5JDzc3OzPIkD3s4IGkoYai4jF3Y+AU/rX5EUr3nX+jIcASFsmePNlH8Le9
5zTJd60znUwfSn+RhWcgl9uAW89LJNpcXiC87Vc6mA6M4tz4Wl0ZRQ5rPcQIKfPJqkagVEV8eXxP
UNoL8N6fv4BlBcyPSyDoBBN4T8seGcDGBa9QQcCGpQ6i3kALkwUY4nmBRsXthAT25pjGuFVd6zSk
qrOdP+B/B2uaWDEt/65H3qh+5duGgv8UgV6nGkqbCelKSj/2QFGq3X5/sdohmoFfz69eN9pY+gwd
qhxZFUkqSnfykz0bVWr8IP3KBYE9UpFanAImw08evJDU2Xnv/8EO2CwtDvl2Kv22JczJDpnpXwtY
F3zDfLn20MFmVVALGX3fcVzDiJJrpfM2H+jnTs0wsKv0MCHq3psNIAl0jSMVA0/jcAZFj4HnXm6t
nmju0TYMsEfLYu+oDLJ/yGEJYG+SM/4XyzqZiiEwnmKSauq5iP9qkPOXUy+y8O6IegQYfdLQGrkL
Hl6gJmJoqw5H9NAf0K3xgAxSsz6M0nMwNaTWXprp2xrvkKR6PN/vvQ/yDS0MNjQYzgxSqnoyWIgA
pNhj+QQJQA8Gee7YSm/roBw3/DX/ktylGkU8DOaYAgCIwlX6ELGJPTxE26gQFslVmTO92oVYUcUQ
F7c4AyrbvkbWVKAYrNg8O7Xu0ro1fD1rJYjZjWUa0LX1ozJyjdrhGbrGL2IJ/hbG6hucKF7L9qqC
KuBeG3sBxF+pTuXuZM6H+Fl82BFcZHRxJoatithLJ/d7ytD4BBVrp7AwAkqrdwAzys1RKvJRa3mC
gKlx4cwN662ptHS48IfSfChmDD2QoXDFu0Sqx5sxOBG12LdkgO8hkZJVRKCGErEzLVdmd6ety6+D
l6wnzm8G+hzGxW/zrND8e/RSDKLCEs2RvfgNyoV4sJdwKImHcyC2vc9dz5v/8AvMPSuEmRQgc5so
/t1auKP0x/IY8DvMCLn6ICiRV7y9H6aCUdboshE7HOcYipjoY8K3G4NcMmtP6HNDW04dnnMBuMiY
8pYxOH9L7Vz0KUhc06XNT8efQht4JILWFUl6VnDz4wI5J+xilEMDbTuU8ZZd9Te2jb58IS7zzqj0
pA+1VqbLjnExYP5SKm58AIFpcFqhCvccaJCr70nkhhPgLlQRVwFPHu/z79gack5/gwzkKFpG3Bnb
yO4xj3T1xm2KDu02ByWSMnLYjgT6myqO6fN260L6nGTVH82Qp/MXVu+E734suMfSLz/ntqBeZVo5
37pLuMziQSTLXyDUIAeediIxa235F88oAO1F25MylGkneN7ICtahN+aWZa7io4uL/u+a3C68Keeb
lmKyHvv4y0bqPOnsqlKZncH95DvzAIJU7w/+t6lxHdvoKH7jZnO/y4Hmz7+aJ1Pze3/Y3EOp6KjK
1xQAAI3511ahGNQxgAGRwhcizDlSWgUf5Oye24F6m1aNr8Zk6ytVle5/6MEdg5H6hP9S9z3jV85s
2iw2OexP90pZKMXvnMTcoJOL7Aopvjop8WBniW0zmsYG03nkPEtcJ9leTxkjnAyypdZ7GVsz4PPd
HFqIhAja74Eg1lwW9GH5ZjB0+6cFLF5UheDLyvB2mXbaLkxph/94c/tRBkHalmTEhpNrdcyzCsiJ
G8cW5b4H4LsGPChrHSruOEb7QusB5BzIsvnfqhn0LftAqIUWeqPtcErPY6KYpfQFI32hNRrvg5tm
yx1t21DNeYWljEaFbjGuEPMywDWD67dFTXhaMETwt2hmtNQY9Ph9EYsgUFbP/w4qSpBmKLtCCXZP
k8cmhdapBwz4w5At7gYOlI5Kxs/SwIpW476JJLMoIB/oDanm99ckbOn1sxEDC7S2s4anu//1nt2L
NnHIqeAQKRBbkVRXycwR8sDYroBt5sfMKjyrGa5LL1rjPYkW4RZaTDYfDyT7FTmmDks/+gPclFkR
C9KQKm5iyjdJToIxYy+s30ISvaQBKhZwzgsl7I0G75dhWMxZ5ZLxjbpBfBEA12O8g8ZwJ0F4AtGs
Fkbg+Qw5z9zBoGJwtroAUVPnSePRtlrFa0KXCbj8WLSgRSaiil3m8Lbdi/TYnKF4ZNeHBZcy7SZa
AwxnX2WWOIXXcKyOsu10CGQu1L8L3kWs39ne9COgwG0QjJQLD8eK9ti7EqgR1L0CSKQckww96bmK
vn8l6FGV1YopXzguHjtegiflngItwkyzkGVWn0P66oOA17B4G94CMxcHBPJV3PtjxLUUdM0q306m
8S3X1bGGpSAp1QJ0jt26AbpnfIBB1poNvtTR4DHBstLBgacAO2yVIParMgY//zlPYC4LbblE/16t
cqVYdU8NGpCSVAd2ixX/xA+S9ixVdO0Gve18kkX3Xy5R+oambi0RKYAA261Ym9WbTNbYaQaoh5oJ
D83BGzwdRs0RbWBdkGTJ2aLBGL3tlZNc9KgBAKoYLp+tpL/5tbkAj0LEt/BVlkLmQTIsg+ajXBt1
kKjFvcG78nX9YDuEY3YEJujl/IEL2UDbMSDOY23ddj3cmmnDFXGiFrofVA7vJEDt0fzpzMQZqpBM
otC5tNxCee0He0+tEMsULarxofufdOIAuXVwkRyIuJwn1XFgHDntZ/86dpGviBg8rEqHGAXYvoh3
Ddb7oJwP3vy5uanjyowK/GltxdF71ypZRpJ+fr94D9hQyoQMz650OY6S9HSY9a94w69hFgJY+q9e
Ekiu8KWxeeiD4qPgoRb0Bo7vNnYaN8JN1lwxljOgf76S1NFNN+Z0zQQjum9+kT5KDJxzEDXENfdV
7tG10X4evyCVODGjOyNQsm4w+ZYkcY7kOvuaaK14LMi1qzsdyCZUZUO8OMt1p6yGVW3aNAsSFp4z
yJiEr7/pygC2NZj+2rf3N0TRNdy7glwtbNwbrGFFDPsKNuzFTriz1rnWeLrt62fuJH20QHfrq+av
Qewb2fN2stW7wqp/5qMmWyIjm38B5f+u4nqAZrW+GqCXw84L7DDMX8D22jEjtjPOu2so7GktVHuE
XGTjOX4s/eGD/o+0tahPaF55L9h025VUdqKZLYRid2nYmJLCLCS5fjNcULk2VE2rFop6QbARgzF2
Y8Bcz3eI2HvFk608oNzlvQEZC7KrPY5Z8O7vqGq/Ng9XRjd8nNB27iI/JqcSEDrpE7NhP+QhsvhR
5WECAHqNN4w8sy/e7f5V1gmF8kU4CLUimRWDncxlAcDSJ7ZElX9YBDHpQEhyyeYv9YHB10FRzJNL
bTZoLfxamGRmIIDxkvDImWtDbDKSIh9diUkVXch09F33FaBpOXURGcd3yfabr8Bklzjvh/FpWqlm
GKsDi6MaqGgsr0Jfh7yJ+eHsZUj5F8SVYx+vnSI90WDOEgzhuTCHnb90/u4BCTyF+AzRXo5CPGrN
pk4G1Ja1plDMCg/MASlU4FOGVWWHBaw4qxzGwukJSCfPhyCdtNgJmpOBKExvsING4p4mqZx+mhL0
D7DDe/CU4/RFD9bghBX4UPUhbjSsDW9TSeBUbiv+iiLLgyJO3u17sAOBf1ts/oe4WDsFrlc4GdIB
/5wI4bG6BHG00oYlVWokT4PgvlObTIcLqbzFO6qtXwhPiVNfXlV4MxLO7NCTYlvcNt/nIlR2kpSS
xZkH4qV7zdBHDTZtV6TEKUDQV4j3JX6JK6fCJxOScvnaB6q41z3w+nEGMSoYx9x6EPnv+QsmA5Ot
ZZbOdTHAxc3GqBi8KPH4+IhW0yCP0SlAYyyh6nO7gWIlT/3fwCpQUayFqtHL+EhQQO/s2c+0Fw5s
RPtuYYmIUP5dyAx35WW6W2m6bNjqBlDvH9AJAzlBSdoL+nhHIItXYfphQ9fFN59Krng1DZGcYQnI
2OSGlBEwUnOV8GLRDfGnUiNo2cuwl7C4wLHTaO4evyutCpNiUDFtsJ3ZJYBpkAzqOMXI5BNSEIpw
YMftyVJXPrMch+NBS5Mu7QlCfRQY9KVJ1ick6BVef3zLaAnWuV9Ktx9Qh8yvy57lv9bINyH2LEeq
Hxy6D4O9+jY3VjTKq5q62gLdTLImsEa4APHCexpeNojjiMcnTHvBk18O9or3GK4A1t5TAKjS7wdh
OIL7PEYWKQocuzHovZhoSYlGHabiiaiiruvkVuq6OXju5MDQm2tF5cxAIGKTYKGx4jYNrdJQygYa
bfwxaKalGHj/WDCGZC5B7DGSPXL4WmyuRC0Vl8HaJJSw7h9xsB6OnvoEwEVaaNssIY29bgJewWaf
e+Jn99qKQ31OQqyejHKF3b6tNQqxb7nkyrgxhcmuOddMc80bk3F3hR7QF8VSEd8Ak1QSxeNzHXSd
FujPzVhJbyjkG0CMPe18vIDvDgrhsUSKw+oG0AaEuYt0TqlP0vrxGA/cheliLwk3flhluxDckBCf
ljwA1YuFLQjXfXH9rihqJU9HlePMU4eHeV9I7FZU/XvNcrQE8Jm7e6qJRIjfAply31/JmXjJ0ggj
nzeAUtLREBBPOa2OvokKMzqFluHpx69h403SCwaYcRhCvSK2wWJtyKEZBq6voPQ2hc5MpsUqJlHH
Z66lIw9XWsrCn5yoSGJFc4f/kF2pn2RSHillOCM+gvbb5Y5VA1U2spOZ/mkL9vZU0K/77zvcgzcc
A/NHLlLSlWucig0Cdg52Gs9ZRq2xCACAAUCfs/7VJ+GdMI2kMNixzU5+Ap10LWBmxFxy4d7OxupO
HRqSz97xLtBsuqBzKPcskKmilBdrD5EwRQHktt2NQJB5XVssEdkzymNc0uarZdeZfElL+BxQbCHU
opF3g6UpzromGgIxsx6kebZHiVJUX8ij+7aqla4bybOCRgTr+A/ulvAGqis3stXOw+dQoeitI04J
VMMjhlx/xxhevX2Iatbt8+X9WYzGyUh82sa47KRyuOQQEWOd2S+LHTgcE9ut3fLiyU8IHjIgjA1x
/xCmEatNyjYYaiPRr8OIKW9VNkvgm/RAB1dX7ZO4POTKsnmgqjOmdFLpW6ZPLSyf3a247SqALJ1P
jZ5ymwkDSm4qWw1JvDuav4/BpZ54dJn8s7cKo9VOLcdjLx9fBk8ZsdilgSYvSCTMGA3fe4pgKees
tB8UwhsYBs6SWUkui6NT5hK2mR33R7DdBiRwQxsnis6rpMcMo9nry4UWSHO8bOnTwsved8Qqw3rv
4w6j2jCg7bTJk4Z5FtyjUwo0WunNrHrGBvIjurMimgXGIWBni9eW9NHBFfvMOLL7PeJlqEA69w9P
qItSY1pNDk4B8pY4XBCZhQBUh2vlOYfzYst73SL32JlLmCqnvMGoGUC03IunOOZ2SLLT3ZJ4n/hI
HMEK2Nkio9apuErNQyVgEcAOLTk9FS5oDrtm3mBYWd6XdCr1n37Xb45zSyD9YZNwmSlVQAdSGDqB
BPexdzzflg+Fd15wFmLYkMawv73HtlMB/wJypa/oe/DkXOeijXdF+wFAPzRzzawBV2UTIR7v89py
fF1ifeFbjHOl+4Mj9H3Pvl0a0GWtRdEzz1SOH8Akmi2Hi6MqoYoSEcEOv4R2MOKNyseEYxy/lNpR
96i0x1UnZnN1/wGJUo3z5agTesjq4Gbb78PTDYKMyvRXDciy/y35l+ZH0RjiQInYJ+bpku5E7zWh
uOjdYNQpK3kbcqhWvuNFmH3IELAPz0I/+DCE0Ik9FGmmcfVfl7lomwS5LS/jlFJVzsuCzw9otdx6
VxTcJ6EINx+CRuOfJbkLivuRi+8U94pbprF9Im8fJ0Jmw78PnpDW4R5AFBhiKcjtYzMI3gItXQ9x
f+1s9C/pnK9v2fJro6RGg7cvv6Ij/ateeyiJFhJj6DUnm0EZ9zJt7rCqcPxXMdr/U3ZcLdyP+Zcp
RssjbDtcypdIInFkEnpgAxWnwdYQiiSqwYHClPRQgES9d2B985zx1X3neaSEIHIGrrQDXxXmv2N3
4SaR6+SK9y2F/YdgUY9T0bB7LZwZ3GxweMQwAigve2/eK/I7K1e8e9GmT7/7TTaa5mLDY4XXUFtp
mNwPaZGSCUPEz3LeV+qCIE0EuBj68EFHJl0/oYbLu2xjuLBdKDwCncfJ+ijNFm4j+ZRONGLTOWDx
51U6fqsImaW8ChHij3+43qWE164EEdfz7V0N9HTP3q54IyToStzQjx+nXuPclAH0/HafgVC9m03m
c1vUinc+vBhDnzU5o8+oo6D99+U0CUdJtcX2VxGl6c0Q7+fpCG/NnPGQYZAagveHRdgia3NYeJ7f
2TCO4eTys9mp2yx0wRSkS6y9bPLU4nwkmy+bly9IvBXTRDDjRJ7FVMmkt4uj11yWsZ5qarj7/1a/
eQ2vhXp07Oi8/VF3PR4/MNGNqsqm6amdpDl9lzxQwTrdtlAipChDwM8KPtxHZNbiJjS/AlyNF1UO
4cnJ0aU9bYnkg4IEAqN9myBBgNXlML9ODTDtCly5aHe9SlNUy/VbI/Lp+LL/Ldy8MCO4dbIhy33h
wKz7MJE3gZmJ0oyG+fDT2Vvr1OEgAAaE0aQOgl41IxJCP4d1pGhUJlKjKN1dmvIb3zZuBAUaqbLb
ZkHHBgvsALKUlEqOF4HUtILd1pyTl4n287Sv0eXP1QuP5e2Nq5lb7zR2aXGRd7VSNNGtYN7Ewn2M
y+PQsnWPRSKYRMfyD1DHeESiyX6zQsr6KrQS7DmaMO01MR1nM3VBZiYVzKMoBCIQkmHitEaWssef
5kuvMh7cc83cuGUmRp8zcu//V8TRousySON+5pBYnyNdj3mee5dIbeqyuWk81z9FDj6DMkDXbHiy
YQGv7S8U8iMXYvxFQGJHJKd6HY1LUBPHCrsL6QDk+0HEAY2erd4FlhOxDGD11vmqLZSbS5DSkkfl
FX6/I4XAloZbaV8rR10FFkCldvQpUGmFBUPzX+FgQ2Lqw38A7LAwe6FTc/AnOc6jHnOywBtncO6a
Md9p8VNR0ecIX+TbUBbA+obdmBfFApqydhtXDLZ3tYxzpRaaVGx/u0uMNm8Qrbnx/q6VoltnFHtl
Huay5JVSvJU40rEJTK91A+AANBqhjKoPtEV7OYy6C2KrT3DFl8mqfVJMQzEjnrc1QMlyKFAZ5POg
hdCPY8Kaz5UFdyaZf0zUWKjbDfDcQQNwkgASZwAH10aPQbYcMXzgSMlGkZGz5OwP2rAN8hBmOQIk
w60m8SD6tgkfjDGGf/qdWIotfPRviHUQLQxqeFjf/732yQxpImxbW5kcnBGIUXg5lMa6qRp8jDmz
x5Y4EYvXBO3Ix0Z7b9EONFkwi3IJ6fdqiA1Vo/yv5hB2okCtwHK0sEBh6YFMnkEb1YQVO2wJ64J5
mYU+wf79JZTKT3TLxC+SJqX2wi7eFL7x+FbogLMJhoQ66XJ9hnciOku+JIN8JPNGVWFwMy8WYaF9
BflRTiWwU9yQ/M17n9PWzkXJAWipUA7lGMQUpaE0XiKFtkbOrnRWiYmCuPfALpGNpNHj2r2RpS+d
eiQX+HLwvhROmEuVezIeQJ5guDSZVwZtVSMRqhQ5n19qZxD8CVK6KZtNxE4x0t/MGl8hYVUY3m39
79RyVJ+gMLrsxzx3364RrrGAIjqHu0YH1+DJH/XnKu4jaS1kynwfIZIo2m5fvkQW+XH3z4JHgOs8
SH1t/G8gypBGOz8Qcsm/g32FIS1BjtUvaOQJmsR4WdUcPxgRhwRKYm5V4HRVAO1FHaDsIRebkk7R
uagFoUYv5LA98COHZXXiYgNCWGF4rQ9AWxtpyji2W0EwToigHoMHo99aI7j/aTp7PTpZf4epaIi7
s4ChcQzAQXpREX+CFmf0QonQ3YYTnMaoGS2l35Qtbqo41Yq2STy4XljQZxloBXpT+qjyFtvThjaZ
5MxQGgfCxUyaE/l1JsUe6XcrtnYFUzwmoeEB4AyAE/Evc11qH1tFFUW/7DzBaIEikf/7ig7ZobaO
l3h42jpsjXynMjc6u3MKtDd1gBqgrYgCsw2K38fB/gYTS2Si7F1RW8+1UN03ZTLCmc2yHelRUXDU
Mn0GkFCPxNZPH6uCNanfwuKcxWCT6Ju0DyztW+soUyiEEUgMZnUTgmeLMFICsTPaVFuRnifQkyz1
JIE22SuMrnuhwTAuJnUCkX9Qk4S1AYHOS0zYu48Xpo6kR+OTvY/OxKa7MAQPg4e9z0GyIAFOB4oi
/XMDeG1HuKXxRDx3i5pOXeUQ64aawx9d70PdsNkwxhgeOOV1Jz8qOAQkAAqfSHjj4vp/ajy0nanV
/TCmAakQfGd/yDIAjrpRab+Vwh5aIF8BCNhA6rEDGk7SGo5V1ZvXoZVFw8X2zas4lHynvBzaC+fR
pgipcJTleXb+ueHncZLc4Y5bWv8r1vfMiMgo2YJs8L7ZMgPXsC2r5qN3VgZyETHypYhckO6i4RcK
wgaclnxw1j85S891Ddf27ghV5GrZcneDTR3B5kDu1k6UGrdzVppImgBTAoj16oVK4cG9aq5zEL88
jk14P0gNpqOK1GCRd63I1MJLjwKUbVNhPu0NH79XOKQX/nM+k1DzOWbT1cPecyXUuEpyv/+/jp25
a7hitMXFbQ/ZEnE8tY2V7v9HGlb/zihE29qOd1FBs8ZOO61ztJsT4AqOh/5DHKyMr0ZPJlxJ0RvP
68BeT64ZXI3XX8eS4KoPvbIHIRPKTiT3YhZPyQ4U2cixcIg4hlagVPCcwd6J1qjCddY3dSM3XHcN
Eb/xYJ12uq0a2jnYMEFGv1xLlAIxiYumG5e2PMqfVTdpZyRlvflk6RPKh+2hyLvRk7YbKQM7uVnd
LAWr0cLAhmVx+75C+YZlVIRvdP4F1TygBTO/hxh1NJPL4W4/etUlQENAHwF3NbA+ofZIovkME3jD
K9+cVaUeEFSby1CHZRV914PtLPjSm5mZ+O0uBBK+aUcYeZr7qDeZ8QO5M/FxSJztei2/V2n1oPip
i5cpR1lxo/XmpdV16AJi6DktSYtgrc00BPPYRzuDwq1BuxiUjU6IfxaE756T5mStP+QW8e/kZN27
RwdzET4nqqsuFbkShYbAi3kjz/rcVc84vkGjuepBEDqrHLFX4tKZXnZCyCmnMLRi3qVtfLQkWjW8
hO94ZhC42EjszXibfV83BjFfSmjv+xPV8pFEaKEAXxobemM1VJlvcnh2U87Qr7rFXDjRjJ6wdMpd
ETdfZX3DLj9qO3OoOhkM2VTv7sMc7bcXg6pxRS0P0LYEMo85CVARzAHpMcY7AKV5Y3O7FETNKIxe
pVIAmd64QRCu88OgG1OPI8a+WaKsDM82NCo8OykYKGjKb3UqQuRGYywtUG5cGEeWsc/WXYOSjbr+
IgWWAYsBIYPXUK2/efdL0OKxTtVzZATTczKlzGQ0SrO//UJovBO3bXCQT39x7C45ZCoyxwPRTxy4
DCPnidjf0/UW29eHQ+TFxrPt4fq+j9yiUqZMSHqWUtJW5JhpAqZV1c0EJ48JMycjYibe69nrjgic
Q/81dy8RoUfP1GVoy44szRMKcJ/4G4oeRU8iwUKFAapic5oPmI835K4fxsgQYEpP1m8gRZMAu/iZ
66Rt3Q/iqs4yLFHoJchmALVFVq25/gotwpvDsJBFhjK7JRftbcBfAJaWwDB1MzvXnzXm9YlYu5y7
c7rPWGXDaqnX0Pj8oRXLBjhHhFlX7NNGKFtVz1XGR/1j7MIGYzxryKNO3KzKFpQZt2G8SHX/8TbB
xFukdHevd7hdEicsCMqDgIsYcn/THBvRwgzttDqnzG8TOMQHUxdLVxBbkrcwvNxobY8oDvvTBAU/
fwRcbiDsMUtPLlxTDoLJ85LNYMVjVMqgPd2Y7SP7qMrsaTeRUFBtuWwkFHrAPn41ZfpymIoKWFxR
4gbFCGZo/OlFBF/rz8iU1/lCdPs3QRdX0OGrgSD4i1hIudnEppx5jacmnPvxvFHR+aL5EN3ik9Uv
qX5GtNfca4w1cvZ1EeH5suflEly6aHV80p9U3VFowth7zHNWJ/M1z5eDPXzGrqe0/Dct6y+VnrVK
8laOZDoX4yKjbxvYL0+iapiJmxJxc7YXkWNHFpbfOclhXI0ctvxRBvEKnPTl4ckI1t6KA7H9Bps4
fUIfhC2/TWTaNa018ZBrqZ+xT72pT3hNVHfhDQvEHsbqWi3JqlzRsAKsQCZiminfnXlyQQmOuIFe
IVYNnaAwdWBsXV1ZU2kvBRSFtRy2W7DbGrO2LxQmH7IyJGLTWkiMW+WojEcTyYnEt3WcTQJcdmlp
kEWkinbHSy4KtReVTmhr+6kcsllYtRAV9AK6zBud4NqTpBzzaaI6XQzLnPV0T+AAJygxO6CQ9CZb
6dpS99kj51c0voqBkOQNKRJSq3B9dx8+Iy6LNq0mdlahghlRXO8xM8SWy+a29spkqCpFDeTljNr9
dXE7zTgj8PBoZMnontVuHILmelq9j0Gnv33P2YanBVi8kXuZJehuxnqsWjVpnAx7AMs5uxC/JTnJ
vfe1F3C6eG2+WJWtZXfk8gPsS3GvhIDl3kohvgnT8zEvXDV9Nhgs4RVrCS6SXzYD4/ar94/+RGcU
/YhuxSMl+UkBnqqwRYPsXRy4+DZMlU7OQ8kSntUOOHQ6aFHZB6GmdPjsRcDfMszGOOMfZTDQSoke
R3/WAMDvueaSrS4PFOALMzemOSFJb/uVP8JEJkMdjQ3m2G5klknmA8idHmbIkOTLt+1tiVbbMwSX
klundR6o51XjD6uqGH8QvjrGx2zTBLsrAJFHDKwwrxYoE16wxxo4BSIZxkk4fZ4gAxs+ZRQEAHfy
rubUxCdVM1AhYqCPCLdwcPx4xeNLXKuvTUI/zRREhnvuA96pqjYs9ocMYhSEHoZidQUgEARs2WG0
zuBcrawhOZTt7GTePvbMrkg9GAwZbQZLqdrBqcSfAtVovH2f2/Pfjk35GiyXyak8bTRzxyVyAYBd
dmbIsYq5JBSzXbkmDRslVzCjovT+4mxcxikOL2l0M7tIMkRpEepMkCbzKkPJeZLr/IQXZkbtZ+dU
ZHQgxFd5f1q8h2q41nT6fCF+JxCkXww5H/0rSXW6usSVsGORVT1kiUkFA06v+6Ic4HL1JTKchPj2
YJWiFxNwZ5wV0w8i9vCcNunLDKyFjfiUV99PgQvl0+2NrJ54RAanGCh3Q+IHappldE+f9mj6RwWk
8W4Q3EUkZMRlVd4XAt7QGScVdWZPqYTFDTEV2vtRzTcFs/AC/XIqMtMf4Fbx5SsDAIT33UGRJdVI
PbaP3STqPIZxWexn1n5X9uBr7GOJEBM2tc6AtrzHQY1Gzze+uY9IDl0s3J8bnZBocIP6VxdwyqI+
RNUq77dP7qXRlT7vlcH0zEPtiHfyS4irRftZgtZKRAANrBdWUmoij5WQtBqxnFtxrU8g1gHniirv
/3Yep7E5eD+H34mHlQuz4fXPNN11N7wW9FzU6RYRSa3GpMEBN3fXoUcb1H2HmV5BW80oTMsIFq6U
hKu5S+40a25codd6zOfqm+eLoKgoeOoSqiucR330hk00tykYFRZD6fqh9c1ePiOjvcYj7r00DwFF
4pUTV4YazPu33W6ZpP1N2IKR4XHW64Ro2rOLRJp/dDficP1NLlH42ioX2QIEXmoEODVmLgECEsik
NX7SaQ7Tboi8vKOEiI4d8iQIHXCY5Evi/B51F1g1+cH/z6Vj5jwkIVTTr6Pok5zUEZXMTeU23/0C
xHhlNEGKweDK5EOfVAl9g4Um9kS34aFm0Nv6kybdYLBER1xL965JwSpO7fv3m05yjQMeaTDt+zA6
u5kbIb7WDFPjnIdcoHqgK8E46d6XlEgnhpWrnjp3kbYdeRTISWVaUaCabraZFm1FTfU881Z1KyiX
wF+fnZ0ehTaTa0l7BttBQnUtLp99oqMUxxOR0Ty5Rnf3i0vVKHoSvHGWI2GKdq4zDkmLsxNKNVPJ
C67uR7AU13AwZUr+vkuBWU7Z/IpGLN8QF8s5l2uuCfIXstqF2/fMX3LaA9cPC1lBJadSvcXVyVWl
YQ4m2HWJrwkfk4/sLWliGEk52ZgfznvzVJ07XqHoamHKNUIRLaYNhexI2J+9urRkKLkVLtjM6hz9
pRcugQpXieqsJBFiNLDggscEYuCRoDrL7WloU7xZlZVNb0wBF5PdLs1X1Cf8/1bFOdCI9zkmVxvd
69fVfraknbdY0KTJE1DS6BtkrcUeMSGFRS6QRIKQycDyCOzrD8MbgVMVkN4WloExKpZIXlkbGY1r
e4ZRt1Aoz4b6XlCnUcigPCLfVeJ+RnzXFWBN36WumHA/4tdbohhjb4ldoTLI9Cn55ntsOZ/6fr2H
yR3SB6luhWpFiNQANEK0/+ZREysDBsrpd9zX2SIUKpHR8egwt86qF8Fj4UhZ/IVyokIcWYv2kl6C
003eVks07wwIwR+Tqvg56vypSjUHBnOGHq3p8A7ypYApj1zEu1wnDeByd8zhS3OfvAAOANXbD0gy
gucsf+5ni15LS2FkA+Outn+xhxuiLkR4dlo2YhpwQlkaeM06vsCOt72VpS500nw1OUCKdprVhnxc
4qQGODbZ5Ygdw0im/BrS+Iq0x12k8wtVsuolj/goyDQdrUSBsp9eBvusTptRsl2r9xjEdzSs/gtB
jVHeLtTXpq8BS+GQIRr1Y6I/zwowMjX4ddv0AjRB4D08PJy0PtDA4ggEOnle3KFm2oRIA2EVj17K
v5T3NA5AcPPSSXWee/cd8IahJCy6zJmUU4zV4BGAiEyOdmqSUuI1ltv3aL6KXMW2CmRqIIjDBWDR
J6GACMpM6bCnwlBBHkk2DUGhYLCnAimQaaddpC9q7gjRW9ABhD7gJxyq0OylYk5UVTFWP1PhEfCe
Zqv2I7BlGmfeGKvGGL39POKOcW9bU9FYfhqBfKUt1AmQPsI/Lgv4B76o0Qzl7najAN/Xsq8VZwri
7p0cq7BUrFcMdqnDP5p6MUsFUw9EOZqnBa12g5BCYO6OmHzvIwMd3Uom+lP7+2oh8wMP7YT2pfKt
0S8xDNC0oE7COhrCMSKsVRd3uGArnOqsnfiBUj32PvBB5Hp/gjoCzFfh2qkFnlTVLIZ40JJboaHI
zvCrst6T+haJ0k9N6Wkj1jdHFeVqbv4jwcQ5QXD1Zsq2bxRVByo+hE81zFtRuSuQm+34Y61Rhk/K
F/V1f2p1SS0dp+ZG4qTmINsK0wrgAWptunCAJaGVmPFzkT7RyyNKuczMIM3a8Kt6sfUmPWUdG0uJ
8LxBFabjGSYtxj1h9flqJbm8sUPH0CifblJIbOXWeLDZhHC1umnh7XssJWwcD1k7T13+q8FY630v
TC1684Fc87h4IhGJBgwdyJVYAog19P/bVSXMHDfs3u89V1ia8EhsHIvl7A1h08EzaOpBZOlfC9iP
8yPRmtLSBWzRZ4ls0r6XO0yJd/mG1SVHHGr/rD/hGPmUZZBc3XlMQDF+wdf1u3HHp0wktsufMVbA
dBQhNMgmtAmYOEPiMMuBKmVEWjtuSVjhSkRXUW2QzxzUYxDQfu1/Nzfbx6QVNwPVb7EbVLLv8Sd/
WCbLmVO2yxbezsthP2WMC3+ZTFlxl0TpD+kogbzKXC16PxMUzkit4ta1hCqUDW1ZtWMQ7EQPb54s
p9COA91hi/VhktDNeio0Vo7Ez9O1sbv+A8JllwqNnC07TydohlzOx+WeKuNQ97RLDwyj+XmjNNAa
VZdL+e1jBDXz3ksoUODXnSrKq9WQGQILkmF2oR/V55AQyZ1UOw0eDnh+6v/TmZqSpIRhgxt/L9eP
pnNQ+0cRlqwRpSxLgUcsAICegz3uhbu4fTSCEkaBPnlevl+xmodB1cpBkQ4KsRyvfidjuoLIf8ft
FuE+lgODIOK61iFphlry4wHtYneitcCOV7dXJ+utw02+nCZHOBjeLvFnDEunW4TtRUVH2br/wlNQ
oGxGUL3IvLSa2R1iQYRGnOkrtn5m1LmauHAPsOfU2mAsVKemE1DUTQtiXTJrh++fF/vsESHYxHe6
at69CMxgV5L6UWLzwCnrli5KJOh7Wpmgfa+BH7HBIvXSpFxlWKVZA9hVPuM786uVAWZpMhcPRtuS
3nTRYOIUI9PWpXaaf4rs0A9dXt1TV67+uJFKWFS7G5Is/LzZ2CcLwcIkRywNaYoSkvnKPrS+JUTc
sDeeqPP9EVGzhqsMBV1NIfPJXsYd7uB/q0zRdfa9IyZeY5Ksw48UGjqSmKchqwQfHgmo8e3OW315
RaJ94QGFwFbZyu+cyQCxWhsS3CnB7SSu1n8KWL3j9nKtfSjjfb3n/UwTkllSQsNKIX/0JIT0t6WO
lh9UxukpjpqTwsbelbvuy6/QpYwI/EBmYh1bxoKrGY/12ZuSnutPgG5w0N7l2CEFnky1q/d5M39L
pPCOhMuHvMZMqNaczQgHQVxc5if2uIBnCh7azhlWMspi9RdBWuCzSc2noRG9TSKvvJfr7AcL3KXC
QKkhocTwtzIMapNpDQhvQdLXy6QOI/e+mq+B2++KrjUGrn27MhyPPCJJauLMHcrKhwnoMeUYnlzz
0G6PMn1AOJ59GTHqXaGf+ksjJPDe0qx6NJs3rf4pLRXm97puC0K0jlDbanwmZD3SP/uAedIG8DHO
XGgUa2pvKngzzdfEYPBuWUI0e93wPnw+o6I5KxO0vcfR0nKOi/G4uJ9iPdI3FirR9SZzHQ+gOQBa
GNNIlyrNYXjltVhnlN24v/yEb66OvNQ+zN5kTezJr6OtoCtDd3jaiuaiKJJZa+5u3M+1ReBh9q6M
fYdEWr9jstpOEEzoTzkwp7kYJ/ST83Zf9EH0/4DlUUat+jSAGPdyrtUyZ7Y4uY5yHi3JuaovLKET
nguy8mg2c+cIumXfKpKUyigHh06vv9c8OUVyUOlAjA7z2tetw0tkgvkTmwlHHby4+qHa4OpxXwEi
fFHKVyXbpcBWbB8lgf529Maglzrc1rOBTzDo5lzkKWniZvw0XQOODJGyMmg//6n00Taw80R7gtT3
1iiy840tiCWl67njlzEjI0bkGMajvyejp8/5aFEI2//9zs6p/nF+eRfY/d9+aN1bPLjRyqx2EHTY
Cz7TcPlZ+1EZ2xSZYIN7ECSBvhwvVLMuATKgp8OD+EDILg4X8PKq665Kmm/wcpwtiBSIvefbm8KD
KQPVKuATlxC59IC1y584hEvBT2lr8nhfqnsyZTiF8xsr6LCajFCBk3+ZsYRDjLY69CEacLmdvs4a
SlGbOLXF+cAvHzocYKnXTksSO8FVRJQsBGIht/lqEbPDhGkhLyjCAZx+xBlIIxYELrjc/Y2lzQss
a+hO4QSH+BjUw/KeJFnSNHDAnIk027F9wl2I2EhZ0kxFT1FGycsGH7Gkx73ytr2qI/dnUho8JmeX
o8idM3FyfKioOCAbamCeqqC7TKSFYHTo/Ftpupe/m8YhX9v2tKn06RQkTKkOdNCg1VA4rYQjm3ro
pKOQ0tifN6ER0mKAKh+9pAHj38R+6SOq8o+vZB4ha+kbQqhKYMTszdqiNoZzQyy228Z60ves5L7C
vPNzkC3AuXQ51RIc3iOloINAmgk4I43iSCCuBOCPA/Yqq6sCyCxvbeS3S1tK3ob6nD3r5mBLaQ6n
MZ7y2Gx9o9isDjX20m+6Slv36Uvwd/5EgklOw7uJOY8lYCnGJSn3C9dw1VoV9liIAYSmtICpOPng
6s+S9EEOvylfo/UtPAMgcR5sVOrhzpKJ6/ehV96pqiZehXjlJUPKf87MKnwRhcWOxKtzbXFCuIf/
kNr4x4X5DJRzzGHC71JubeQIyWlahSmMzgt3vo+NpP9lQOKmySAeeDPH+YizhnAOtT/r9U0qB1mL
A25xFzr9neCZ1eL36ogIQkwrM9Z0RwfNf0vWM5QCobo0fHH9ycUlCY+HZ0ihMUA1c9xNQ6Xhv1r6
38Vg/egw/9+S3cJPtjfDssPgrJznnfxuOteARxtxGyQpDELNgWyETKf5jKRYziFfy9HnmwcoL9xi
LCpys2TU1pdA036GjNSzNT/lI4TWLUpLOxVEy59K0xQB3BivaAUUCThvrRgjkikO2j9IiHEF2yB2
+ohH2SdUdAUXEXSxPh8CP9El71wApBieP2jEW6bub39NFo5m6vThSTSZeOjcgowGEa3YLxODp7yR
rVUBgpv3ttfNLazj/oZX1RU48ZxdYXXFY4mOC2PI1QLr0vLtJFZZavFQJuVebtW7otLQUPD2buT6
C3Mh8KCyGB2nXv90DAiystC4LyXxBDYu2UFxiPZXbthZXbB6SigDN0wxbcfpVDsNqDvbuPdbaiaI
mbEven6i11oGrzYNsZXxOLgAkTQVLf5lf4cxQaFznpouCUx+3AB8nqiF3bTTZy5SZb6Wv3wihhd6
+lmGGMs6HjBER5PNtNEDwmIoLYv+fzAHM14beDqGxI2YdIT9oNSnISewB6v20xgIgfjEcettHOTr
XxR4gp3HDMAcnWkZRnAzJxybWvKfIU7fQdFmbGJUWngkUdJccUkEuv/RTrWXLtp6YHZ3WZL2jmOV
eXH/QomfXL/onP3Bj9Bp64lT8QMT9RWEkpZdavVz5EnFV1V/V0SYBVuSYYkzS82b9dbMStsGiDuz
DdAV9nY5tC5gXUdKFiaTgBjE9mF6fJGRW9/72Hrj9wu1xRGK02qthpdsCZRuUUk0pBIZpbdCXgKy
gr0EYh8QjH35BBJ7RXK1HbEfjkZ4aRPhXftjNUc75l/WkGqlKkbTPfbVxIqOjjI+8YDKzI0GO4ST
rt6gjI6kpLuVPR4mKR9VGczE3xIGhK+/gt5MqPah9zn+HtYgpMU/fK1+++kUUKR8H0S2oHnzD6ZC
sg9F2RVQgkoX2UATtj0Dy2WZmYhJdgZlYdRO5imeLahHLZLhruNxZ13ZOjGmBtvlHvzLLDaee354
po33I5AboHMFhx6e14+p0wJXc8oCUWaBgJnwRYtuL1ASpGakf9zjDly1e6VzttU7+0UVkzXWwIZS
2DNSgr1DWFzwUMeezfOIPAMr7kCW3BodLgUdtxMEB+DpsnPMKMeN7E6slAqjKJh69+R7cGJMHC7j
Yp7bYT7h6+LFn+aLRFY/zNHZJ77fPj41P4LCM5/w/WNo7dYwRey0PU6iPVyBJXHtPua79l1EX5En
geJLACYjwUqFaIkH+nKpmztviwYyefpc1fnvuWpUQMi7W14QL7qTC/83+sVYQHIK+rG0NNW8H2wF
P/OHUmkBzGiO4Z13e8BDcYJEZF0WQZdeHanJdxWOzR4Er4Wh0KhAmlMhqCbVgdNR16G1OYVJwECG
jiO+rcva07Ld/N9ALtGTlDRF38BBFCKavx+Dalx0+15l6CcWs0gA1wIVq3YOXZdilJx5RJ+pUrMx
9b5SsTTdgpF2Vimp1buDXv4wNXbrP/de1Lc34tTY84pLSsSdvsze81unSdNN43KiR8qBeSXyeu0X
0M6JLZLpHYariaS96cXM/RfC6CZARoirU0BN1q+/0WU9Z3eNO7TqW465dFEf2tNi9/v7zLLgIPO0
U1egzTDYWdQ/0h83vWA/Nvlu/At86uosL4Uiws3Ya/Hey9g6f8mbE4aZnwbYtOFrdS53tretFW5b
UJyGbcd38nhknf0IdibbeIrvQ8mLm7awY9aw/zhjPslMHLRZGXBeSVd3cDdI6uFGVOJGT22FzYFY
o69uzQtqejir0PxpiZBHP6P2u5n3Q3UmEtEW4kd8zh77FHUUwkwvL30t7O2GmgoLoWOLeJRwZl9R
mg+TrRmDF8qTIgX2yWvFmjd4qKNm/whY5Bo/CIyoPsVmrTVt6x9Rog8XCqpdfIBJgcOPx0kn2Q4y
uarkZNk3r1GKnAw4aX69RXYCPa80D/0YUM72WKQjM+9prhw4VCakQqLvOMI890ffGaqY7zs4veZz
lDFXmMh6bJSE+NyZHqRwA8WxidEcoy9D0PG3G6M7JzC2oXOsEPw43F04HVv7DprDtbQHqQoHtcMW
AxuHgNT48mvkRpB5bofiXNRTwdu+tYcXk7HG10F3XmBzFJtrPBsE7EbdoQyEE8Slhn2yYGS6QJWx
NIQHKv/7vqw0kYmqd/Qe0PJrzxAaWCRJ2p4dI8GQVTCQeR38AivyoVrvVEutXSMngA1OocjknRqb
78zFsOmijqE0xvF/HyIdcpQtTZCpBk8F6PZf+WRoUHJdjqNWp/nblziz7sWqkalcP+h+qeLg34yJ
XFL/kpHT8o0BjTRqVH/j96OBOGY9/m4xD4lXRAzufFz5dQvLCnde3wgIXd3WuuNpw0M6YsoDGwIh
SPGw/0LT2BKEaiPzWgAbWLVKpUVs9eGkH6PEskAFyUtz33sVSJ5LKnkOUhgpP+oASc+Fv0Zx9PZr
HOzHBjLMMKXCQnSKBO6nY1lPx1gBXoyRLRCsF+3sdPZp35NZgJ4/HiwLe2xkxYksn7EYDCXDjk3i
FPJL3Mf8fA6wh6jxjRS6QJFpv4fxtk9BEgoQW38hleHsbkaetqCHUCYGZPzyWzZ7hDRriHqphsS8
pzguj43GZvzugin7wfDHo7CpuG0R9+8EAEXZBS636tuVh3cKZQTv3a6HOtaarIgJtlDhCWw/03q9
eE6kZDPG/5+dpwQSFWpvp6iLTLZO95bXl8VJFp2wa3LS/+I74Sl26hDzc+0WqKSSvmrkskDYb5EE
r27zTm1DpjSuGKJZFmIpr7jtLpLszBwbok5vgABoyQaykusHs7EKWrlmZy9Ioq9NsDLAjzlQSyy+
f9IzKxzsmY/oqCkDJTmX1Pomkk4eSV5AdAA/wO7m5+P0nkFi6lpPMmUtE9Z7uASM4S26/4B00mku
2oRuZIdmrt5nuP2T3yJYhD0mCAKZb1wkP+CNaGR86AIoJcqH7BECt7WCzRbKIHU8Q3SctU1PWy3Q
UcKXoHlb6ZHZIEeMbLWjjLaAYLhWF7xaZ/fOjRHOZI8Uyjl4zhY3omSfhEmBjTS3maHGGSufIgbs
NOg47Q/HYvOy3BTDkzXPQIWdJVw4OKY4ztCE8cqwwAb5qtEhDWhFvzEVDn5gLfokrenj4WfPkE06
TaDQDLehCnesLIPOxz33of9utbUsSEDZ+AvIu4EjMZN7jwva93vOqH/H0Ip7AGIXACG5P5ASt0A9
unyjDdsLvhSwmLMqdrzp0wfTTyI3/I1HJEmy8K7EBZaKs4NIir7Pn2N0qrcQYPrwv4eDQOCxFM9k
w5mGtxi6CfDWvJGYBKTi+5SvTJ5Cikc2Z34YvtTG7YXFRkVgNm47cpKaQg4jjqa06WhimadZ4z8h
FC5DNZdTPMuk2wHQa8+r5YtcizcT0+iaXwpgeRi7WmDpDpjiKU/NKASBGy/4gK7sG5mgGWuZmdrD
Ci360Fj/tlq4gwi1x8ktlQdgNGy3YkzlQMA6RDqmK2tSX0ynaSGiUI9tVzu1ESobzsmVXaHyyiPZ
Ros31GIQYolCo4/AKB8ASYndRQKi2ECcliUZKkG3Lar6h+6VcipeJn7akZb28NTDFoq0KKsfvw6P
xhRgMCDEIuztVUoXjJLOitu8+UyLWGXo7BlANDaMe/+mJ/8u6QhhoeRAW8w2ageJPT4aIeOY1T48
ysgThTJFCTzpMJ4dVrzrCIfSciZ0fgwZjlSkPn1l8kGQnsQLfBkzzSTBxIUE02fPDBY48MijMXpf
NFpiHiFaPfNKkU/W8D/HE8SIfRPgW87KsjT1krNFLq1CON4/cUs85E0jmbrUxITv+IjfFhrpXV9K
gqPWHd2lNpn7fDqE+YMxmdogu6mMq56+8K933oX0kWr0Aj3OKacEVyN+f4fddKB00Orl7E+HFe3O
UaOqDhBUIYcKP14l/gq9bc4MxsX7h4/TRTgKFRy3xMzcwR9jPDEUceAM2LToz6Kyt/DNpZ1xWuk5
1/f0gu8Gl6/a/Hk9GWINYihlkNgSKg8PEDXIUagnNfSDwWst4Ra0+bIZqoOJ9bhOhRxBgW6d4G7q
ES8vF+ZcDhg5+tOIeZ7nMWo0ccnUFNWafa2n2qe7K2pHGy3kq6HlicY2JPHrGV8zaPXtuCJZamzf
eRe2k6o25hrRVJZChRf5kgf+nxKU2GPLf9Se+xY0ODwFQJ5M9fNnYXx2tlTYoPjavahQw0OcKGIn
lHaMLZ+Nl/Qi9kPyemfKDoiQTVhrINxZjic0O9J9RVvDEWT+pMoypt6PrIi3xNWd7/lnfy+IuVNq
Aapys7xPPMnpMh1Yffg7TTUOT/BMZevOzRPVzEe8KxNWZSI5mGqkXc+jY8uszHDyuJwQegq0Kdnv
KVx14g6EAj7/WtnRgTkdMsRmYrfqPb9W3QWr4IzLWhGPbj2ZW2JOXfoWU7z15nvkwl+ZnHjsLiDH
xSE1/cliOv68qztOZtn5T8nXMb8yAeTI5UoN8cHmRKwlLuubQ8Wpw8f8JazvJqS0x1gfArDmzxGS
S+HZDZjzmZS3MiVsbfrIo+P6TBMK6giUXuJcUfPJ0akK3svY2uMbdE5WrZUP0P2+Yfk2mPobwyUO
zCNgsQ3LmIce6T2pYsZxgoZeY5ergzJT1wdztL/pK4sGvWG2y9LEEn+Yh1ty7ovBdb3fR01aoyJq
tA0ubsNAbda0/8PywQLO3zmgQaIq5R2qqYU8F988i+QnWc2T8HFDdZ+LJ4C3nUVVtddi/vTInerX
Q/JGKl+485AvkJq5fVXV74oogDXDR5EmltrK1uEWVO0IotleI38IC6omsIHNg6GGA/fs8LZ2LEJ9
sjaepelI/i69VI6r9B7tGcypyOWjFgO57mqkzvhVLxHGh8GXkianUmaqB23nxKUOhI/ygcjzwf3D
TwjYQVnWAj+iTvb8yqNi7lYqurdSWg2Mw8q/2irqRbpJdPupvoCkSX+4hav8NiXaI14bIwgK25uI
I10froDJk2aPPqy5Ep38pyBinC3xt6tGFQdjj/0a5rZP0FAig5ZuKZwIJte3W30wzDeVs0XI+R9N
S9E7nj+JC7qDME06A8+j8oGnfZY27HIa5N/rhvEoq1g358wr9El674huo7O2qqBBidNK26muVAVa
KZMLdNHWpZUW8OOMDrzwGTcTBTlFe7gR1jP8pyveo5Qdwxx1cJgbyMB7WRQBDL/fTm0dbEDu9Nsi
lGY9LGXyexAXqUUWeUOx02h/KW0coFi4BFHEba2B8qx81J6W+Btha7+Lpuoc65Dm0nZ63gr6dHP8
XxsVkLacrI+h7ytVfTA5NtWmWPYRrX+0bJRvRnEr1Y7UR76wqkYp+CwchwUPurNpELK9ckBViFgQ
WNL0EcQHJTfTsdAL9QIN38NOU65d2LL3xRcOgqNgYWITQzXmivt2Iq3vX3W1AxWF5NvU7N1pUaid
nmtIcmZnU5ld2P4zYkzMXiCDuUoFGjJmCZElsPX9xnTm6HpgcHc/hxwCAGkBMIs97Po5d+7LHkCO
EW6aknY8rSLSSvuTXbz1GCVxuvWmSFDe2hO87B7sFZPjwF2d/dOp1tYiy5Cvx9XV2CQzMDf7QKB/
HbfdJdpgajR61BzoiDB6EeXA8whz0OcAYqiMriDgLzauqJEUiav7kjLgiNSCOctbl4dc2yjvOf0l
AuZIXmRDphnBpkAqCSphZyGz++OssF1eAjvRlCRWY8DQ0dnFG67SydONpwZkb4t4s+N9UliHmOnH
mWN3QIMkmmcH/SvlHvdNTJb9xK8rRTl2ezt0QPrw/c7PrkgGW1WKNmqNf+IUAwdnTXrNLv/R0Bfw
8RQSaQN6S+nm2ZC6VCRaKAK4FJNZw6GYp+ZET+RdWOY6EFa4rlJhSrncHGpYAyxLibtnmuzFjHkP
hvKa3WZKS9+2WeoLeeRtJQKvuef6CXC7ylIsRd0/sKxWT5RFeKnG8OAGak8Ded3WPVKEWdX376d2
BwdcpXbNBTgpVZCKOyZgF8ghbui6lRoF1u6zwzdGUyEqoW5iW0LxUevZbz1F9+vkud+W40IhRzzt
JSAQAadV1rJVCgvdycihuK0tPeaaBVSwCblL5mjK4tr+qcMJ59nWUlDk40dNZmSpG6XdmiRkB56P
ZOKM4hWi2DfrmSKBK54gslPZBIn2OvBO+FKNp6BIMClhkl5BJhM96RZChS5PIgvqSZgO3sLaAlGe
ZQXZfZcirdA8LQtUvtJ2DOufKNkXL/VEeY6TMnnMPUeRypl4CoOSTJFAQgFrYVb30qsR7OxN8ird
GAPfYDRVB+Nb4VkRGkyOV04+KkJBOfUUJkEmmQsUif8Hsomh6M0IT5O/aK6rlCiRUGyXQP0IFmTY
NcnHIbWQs5kzz47tpQuJ8ULPBORsyvKqIOVgU7JrOlHMCiFsKjUVMZgyWbnuGtz5XI0FswRF33Rx
hfvtexoxK9bhbO1nvZown09t99MMFW65sy5PE8Z7j7RAUE0Wx0QnedkETjwHjXY4KYROUcAAZvJ6
Qsgmed5WJhoZk4AmoC36YghtNfCe5TV0ps6DeYtgyRAKbaVJ/ugOCiCbXux9AMZnpTrB4iw1bWy/
SIkRPvLbiL76NXv5bfC2XdqaHNfrIY4IHDkZuQW/6Uykl+j8pGyX5t7A1+UNF6O/RoKkX3sPPpU8
RWJ5sn8Tv6gaIKygrPbQvxUts7stUutojdVnlXfjsZ7jHz9jJNSX9kDyjRRt1B0D55sInUgjvQ/X
9ZAIDJ3NtB2IbAtugH9lV9lEU1GHlfJMel83p5LFSDdzOJJ8w+hKp7ZlskJ4I9xCFHsGqbC9P8nB
D/uvCO88M7Db/LvS3XpypYeq6YPrfiAvyQt5Pxbu96svqgphJrnTF0APegSxD+fu7UXCz1LqFmFO
yBbvOBZrHpvgngaLHARNk6GwMoay4V5LUKH/IF0MEtAHiY1tziGJfVGSqETrsiCVTDFlRv7qGG4C
0xR80ZtAvXS2oaoGXpWq7V2Nb3vELh3bsOUxT8amekoh+ZuEFSnaYjoSE3K0etTqM1OIKLhl0QWD
XBp1nDT0uF9/j/UDsIe5ZU6lYdUilnmZ7cKBnrL83gdo6xqFu6oF1TQ2Kpgm4GsYdvJ6XSYqXoME
6A4mSDaw78C9oCTOBrO6zNCvuGbCmJBAFYjtvafNFG5h0IuyWyVqhlLRvPmQ2iBKTl4Grk38mpMF
9zE1AAcIBeeiGZn2dY6xwXiJWIMCeMRxPUKR/TsCMGcJ0Xe64TI6X/zhobSFq1j0fOHaJVv0iW18
+7qAJNEgfUvsDfevjMBldPxw90HKd4DUy3Hvax10MVnOMFkpLCBDJmqksiJp6Z/OysnQ8kweJjAU
4xUE7+NQId9XKULB5Les6ZSVd1xMjEsZAnxGUamJ/q/gTuzkgR+OwO+T8Ozf6193+dAG2TVCG4dx
lR5En+SUumqR4215amAfZEJuQrqlcFisejWtA3K7/Q7Vdn8BBiuUjOKGi3RN2KAwlQnARP5LFXUa
cLJG0Ey6tKrCBZdD7aGy3FD+Iq4cWXGjGIGDVgs6PEYfu8VBGTAARmFZa1KPHbKHvXx9kcFORuqX
uAWrVEyWzkeEgCgDVnSJMyIG+2mi+XLL5TjRSpA01KSUgcLGo1JO+F9Tes58aW7gvils8VPo+Aei
gHKAxzwFyuSO9JzHjYqSHohNkRDyld2tE8bS8q257InBycWMz25RkADy03Qjtgm6VzfwNy8BZy4N
Lltr4vGuXTs3RtMGH5g8uG20cqu7UFhh/qZTzschP6Yx5UOQyfhJAEMtvwFCxTl6iR20yqEnGYuG
V4/lZ3Qmg6J//MKhF7vJprQreVCJi2EasKn5dlOLjX8E5nrGm3MdPItbQTmTwlcabQfWVS7xWHNa
pi1CVrvMR3KzEAzhTmZQ8mR71Yfk3ih6c5qxG4m4LJrrNh6RoLU6g7CTeO/lNmLuAQ/hrBaaLDzj
+JgIFGV8bWpWb74Lg2okOuA2hb0OKM3JeCJo52KVSyAj2AkB+0ZBnUcz09VuOlwciGDdBLTWT0OS
VH1VRFY5dVELF9G82I3/w4ovSHxq2lKSeg4kSJYBdiL/bdrhMG0wqf7FS0t2tPizY/XcNsc4RnNI
GMGcnh//DcW+NrwK4mwQiyq9qM05hGK2hWdEAGXcc5Ic7K4brFZg6XPyjezTzYW8ffStjn3Pz6kh
SdgI9N6cK1ePf1SUEPJSMGYq9EWqH0KyH/MIEvt5deud/4dad3nxd/T7tRzcD4P2TVFOYV7xpEsd
/2MVdORCXZk+JRDX6InT4FqHy2unTx4amE5Yccv6vdA1KuIWBHsih6iTGBZzfOz1gnz7UoAyZREz
ixHsKnFVybktOlDZ4nOEEYTeeNB8ebQ1g/LjdNjVbpeD64Wm7jplafd+OmRLx8anZhyyTeU3561S
y4el+Ufnv4L1mLAWf9Q3UaEflnie7zlmXTdROALYBQMoWPf0ZFhzMok7vMK8YaQznfZ1W022Ocza
0NQzwfBpwthIP/SGOrwTSxGFmmbroThhaKDfliFfWo+jCOt4bWZ36qP50EimVTj+O8HoZFv6mpdf
m93kfoKPnMB3Ea6dCr/i0RgVldntFR+d6HlhJ+gkg0D+q4qxBFCfcZZydIlVp3DGZAlgXM7khdBw
arGvk8R6w6Dr4DByrF7Ss4z7BoatKZcZakCYIpAIIdWOCA2+TJG+Xmwk1z57SArjJLkPcdF+A91b
wY/Qzqi/tsK67pDB92SlPrlBntP5BrS200umk2ooJcrFIdso/Y1oT9dXG9yYEXEVYbtQT8o+f8NO
2XJ+9yVqn4BPvxj1ih99D30uQ5wTs3dgyPjkg/BQP/K4DlL29TZz/Xy6n81hBCiI+J78zPMX17zO
GF9UWQ+117bLVEX9SYhDVqLvEuqnm0rNO3dvL99pC0oMo2u2uR5scjxzDbidfEWHQpXlRvMHiwXM
zicAdkeqOsJ336DLwyPG9mauuZ9TcHbGzBgr7oI3titUl2P280yYt4NXeiLVszUbFOGuhTqcxSSL
2/7pW3cF6CdcO35vXL225IIIiu+AqsZ/cWW3+k/CmmEvJ6Fn8D3DStFUM793QXjt3JnLy9jLNN21
waLCC96dbI9BOEKF7parnJpNl9EBt6KLPvkaAwtq9EGszhd7aYmiQ+DwX9+tqqFjhHHkna55TTg9
QTMP606Y2pPRPwtAyX3snUeva9NQD8YMShSPtdy8uuDQIeTHkmUoOTv4/0GKkNvNqNaeMtolhO90
wvJZQHudJ983HPcXFmwa2I0CYbBP53olg4kXf7R4tIAytaPveMPgjH0lHaE1+4b7RIB7A3BeANfH
2Mn2B4FL0J02vud3vKHptUxChd6son4vQOYqIAdvFIfitlr6zq1TJETs7TT1DAqvoUBKmB4gji/l
TVsTB8vk23+aN/TxX/gpv962AIxifT0Xbz9O9DM6pCehxadcc2PL/BqiIL7IzaVz7suGWkrSIjej
H+z3iSPH29oe51RmLk8u+vVCXpm6vlJQ+5IM2bKvx13Xz+5iGJh5cbG2HA1DcvUcWCJgf8+OOYly
P+Ikvpdm0R1ldhSpE9dmWkce1WcXhwl+SHff6lZNhgyGVibEr/BlIfr20xSgixYIiyr9TfvdZ/7J
pPdB+GjeQFbKCFFKnu8ugHvqQzAu4QIvrc6e0W40AjXbscQYGq9QYwjy5dAnQb35v4+hOrARx+hS
T6FD3QY2Ca+e4euN1euMfb6Sv+LoQiLtfsIM+tw7o4MwN0CTcengkWt3KLpYSZxbNjtEaeJeFkEf
bhYvs+fBC+8486jig8+e7C16PIj8o0w8taC0qKNeIEMUYbRahoUSG6vxGirHz3IYSmG7V0yV/2cI
YEN+E8RFv6PaWgPA7/ybERYyQgndmZiexjMA9xUkVoNv4/mXsct1LPmIvns02elZ+fL4fTpALnDr
JEBDGhvQIfv/Ii+NwzfDkJ6oWnM5W48AJZ78ru1+4BZrhuLMn57o9O5+hjz8mCgCkNCG2UIkiiUj
WzQKf7rKVkhf2g056cekUs43Os8QxhCshtfNcZXGx5lJXN/2HfkHe+ggQp6IdfF06j6XRoV7R96I
Ewi6zbocQQgpFAeFh48iOa4J+xdhEkNdTT+trH44sz3cDFGCKbppFgTvhcWt68VassjDYG/lNf6A
+6AQL+U/v7YqwVnObrPWHP9ZR6wPSE8YuRfmIf+88dp1c2vwab9CN0uCQt0kC0FpRHQORH4Heu0P
Gv2VMrwG51IzkCjAU3ESZT6KenJgfuEDvA3rixHcjFzmo0OniphBVJZAjPicR7cZ795QX40uu0Ct
K++mJqqQKaDWbOtQgWmKSBo1XvlqAzo72NM3Rz7zYIxH9l9irfyqqAjcVqEE0G30UF4JQF2miacO
daRj5VauDw5tc+sIsFZLgyIVxRc/0kvrLZG+OQazLW65uInnLPFF3EJoMeyCRpvBChfzKzO3EJ+e
i13RDSoPTK9EQj2tjE82Eqmy2krhRDmRgBLCRXnr7HKCAjpu0flqr2SaneN4/0aGc9i1H8JWkwLq
RaeLOXriG2uO/3vR76WXRLkc6TwgGItij+rHF/RVc9kDvY3mElfKy0g8b4c86cWzdMSWqnWBjMNG
KJ/GzKQj+zdCPJ6f5Y721GLYo2YuWH32hDCOPn1lJz34ie24FyfPPF75FIHnHCzcn6PHHibNKemE
q0RR/v1t6KC5x6fk3DB8RNyf0w09XgKc7CvYMylJ3xRBDryi9Q0Vx51F2rP2xFPONxM2iIugMWm1
PWUjhGNioD/WrkDBLSoYxNGOILX6vNeFcSmXEFN1wCRR7z0UiXwoVifFYMSX2ZOQaP+nICzavb/D
xad/udRR7Gq/vA/FgklNmVtGA48HGuET/O+azZLDzXukeEPFV1Vwqrjw4HeyBqTwKcQIkVAkalzG
JmWiGk+yHNpS/dniLvNd5vzE48+nsUY1yMGFwzX/kryBUa5IdYv79vXhtdRg2qRKSSlSaM8wptR4
Bu0DAzFAQn5OlYBNLK20KL94h/E1hb0LaFkJawWXoqxWcvPqy84pcmbMEbZQq6//bMMSaIlK5ca4
knJaDWRA/AdbPr15BoM1Gkj6/CfUA3dFcUzgLRCFlQHx94DPmqcUdJomKxGQdEG2s49i68ujzbh5
hwe+vHSuUodSxhAEKqrsHIYDDDmf70vDIrtm6l4LetAMbOljznriVTO043VwuQ7oOcGeZtybsSvD
6Q8NRzF7YDspCAVaCFxakot9vH2kFBnP4JDG8fxLcLNAfwX+pBReN/6Q40HHGCx6EOslRErCAIVI
sO3zSK7kB+Rsn6PiGCGDqZc/YzD8kJ1+5VbW7eYD8B/2O29hjG+fkZgAgYgU1vMpX+TBKVT/wojd
gP9DnZKlTCcZiDxY2PiIsus6futfl9DgYbxCvyVDEr/gsCkubGwlK7kM/Y25pZg00i/DriStLADY
6PhEMaUjlVmIacmzi/i6Hu6TzTOP0hTIa8HTxzjYWjfvZTLQS87lfsum3UL39oyYHfeALW7SNx7c
FpISvq3Dr1APsW9Nn4tSVourLY0Raykw12oJlbHi0T+HYOjIGmhByytRUU/7/lgjvByYKVtSefpg
zrYt2P8OpFffgguLaV24IafUKbpsalFkK8tUKc/8gPOUSvdgLpo/Qn2tDoBx5kKfjTx13j1e/H52
cvEByb/4g8es40sO7sCKRCf9YYQ85L5L2fZ5V993QssZVT5saRBgR4M77FvsmjmCJCBtbNfTtlaJ
iFNGK7maJFB2IbvNPBKvZTKpYbiyMsG8wlBEsokFWRrEjDTOMw5SKSzbjPDgX6r0wPPUML2fsr+s
xN4eL0CzDXokiumFMT9kc2WPajP8Iyt6TLsUfT1XVMCznhdLx1ictDn+qyqtjRtmW/Q0zq/Nzv6y
lA4RVGvH7LvfTAgf8O7KkaEGpeCOYuFZ2WXCbksUrts9i1VQmvYtV2pxiAhbUn/K4ycbAK1iFfTp
mo+UwBJ8MPpnDkj+GdSveaWaykOThMNLBl0jjRf7jp5VPvahoDLws0z+Ppm+HabgG7Yio0EbdvAd
nMm67Pkr1KoaPc/8WZ+U9CYuKuVNrMixfZ0Dc4YsUbgBOeEb8tuTnRcV3OnpKU0qQaSZ5MY5M4fR
i8WnxJpU2w0lYrZC460vWhQvlriidjsyJ4QS6RDmPZyAxhNRsVZAh+yYMZt++Q3wdvdVaWUrRVxa
JKaCS39pdhT3uOL2CIA9V61n0+j89i4onIq3S9GC8NKjQAbJ8YPOUPscmoRlvftYQ6karfWH7bxW
8Q2E9rH/jZJoic9F/RBbwncsqyrojiqmHpo2Tc8Qf6V6uJrwevo/1a+7vFXL7qYMeZ9e8VknG55+
+NNyDMMp2Z9lVBsiB5u/0pqz4sxIxkQqYwoXSSxx928Rg0AivDBtWCnrQ7xDIAEM73uyF8ZFvBco
791iVkUJQ7iXkMH6CtHLFrztcoMf+vUManpIAkNKlzx/Iq94aa4Gem73famgX18LpFomUYLik/pq
7RrdZbcLWBtufEZssnqrWN+Uglpc23ZQSrhrsGq7wqw52B0YkYyKomH22wEOifKZk7avfK9iObVV
5ZZJhz1hTFsOXsOiZXjn0MS2PhKAaj+ys/fR3CIZ6tc99Rs/0OmnHTvTvgnrv8PtwwGTyRE+KhaK
tB8OicAn6l+zvKQQz5zVticB1V4ZQPkNvh9Oe0FXbmcEPrLUGdeiai9V6+a+swGe0zBw+BMaaA+O
SnlTCuF6HK94U/lwqwpWm1sF1+KAcEQRlp3dBcqhc5sLbyTl1sH2iyTOAu1EX59dkA5uWNtWwBgY
zDgXckmEKVkcDBNYrRWvEW4DgmDwOATN0pw4pfRSvzWdvbwrkeVkjPZxtf+VDufRK4Hxn3rR4Cr9
azpYC7SS78pajJh8yhjMeVeE8XFHTsj2tAo36iaz7YLOVfsuk4WOOWJX/N4JTc/xqp+RUOzJHzAG
lxruX5H6GzvFdRaWCRgi48zEZQT107NmelBlKa/y++NPZrPkew3ryJDjSQkmCLurwhpkDGgFvav1
+7Ozwx2lRrlWkdTb4l8cVbLNQbUrDxtGOpO2sn2SIfUE9IZFxA0ZQYQyQtM6sr5tm4TmCsJunWeE
iTknzWzu0AtwTZLq/n2MYoW81/y5dw/bIIoK7Wgs8C+BZ8FVtsNgkTB1l7ftkN4tAv7JwCHJ8Mx5
SArwVUzDFne1rpoo5URE3yPLx8Yj1pHEvLVfkTuQKq01+8cGGA3cUuc8o9H0o1xAHBYXHR8OdODN
oRRWXRlhtzHrSIY1zv1QhflL8CoYeQhmxLZnLitsqqwClAcrXKltkf2g8oLqeTk6tajmBK1OiI33
LAihyET1sOpdAbnogkg4oiEFOZQ2CzlETolXxckL4Ov8flfrSxTws8RZ0LbW3HnEPn0rxB3iu1Ba
3Wf2nNCV628h/rUdfQGeH0S3FUahuhRTSSXASlJXrBfnpoxGdGSyIj7rWzyzBog4uSf/q9DeKXvc
3jV43ncXSUDr/tfarLWpty5fZffa31wKdnWI7nFonuKVlERWccZRHIQ31xmwv7sslEuN6bWy7j0N
KpS0qDw16PyxCzAyxYdhzN906Oel9ZKe0ko4SjuajjSmt+zVB6gcrosiAnn+R1Rwd3eEtSWOB7Yg
ANMdRA5bIhF9DtuZPezXSCC7NE9SxiJ4oN+34IY/ukZqjwXuzoMJxGzdzIXk26yGdfAcGYUv5ZRL
hfTMFmvEMPK68705IWBtvkMEzMETVZGYysw5z0RK+oHjUJcbyvF6hM53x+fML0L9Dyxsj8CK55I/
l7q7VCZYG+9D4FpFQCiVISzAwl1U+JgRLOjwP2KWIZbUHOnSjKO/iDZRnmi8xXE7Kn534c6VpXk9
rXpJQstF+HH/dsAl8YbgQCMzjB1YfjE3HT/piNVRg22VJVRl9li4VyOHVAROq6ZymOOlwaFFO3BH
Jt5xq66IMzwalbdeybu6eWdnqOQajLNm4PfJ+fHE9j14VJaBDQCI4FwUrkF+xQTmnaYrAlDZt7I7
CiuAL8J1VPfmgn4V34YsyzTOlMkiCKJhR8l/hNcUU/Kcl6O7tcf2sGbB7eoFJxGLMU/ppyeC93uC
5lyLGPvhbQWBg+14HX3c2jZhavr9/ZkzQilyQ51j1SsI/v5AFurjxxQocTGBcuOy+H/6lkmPqOux
uhi20ctOYYWlY8Z49BxhsA7uJxIN++CWzZq2NIIWNJVaqywfOYOtaXsc8tS3cf4HoazLJNwGpQG6
EMot0tf6WAuritehSVMhDdghtol/6/RztrME7KsHFG6qVY3uMHkIMXAq4Xf0caQgoaTc1HtakduY
nqIgBUyOLvqf8q1PKl9778UahDeL2scPe14Vrwzo1PhMQNekbEa5T1qGBiYFHB+yIHlniSRiWyiq
e1T2Ot3i7N4zHPvA7t6bfnbFPo3p48XJKR2pfViwY+MwpUF3rqywQDQ6zUQQQoHhgJH+LHUyvHhx
fDnW4HI7GcdgbzMeLQFa0cCz+fL7R/l0MPZFdCrvYkz0+04UkJfkFR/8CwugnWZMxoX9zUv9HQ6o
7g6C3x+O4Pc5voK/w7SmeGBAqva0AcIpaIRDO/SzpmJ2Xnchpyd4VhMAZHr4K0O0Kd6VuUclZnu/
gAi+oIRyuQlkZrl7wtooqpliDp5l8KZc0JlQo/L1eTT5b+8Nd+aOCXuAgJ3FzrX7dVt/qJVOBRq7
9S6gybjv/vx84MIJqCJqhoLZFpISoG4qEjejJRchMX1Xs0LQjvbnBzmBNBBUoYuhVfJEsBTSx1It
krOOXgdt5GkyoccBtxYifc+PgDajg0KxBklZGLQUH+BFwrWV36UosAQRzaILbdls5mG7cOkRQYbu
try3GBU1FGEXZf1YNrUFEsxCWo/0M1WYqVAy0qhSp2j9kmy5MUIT/6XJTowkWpE1L3WWhW6PQjS5
fQncQFM9my9bdw4VxbdUthfV4dvJLw0/apfkqN9Lk4yS52k2WEzXkh94iVMa2c5rEmoxVaHrHyKl
7QVc+/20ZJvyB+TnkPgiumYZ6OKJXL4TGs/EX+MTSG3d2y/AKsRVE9dKmK2vM6ADwE6Wuw+eP3OQ
XM/4jYuwwoqvRVsOGCfNOqrpEcyU5ikML/bKukX6qU7ghlUzxjXjkl0lH/0aNAnxS2b0DS9FWPkI
cRAj28PRYQCPwVWcUgHu12pCmDmsxtnX1GxHCuIAGkTjJ/3Mlu/OiDDK0hnEOoHhF7qnmaaGKIvK
gl8ubwLzBsS2UhXpiutqYSXJSycEO9ClKnwgBhjSuKz3rrINfTUpo4Ty+LYBCNZ/zV6TIAGrthE5
z4H+kPH0GZIzgB8BVCmzkfkp2pik53y1/gHczFr9Zn2vJ40LhkPTU1zx2yyz1zRnpoYDqvLYlAtq
I1Ya5vn+OUwT5ArmRoKo3tJ+82iTSOz6wYPDdP/OcQ6csgyZAXWaOPg6DZcPy+STsYO25c9wWnIa
6nlquEj2tz71F3iz+TwgCQgvqTIHTkvYF+FNgiBy8/l2Cw/AzaLKcYAiMfXfsuCIUgQIjuZ9gJYY
+nMdUZ8myxXrdh5St+7YoluTMHScZEpd61HXwhDcOjTyENQb9HwpR/tZuGZ3Llcg0AnDUO0a9QTx
s848gc5R8oPRCXoKvMG6DulbyGyeIvEEkWAs+JjHTOWw5I/iv+hG11Z7yydOBreXQxqvJDlKj1Im
Kob6kW+4or7DKYA6cJ1AVFWgBvYD/djcUDLKozRZem/qLTHp7p1dfK7cPen/UIftaBGwqTlk0mmq
AACNLD5TvCdDJapPQxedCFZwSqhLO061Xie8Q0hUv4FXVQzt84q7weBuKwo6RoAv0Bw0QVaKg+Dq
k/1ZUbDLzccJvlaOU0/h83IXf2dyVE4ToGZn0PCcASktigND7EQrTNvq2dZS6l7B+rBMrq8EWWZc
US0wDnlI7CYOuWE8JdwDTGp53pE0kl5HPZJAsSoYM7F/C6KcrLYaWhORfLW1rqPA2oO7JzXRsKl2
j4epctQxXid/rTNGxqYhTJvXUdUveu4+kFFV+F4Ktd9IAdI+m6YZib1h0s/d1E3gahUhcs5fz8iL
FfA80ydG0mFv5cjtqSw/8FEUEjo1WlibKBREsk2l7wZUy6h6uWCLx1TF9V4g8imTUuZqlL+6Rr5B
aBR0uarMsiD7zC6hHRcQSI9epFT2YpV+UxRU+DB+40vIvYYPno+aNPMQYRC0y4DEd/EoC1W4QHHx
zsQq0PfmIuPCfsxvouji6kDacL6XV5by/zi3LirvfXs4u7Itv4/pRQULNNgAt41wN2nMclc4OVT6
vVa04oC/KrYSgFXDunduAkKyAVYg46a7VHGo2slKxg/1xB+wmXcpKBnlizBoe6E8R/p70WYtUbjB
O6iiCXzl6BbwN7drf2uhlHHMOSznRhlfiQ3LRzlqj2g3sVujhTvrhyD4/6GxK9rTpWTojaNTYdC3
PKukgDbnWQ98Q9a4FCfuIy853KHkQcAlyynDl/cv4xaQ9TLBmUwUJHtLGTAu6vHNRQbVYOa1NUED
N4179LFyI1uiUoONaG2VxYtIfjTfjLrHpzjQGbD3FpBiuaBjKTpYrgOjQO/fXJA0CKhsA+usFPiM
fiGGRNqsVW8GxBlkJul4ingMU5Wc7qoGqXIbo16gjkoloWthO4cq4GQOTZ0S3rKKrGpJM5c4u/A5
8vZtE712GX+pHAvM5XgZCAD3M08Z5tP4SGKuCQ2GfUxCmge70lfU9m9Jzjik+gSthlumYYDO9QYq
pQvsl6WcUtHx6rl7/Asuykieh+3mWDNLnjxK6rwMxIFu43bbal+O8LQKWWHlHJFV1C0fEB9gPpR4
zuvbjgEX5EsGLgS00sh1zdvuthY1u8Y9iyrfCGHbWMqEMiRGZPSg69c9hJ4NQclMqtHi/CNFA+VS
7bUUqKiFNoDdTNpkd4EhQzDKNeej2vNXw/uW+5u4c6qu3L09ipoVs09w/x+JXDn/BVk5URxoXdM/
/OeY1NrXqYKVSZfu2vW89zUjw89UpHVoeo3kfkpOJS+X4CvwxaEvPJrWfGkcQrT2rxfUlHFDq0EZ
brCecBPuiOvl2mPCeIpJ7S4NOCmF5qMvyZYTeagpz9Td2I0CvDYZJvXQxMo3HzAHJNvD93QKqfBs
inh1PfIIFUFR/hsTk6zGn+osM0/yXUIQ5zph3imEmZ61aKoxbBTAgipWe76GrK72Xz721NoyP5sk
zRj7cykum+IzOQFF8oIuH7taRL5nOLgokls3UVktHfakQDBn9j9JgdjLCPP+6wmSoGz7780fXmBm
ayNwyCGEvKPe6+n1NW2pIQmFECyAUJtgyxyLjy/WHKCqUjEVaIKgPylNqY3br5dAYa0gf0vWWjff
Tf7aEuuSYcFHj+5sNFRGRpJP9rySMb9DJLkMC+cSuCWALpmdZVbo7Dvhv18HXSZJti2tO01wpJM5
2HZekpf6yBWo1ISaQruXVuI9yl6tEL6VFaqjBo80vE+cDTEpxepPY5d4esrV5aG9bLzEgNxaAhN4
1rJA+QtVi2lPGRqi9A0L1R7iV3R1pLC9u7lMFZGMFzj8oYgjOrc5F657BMZEE2wkq9dKsvs5FVJX
ti1utzWb5NUkiRU9Jd8+7CL9BQwDUKPaxswngcZroSHkQT5gV8DUWmYjrdc8GOp/xm/YRPsjHcTi
eBaCxZoNmLs9DcHukdL2LAR12kyPDwAL4FcrL5xwlekEwf86TmOMvHF1gPKndqe6TDGUjYKdr78N
tNWv+E/l6iNs/m5TD2wgagvzcFAbjGsH/0bsOnqn1VtbYe9SD6BeJR4m8h6qkqVnjDqdFpSRvfXO
I97XFMJvwQnehuuHJnrUM7NfO/54+yjvZaagOHRx3Z1QfsNNBQYsfA2US3r2QaAT8AFhz/FKpu6L
zxITh4rgDIRSsnaxB0cY7mC5jJ+Bk05zIOUm2g/yC0AKXhcDjfSWWiAlypXWxCMpZLJKRnLGZQ6x
qxETRKeDHOZaUOpovOY9mIDN8MWrf9tSsM/wiCEnxykFQ5lD0Urn/YSCbXtwtQKoaZZk98YkO1z0
ungUUSrCVLEsWN3eLqYgSJ72oXXXewmSPgwKwT0CgAWzv68BNqsby2u62FTpPIsXTzsgqUOZ2WY2
IgHfdEDfKlXCOhUBwcjBIP5NeOt/2SRZQWTEsuxozEwGHdu9GB/pBCtxnZnwwhFvf4LWbR/q2GxL
GBzsUzYGqpCxK62srpej/rXGeYqKNSUpEtyRiEl1gM976jphC4a3sLcTRMBYHqyIwn2ahxHXP1Vd
abRdbM7rCWwmGCGqMWxgI5eNASZ5KMZJJvqQLkRA6AeWFe93QQRUyY61oWie+OnR9ky5XQSTGhF/
UG4Ycde/2RqxUlbYuRDm5FAhCaIIO38ACAi1vJerT9AZ3vMeBa42ETq9uecWsjw2DMV7WoAsrq/R
80JsRqHPlv1xl2a5fbjCb/YCXgqJBSy1WL5nzSP+edcpeNLVMoQbmObQqceaaTX9aqtGqS6rZT1G
6iLb32XV2Sq+YhTQuF+pA+WGtIJN2iWZKJqU3eJbwXu7ri+vJIdulzvFEU6q9uoi85cDCPv5UpzO
orWdqCXlYRIHl5BH8vxkX6yPMvz8aLAPcrAKRaJ++eOQWbKvd1xCtHe6reLeNdV896CrLEo31p4w
/XvzytWtoUuojYdsjBtkZOoyo0psQz03D4xCuugz7Zrdi/LNLZ9VDRBd8vT7jUaB1TwORBXn6o/C
gBn/HN+3c9e1L2n9Skum6Iof1aTIizciAoQ2cystoIK7VMXcUkZDtYMfMTX0fIJmpiqL+ibG5uba
AHr1zJttBK1rDlK+mZs2oZPug/AgGc/GRO/FNBdhSVtRiviS+IVJZijY4WBWBtYj61vqtJfOsGGo
b8moYYS5XSAKolakogMBNTgYGyX8aQdQPqG8GodPwRs/rAHTjuRfPwQlxW3nZYvDVmq2hXWf5yG/
+FJNG5eFt6Bhair/UqsmoGkCwf0tM2cfwMpnNp0YAYxt/ev3jKD06hdRBYxJ7dV1jCEQYEEgFjry
qIUxH+gK95H/J/2JldwVmXkMOCAEp6Hh8JI/YglrLbCVkMNphalDvhFB1L3YxVQ2akcJzZQ7TJkN
2z9fnwixNn5BY6CZrFr1vrZEGzTM78lrfVeYFrXs+TW9LYuqCifk68pbZ086R992LDwktoMCSWjs
BcZLonp1ux9yIrlO9uIyDvPqKKOT7NZIpfNVwLFLfRvUGhSnilzZ8GjtP7f+XxazE63SXdWCPIb4
J6gPRSmdGBMgJQxEbHmdiNutv0P85jZBj7AUulCSv4kSeJNfejHxnVIpwKTg533GIix5zGIJyjIR
rfpvLPOLzNwLhC4O8cWhLxN3ftrQPPfwoBRCYtNN6vFmbW2vUV+wwjXRn/8I7Ocl3Elj/EUtACgj
/98wva0cGSJ36nS9sBRMdyiRcDfrbB7pCHFKmzzuT64pZxd//0qAMG+eBHgYPoZ2k8Xb+KxAjYR1
ZkQKa9ZSiNBBeyryf5VygxJ8Ah8rRx+JkodOLKTrfsnzu28S35GizUVEMknboTGa+lG2woR5amiC
3rgUY2Z5Qb5z1QpVoVG4qLyfmBmrzA927Aw7peGLsDw+ODPDYk2nVV8uqp/RFkZdAU2nrGIl/8TM
hi2MLw5lynC9xn3sZbDfZxfCtvjnY2OaRohPtA2OyJDZS3jlhYxRvGqikKGKNuoZMTU96FKKaJns
3gvq6JCiyt1dc9Qn89h/b2mCVFT7swBhXAshvS9gXx2+9Qcuy8sKJkXmevfrolLgqDtArbRl/igh
MXL0/p8akNkJO4CwC8tHP5UbBJzF7FrcC/BZ7spqPivirKyXdngtWOXCV+DU2o7zRXyDiU6JF7XW
xV29GQ5aBREUjnKt/dbBHb6CYNLSZ0jqx+B31NZJTxyYxOH408pOBAsUejPPg8X9ForDAob1xxo4
Kc8RuyR7YysQa0z70C43eJAqyt86b7idRJMp+9RFUxDPhOtCZT0g9OU3jJ9dfkIo/IEQ9R7gLxu+
xZFNabJ8Y9Xm4aOCe3oHxyCEiTRQdZ6vzMhLWpRCbYm0y7rGTnRyMgKWQXTBdFnvxXMv0EoOHm4n
4MODKJ0FIyi5e0ROX9kjRnSX39Y5RLO6VUwqQWaZyTynUU6+XozwHrJkQyxeSvbQRxjxPPRbpthU
IFKGygKyyahSdrj19tFwCaKNT938OLP5VES25fVYXDRUhVgyA34aHOmibAE4f0Cq+YDzxG6mLChQ
zJloKPRVcc19uQPA5ja9NBKiRDOr9+sndU99s06/yHfEoUuDYnAWcG3lR2LYoADtSa3eDXJJidqj
FbKiOtMjPnk6TDVv2xwycjlljenxqRCJOdBLvvUQBRDKleJvISRxar05BdsBKQRYgVcBXssA+Zl0
byxrkWSxkdb9etoyaTiRvuoQt3ruS5wCTHo/DO5vd92ehgXKbJUswURNTW7V9K+q34SItci3TRtn
rY+aOyhdCw+7XKvEoGAXxU9Lt8R0TlAAKgUIbPguQY8f0w6oKyZ0k8NKwRNsEbryWdbp/xsvj1fW
3F6kKsOdSkQM31GNccG/vGgFlnBNti+16OWNfbSZLo5QzxTcqvCRcBPg0VxQDwynPk1Dybjb18B+
osALbaREWRranz/1NrZvRlpuX6DK8gFcA8fKUgd9sPMutXxBWKb5IgGY02SiWYKPjY6s7jlNPMuD
KLaO5MrgPEnHAagC4qcoKsP10pI4G1GZ++EuYP3YIxIidLIWR9T/j0w2ywWnHOJhHU4W3ikvVE+B
Dt0lRHAbVVqXwG4K0yxxDMeVkjpwrgMTzFwjWNxePovV0yahXQ+RAGavdfsQ6Vm8wdbVx0kIPB22
zGjvjzuxft9xm6L1QJ0IgXTY5zeEihgq2U0XXyEEQ2E7Shtqt/51v1OZ1yCAewPdTciFyWkj00WD
BbJXOCoEu3eiyAIzlBb4/8p97joDV7BD3FBxMpqLGszfiuIvZLkbYGyFhuhLeTTLCLauRv92WuUy
vaUZHJRWiJW/feBRn4i/SKFzACxQ2WnmizwxNdoZuIcf+MNv9VL0P23d/+w0D9kZGAqf7iQ5lOeU
mRlX/Ukt44uFSNqZs4+JGCNIFF7zO6imMbGg5R81tTVrdzJKXy8JXDjEzLZ5qyW/O/OTlamNVv6l
nzXIhVOSheKjO/h8g9KDb0ONSekadl5ACt/UzUhdJlJtScpNdz7e+eXe7RRmRirBx3E5Lynt/8s5
jL3rudVO+omxrYIAjxnaaOyu77zd2w3DPwq2oD2gf4TJof9jw3KMZkLA3UrE2nXURmIBdVDxG+nK
254s0DV9appd9zH1E9KooDvttfbBu+Sy4DpMFuEe2PjAOTcRkkDe+bz9/fkqhQJTPRsswY40QV5M
n17oRS4FJ5HLIOI9Uw6hXf7XowX7QqqIqHDypu7xt9YfLiPcsq+3vatSt+0XOhcHkfekqvbXp0c/
Gx8nvZr4nIs+kx3ATwfazucpktUAQQAaqDLdqt6PUUHgnl6QQ2HxoofGzncnQvEIOIaa7h5UHgo2
HGX9UcntfkHO/CEWNM7sJdDnxpfzXPmmIgoVLn+AJdIqVxF2OSdvqyVp7PTTq1gDlPiuZ+MxDnAJ
xgMREfH5W8BQ4BgmiJKRhakNEZlEWjSohelACnG9LV2Xh0m9tJEgtTHArYk2v8hDIMJMz6cOo9Q6
W4StrUacsgQ8P3DmcVMwiZ1IwIiQJ+pCqSucfx0vScG7baZNqLaexo2/gwtNYTY/C3XsCd0ERJe8
bDucfFXpkdPvjXqAyPJLJINJfz/CuPYRuX6nGO1c9+JSUwoByB2XHZxTiX2g9n10pHWmRYNnkde2
3p4lcA6xYtXOZFleP1mqs+Fayt2ifcXd1mBVxvpVDleQ6asVDlNts8to5ZWPAHtI7A+lUvdEoxE4
a9AYqLKIm/IYiKSrwX9SQGTCxFRoYs1/hZozz/f+II7g+rAP6DPdkQYmb9ArWhO0CqHXdIMLsNfs
RmtMz1xK79Kfnq9S6CS0N6dfO5TENhBiwB9c6dhYWL09sDFFOsP6nt1KDmh7TFlM7LqvqQTFZ18g
2g81rbgQCCW9X1dNfj5FFb009bLNwvRZaxCuZdJEd4hMWQ/OQGR4oiPvnw+xjibkt2OjzFXVfiPE
XGuUQC/NqiUUpYW+2MKmg/WuedPZB1fnPWZFydjYOJ+IVrfBHbr/khfYXErv+LtMU/iPFBbBUlb+
Xq6LimOCsIM3uMyKxFkvn6zVz2TTlFICNIflr4d1OG29da7wTjsza9H6NkkqJzpsrZhgwGn7hOAg
Myh9fHAZu5ywhc55zxc8Lk1wk52Xh2Wm6nL31PeatBjrK4qgP2A0e0uLwDSDqRLdMYGGdkuKN/I/
OxDBdUHhVV9M9rTR9YjUcoJva+9PZzCRiuBqwBuVWXqB2ysXf2xeZlDCFx6IJ58ewqquF88XN1eZ
Sz/0jwQ3lKVW22cXCLfUhyI3mtea3Gi9prtqFpdfPYbGlNlMe9OiSS1XDO2nNL1NkMb7APGpNfuW
5mTB51StzCflXFwuP9tcW+ljOTubmd9QtRWdfIypik0kQjbvuM+OTEt1x+yBxn3ivCan0vgPBBPq
UhaZvEQtQQU3Gj8BLcu1aiBzHkpXJ3Dm+H++gvmoodEyN3E/RUAfguXWM+M8k58/E9ZfEasCjrfC
AzzrJmNlbun6ZQ8knTGsyGolGVH0AEJcWZUGjCH4KMWH3kPnJGRt1z+fNDk/B6m1UfEBb3GFJA+J
Zpu7S5OfYUw5IdHJ0wVOYySmh80HAOJHPdYcivhEpuBi/YYk2VhU+ObyR7JKAGOxBXsARvMPlpVm
CvgZjtenX+muL1O4mHwpGse7scyCVcykytaSLzLrjqUlji8raZx0yM9iwFx+T5OYTYfM/Myw8PIK
0IF9Unl1HCer4Y8EQb6j+7nhdvLxRMLe+fkC+N3n4/KptDe1F2OtuKoYohnhPVB9gqgJ+9vSN5E3
GiQmzUeQoEUq3JjJZpEOiYFH66TbIGYeWt4a5GVtRvScAWp63203xNvV3aMg8ko7qtr/xWkcRhey
tX25sjwKvotAujrOvfegQwhWzExBFS7MGCr6pUuKfP9NaAS7QpYOGV7EdqdhD+k2p1paT95Pmqd3
WmU+N9vMo41WxuoPt3+zGVPX9t18HFgRxDfHxXGIgR4cCHMQ9arBaNJqiu+aiaY9sjNR1mVA5g08
F3cfN4iz0KeTC+S/LCJH6Jdhs8wrKoXxXfpiGQzttYQDMWCw9UPKMtwYAQNrj7v1Aiq/FlbaHGws
Jl5lGfYbMP5J90uADj2EJlZKlbXmpXCJqorhgkjGxeDwiiWRszj4wCAdQquRTHHIXRRl7YM6Jk0W
rd70LlaZJKJlQ4Po1kazHOnBaZu35d9c3loVOrmlAGRDekP3M0hizKwe0U3ifY+/5YJ1/6elkaVN
Vy+5Lq1Byu6+zBkGAdO1lqyvws1CsRR6XEq6WQFntkDgddnmQYJ2OlYlDdpCNBf3o0M+pZCqEgnq
hRN0m0Q6rKVM816+aPyqoIiJsBvSqjMliCxUVOfMvt2X1lUnRb0KTu0uo/M24PBKK62Neiz3qQPI
CRBhk8AtSAZ/2oqqnbPte+rc0fx0Oyh3C10FoIretFzf3s11NscWk7aZN6X2L/6Ydvddl5+QhD33
xa+zL2mMIRYtUnrH3VRNJWE6iSuHY2RXLLkGVOcmG61pWfoAA1vhb6F24jH/5m9PQQ9ieGUgjJK+
TtVuiTx6Gzyos16OYsBEPu4WRW4rhzgvS/telb3ZjPrqJP21x69KQ6RgHsHI99JdON8eVh3T9c7u
5VCqdx+F4Fw0MR322owu4p97n0uXRFdOVKzAkOLhe+8kqwVWLFRhjOr22C8XAM1WFSHbkoTOBp4z
U+8VSlj3ohtG1NEHcRB9Ev4wlnxT6SqKYxpECdnvuftp6MmC0IuHLL3wFUN5GBbmZw/Fqk1ntKEK
YkiRhbgiKGUC+5MBNZqb1flRmwQN3NZs5gVsD3cUtRg49iwbC46SiG76nE6vgT1jbzCEo6dcPitF
+ejD9ulnAcC+f0nTNLTxuSEI5ToLgeRMVEibAkJxRfj8OPSg0MIVpT2gA6mXgEDOdbxwYBfatLrQ
j2kCATjqUdQ+mTJVhI2e6NbpV2Bft0km7+qkInnPGCHr1/TPfeDMeugpKqtKBRfsgAp1U1oi5Tc5
4ghBxb8LLGTE574RIU3Bvd0ONtbj1VwqiydqXS/jgENm+D8jDyu/pAbHv52GXJdRRs4Wfi02xqwq
+B54yk1OOFurt5Uq7PSVXbo3Jg7EspkFkfM4WTJoKT3yvuWBymW7rcQD3PPYB4SwKDa6IIuUx+wY
MPK0jLtw4xFcbsUlBO1O70cCGmCdLLp2N5cwKlAAvyftQKOkSAu1x7g27pyieLZpo+6BrdlGtbBh
yr3TI6pSWXS/CtGQx+R5BD9l2I6keA16KnJMC0EgBnHdoAdW6Vi0a/4b2FLfroyF/Wu6sK3935bV
EB1ZL9M2wdiFQrZ8za6lz1N1WEqyPkJZ296sn11p+8onDRZ7uTv8zpxtwWu5iuqs9SkEz/Kwqn9q
yX5laLJp0c+zPFijO1TWc61PpFKHP3gZk6LrV7HjL2O1RO8ZXVcasvjEwYS7BmNmtJQYhN3SAQlp
QfkG9MCilcBwixd83CPL2bebqYx9nKm6GyUCk8fPwXC6ext8g4FU6EyQ5OHN+sxq2uB43GT7z4oP
L4/GIQk6pUVhKz+GY5RRg5kzWyYbQQG55Sg6p1hnyztRrnOJaTG6ZQwM6vlEqCQMh2ooFv1wIFzX
QvzHlF1VvY34x/wYDQUIPMVTXP6rXL4u7f1PfKXdYPf0fgpz73w9TnGtJZHziEOMI9q3oGndh/Qj
Fu9e9m7pphQ7ODVG9sm9eLUMCbGw+iXCDGmnJtPtqMRbZQ8IIZO4wiLRdTZteTcw8Lsv0PYpQiP8
kHAZvUmtNqtyRHXyJzEsyxs/ZkW7IExIAcyNuA0HbGUM1FJYZUbLI771Kfz7wWrrK/GvpNt6kvvc
CKfTdpz1IwuC5YApHGf06xSUJxJ7AVMB5oQrjs53pPqWeWTwixyomFt6ZC72y79Vq7tz1poTggoa
ANahx4y31eHyOUM4o6aH5xOS/WhE51oyTjKAVN4gqrRJseATstPoqFKtp0O4SX6TgQTdfvGednHH
3MfkhbHdfqmbqG0QDp4WayJOmLVVCIkR47xz4kyrb9n2XqjQxbeiLlErb12FoV2M79/4D/NkRkwt
o4s+HdL58vtyuvIh8Zxzwez7O47S8HoYdre2StszcnQDaoto7g/xQP85BUbvs9uFNsgceHqqWyb2
JNjETKhYnQdTjEvBfQqxuoMnioSgc9RebUyH30Xw9OcV/ZW8KRJeTR6b90b+PGdPbzgJkBMeWdrt
8PtUyRl3ZB4DIiN6Utso5xgmrhRnz8gYCBdTW556L/YRjfRE7SZgPUft9/Yv2FJWSoGJbqMvhhDR
zu8QkhdD15vvM65rqHj72Xau2M5cnxJoiRJ6ufwQBq7Hosj/7gBWgOQJeyWf51AI3/7aJXY5bhKj
GWFdFdB7NH19g/v6/FZlbeUAp4RBEloSyEeyBbXLN2zWdmf2Uu1fvPAfS0BAOcHTBpSVhPRBNZ1/
oqHMLRhbrhBrAL49xDckQt7z1sBNJXTl7zBNsL2amgFTGe/DakWE3hMLtuCHs9GNxTFHPW8uMvCG
v9fFoFbSYtjmK99UmXGR7rk1pX1GYvmwXVENDjrR8u+dh0el040eDUfPKSMiHlp8WyGO0//y8kp1
eeP8n9jCdUQSJDBVba0A6aM2g7B2D4kP+MWamkbYCf+9/Bqph2t8/T3tJgZmh6eyBbHLCh2miU4T
vO62WFLa+xzwIdfYnza64GGSPQvCL9E5m8Z2J1whgganaIfUmoCOYK+qO//qikWX9ernt4Za6j6b
A0Obm8xmvFBmisKj5xvAP1a0bf4Eve9Ik+WpRvM+RewNVPZTiSnZn/GpHnpYZD5MDSiSoylVw+wR
LtsVJIdv3gi4uZLOrmygMOi9o5xDQz9l9HjBco4kK5CbW1Fi1ucVq680vRmQflS4KECH03zNvHQh
/mxfO3c/Vvat01+0+2SEa43RBSfDpwPGzr8Dz2f6539Lj8rVx2b4u+OB3XSB9mKBwKGhket8WmQB
S2uRAF24CjC+nVh+mR6tq1gUJDA2+Swa87e3vflSi2ILEWlTTEu/8MptCQ0If8m9w3N6Q0jqA7fm
uM/HlXspjcYpt8aj5GySP+bIoVcHygOyZYPmSRKd3dcxw63EjoO+NY725sDgp6iMp0aWlLeIE7X6
zCASNx7nHyAqnLQh1KF0+ixC1nDuH3SuwqjMzyjibHUGkjWg13W0s2N/u4nRXZ6lN6962/bgmUxY
J+V0+3uraBg2g4AfRcjBLhK8yU8i1CiyFfQmrs3DHziuN6qWqiMfMXNVIrrbmuwL3QHsoCGp30wC
mO8emzWDAmntK6EpsiQ+HK3y5J2WmHviTgUWW8koGJIZiyzOGPDDQ03HM5UQh0fQrz9iegjypB4Q
HoDfLerJqt+aa6Pzu/e1pDcDVk744UEndDCGHrkSYmArXYUcdD+1bIhf9LYC0cGdCOE4mGQPoFBD
AAeCEMhtJHJgms2CxfHpK0qPSTqPmEEZwzX9EITuNzEl6Nzdv8EJmuKSlzivXg7txmuexWPF6JS1
7/C0rMqeQIJskHl9L7qba1bd7jNBpPARftqdwIgY2nbMfFVmrvLfS1k0/A42cCNPfjdcBRzxRCZA
0AG56xGqrmNOh2kQSLaKJdPaXRu1rsFgayXkWjvMK7iR5KVa4LhXiQPXk/aKjInv/Ds9e8PTrFxd
9zsKTn2vZXS8081aoMoTbt0CQIaGQ0q1QDbrLlIqK99IQLa1tLJfEsHZjXYOCDCtOIMRw6AqCJky
CTAQIActLvrdbx/Ij4JaazaDGqBNwVvCQS84osWobT8YouvJ1c+rVzI1XCUis8mHP2vI7DBojBd/
haY8mN71H02SQ/J4muEhrC05lyM0i1firb4ZD7I6ZS59oimQUK0i9ouDwbxwFOmoj3UD1v1T8jB0
YjSTzxUvOJhBV5HkjYuvZuncmzm6yKgLZFXlG6Xf3Enf0xEbAHHnsGNhbz/bY4KCDu9z3PIAfo7t
olHPEAvEoppVb29IvTVGMTbEf8UGPN8tYAJif9zzsvUfa3MvBSgcYNygsUEQV5RROwnypZff9Y69
WhB1bmwQbf5NvqXvrBLhAkGAcZlyFs6cUhGnXiLnefCUCMetbPJoi+WKUHVpNcMUaMjIn2Qdnm3A
ndDpZPxyN6U0ErZKwb8O4tpQcV10zlgFtpWnkNphOK+c/JgXQ1x7FTHE8RN4RAvtde/fZ8SC/vAl
fmrlsGv3xZNX/ImIpw8aGb1g/x/5qU94IboGWnBzwxcyZGfQyX7cFt1a3ABaQRtAdMlRrohN3FWp
MgDTYYefEtS7YBVzgyTKEpf5s4+RCUNJRYoSGzVrhP3+CaxEaA49TwB4KZobwgdpSpZ+MY4VhrxM
vCvqruh5y0ACvgA+HzMRfXNDbehjCz2JsWwv620l3euJmmFj7e5D5zE/wfI6IgV/Mh4q+lJwUOKV
yueBjs7mIWZN9BCWWend8a2ZhwsmZzh4yHcub9PHGva0SNXfyN8DFvxMdk877Vxz9sDuWhczdKeq
7MfWlwN6jSlBqWpP308sLLiYREYirx9ii2apydMdzCF7HATU8u/PFt/gNGY4AJcLUEN4zDlUAenf
PQUi+yLok6qbUDokJPEpjAw1qGD9CO59q1UJ41wVlh0oHxwkY9kMXGq2z81KfHgpAs1KTZdaRVNv
t1/A5K1TVeiIOwy78yvLSVD49+VonIub7OKTfXHCO1by0yDJ/rFmUKW85QK2EX6YwToUDZHxloS1
pXoIvwC8Hg02seQcocHKT1yJ/0xdQxSx8z7y2a5YY6n3i016p7N5wYpCLrZ2xvjODL23F7nEd2uW
2z4SOVx1vLaAwZQBQ6UCGglvPNyl1AmBLwcw1w1DP6Fktt18h//NiLeYVNfHvZGlJQgF67uhiIRQ
QCsZ6OZfTh7jg2YoakoGYhPXX8JBQxfxwOgzPZmhMCEuoG5VdiZ5DEZwIiMDj140Bo+j60pLkAAk
eeSibaGkp9WfPT4+eTJcxoGr/X+HwL/EU9ZDRHQkgObegfwHFvY3Jtfo4HXpX9oNPWkAx1pM8Vw0
0JSAjtBytnK3c/7wxJw8hb/WloR9CpDTmGHnAQJWqdYhlLu1011uNf7zQYh8o1mkwmq/YPaHxnzS
4HElDorho6nx3ZY9zGXNcU1b94dsLfPR9Ppzv1BMddZpmtZ+E/7kZpoNOeoDiG+9DlR6kRplRv5R
no2G21w5iGnAhL8eu7ezsO8dIiyxgS+PW9nxnqEKyj+aAehuk5ArI7AL7nCyHgAZqzRh+rK8XMJr
ftNPlVk3fJvyEDpV47R69wp3TxEpuuGgXKX5iDxbf9XyjaloCcJqt5LC4trNcuf9mDCQ/BoMwypf
zy1egm4RHWWlQd+GucndfMYcEJ/WlFYYpXj+iBtybFPq9HeWw+77icGBdyUu/FFX/vKxm4DsgY/n
j+SscjrRwC2z69LingZs9ttJxTJ9/wZxNnCIomUY6cd3Ls3W5V4ppKM6xZOl+BfLbdzW+pMYCXXH
qkFMwBCteEIf5NK2wxWT3g4ezZqH70mkZLHMZphvzh/0u+GbMTtzXglBvTxdY2F+K60wtFAqeeFK
b5Ry8Pg6n8jyT0QirgxGX234qhm24n+eB2l5uBzALsrpam0JAVB8em0MxQezIGXRrGrsoz3+s7Ru
pHdR48km72lSmJzuiVflkk7EvKGtXdYp3d32pGNYff6CzFQO7V8EcCRPcGrejNZGxIdL7C5MLDmP
ZB/SlgSe+pyZ8hnEFQRrBRmuflCfogGCNNm6qigIUPTf80uL4tenz+S6Eoe01hbMoBafeuTBuHQ9
rCof3HId8oi/NiD1Ij/KBpd6JI3inrjds7FHg4qx5jP0wMBLmk/Vf/EV0EnIsoYrdGJlquXCae1a
sNqsvBzt+KwnP1VQ4tFsG0bo4f/8uwAOx8ZzyT7qhBayjD/MHQmNsB9TVioyh1iZQxDkNf8eI2+W
yGZJFpKfehlQraJ+mfm8xIjF2QzLLw8vHGEh6dtr5DyOrnNLG6gZxEI2eztnGols4paGBCdM643l
GOQrjLCrZm0jnvyrNAWIh0utK472/c2EIVqbPhje/Fw5Yi/GYNr6JRSV8mJczKwjmGq+f3mta/OJ
kYSao/A127lyro/yXyVJ6xz6pwFy9U/lA8cDVZpwZrlMB2ea75ihaVL72Q5E9ZA8Cw32oRHWvPH2
ZOQsLOXjd73CmIrJpt3thGxNT/wXxzrZ5VnOXGmFAXO/1VEaJy5vrplegsv0tDYc//HxqUkVxTbz
Qec8e3LkEkMlYw954PWnK+cFhW5PSDeBaxdbQreIykq7+Z33Bz1dZk2ICA8KFmL1mTNYGRFEiSov
DroRMKkurRvkseW8OYzVVeCZ1PIlkwelhKfgGLG0M/ylTddCg02JB0xFxyXqrwdUC1QFCklv95Qc
7T4uAqtOH61nPp9q3gziwugKHh7aeSmTkxHfC7ZsG8bVCPaHHf8Ps3hyCRzNy+5IDeDs+ymSVa4S
CSS5Z1y+757+Wesw3jJhhxnghf3ENLH6d/mufRDH0iFOigkIJ2KUQEpdC33Rtr50xRBUySZKnopO
PHXpzh7Za8tj0AgQTkmEupOEdSL6mZ1wDcsjRecUnZ6wCf3/bQEwpVZGThr6P21OrmdDDRQhRVOB
96g3RFtfxjTahVeyGPabN/uaWLPbyjLrQvQpWVbeXfm10xBMA/GxLYw3g7NdohozSf02evCmQI6X
ZT2gcg8oxR5JEBP7JVM/qSQ8kvNCAv8HuUf6ac0umMvXwD42IcRAFaJkYy1piSdgtnvSm7+/P53V
WJY5WtqMzLdgCeTV+GOnZVky13a1zYJ3sc6J+CyF52bU1p0NFd+8OKx/ymWwJ1BwxRhKXI/KH4zb
dd7ODYEFvPyk4DN54o5KwEyW5daOqcwyrr3DhZkV6x3MlLpb/Bg0rzRAXEkzh/GNg35jSG1QXkfT
F2wQTHSOnsHEogr0UiwTg0Fh6vspP0X5qoYmdVJEjWfMraTtHR0PifD1dawBukrcaRHigxOHP6iN
/dFmeNiaWw6pS545wPULwY6qMaE3PRk5MG9c9cojnrH+G9MvUDXdGyKqr0ip+UhWQsqpVpnKa330
PW3YyvuvVamKE8IJWKpyBAWHuR2J+K5ySCuLneYy6BUJ21lji7rwg2r9Jbva+++FhetxuBY1Qefm
fbUiRGb+F+0OGeQQPykTi4RdtE4uVz39Wqs/XKZRMlWf3VQ9r7Wox3F73PnGMm9V17cbR+CclEh7
B/qJ8Darx4MjBC5MV1cn0wAOkkDNzEu09+sIHor74dvs0pgc9Hf7C9VBFzj1ATbCH9mtCCL5Phv0
s47Qxz9BZhUq6kZzhDaLWaWYfsZzlveAMxxPwdz+tu0oJzctFabNwmvHdqhmt9Uoy5BGZ+n0jfXb
hJszZV+DwDNxIBCPUiPzsPvp1Cbm/YpMJTC2rwghvWrfNUSbC+Y/4RdAB0l0umE/CoonSPwtlZOR
06tmUXht0p63V5Dq8jA2RnutCi3FS2+0OtD5aHkPwihG+lbdKyq11RKNTZSp2YKrIzvUHW/NfKZj
e68qFCfZzHLD8yOxNhadwmzKrMQXQKgU6cWUYwFSMpmsU6BbCIF+WhtQp2F+JoCR33sr3JeMepaB
8KnSwGQCPeLd8Oi0Qu0iVyOxK13TUsDwEAJ6xObJntYof8ksyBl+YKVFMc6mj8EIfONZVnbJUBjS
YrEMMM0VhJl/oYU0+l8bUDsRqPy2tay+7LFpcYCOYqZh9aOkeE6cAqBgSynC3YmMzClNaHDZkKow
YOAgCDU2UxME6Ric/2xmHC6qOkOBgiAyoncPKOPLiSRY8RcIk0M0RMBjOOsepzP2b+OyJcDhf8Nr
tVc6IW/pHzov8RTVTD1DG0AO90TbOfsIe/2pP1MvDElIhlnaR8dQ76J0hLx+nAu5HB6wxVA4vtpl
bA6xiXbTwC6Whqql2gihnvm0ZHbF2vM7aYrncp7glHoned1qij4gF2T8loxU/E7uNjck/eg7ZTmp
cwOxOaOvg0HlrpEuKt5tnWS0c99diiZ4p4/oXKPqIB2KY4g0uhUegMo7gd/1WlUSHa7cMZju+tzK
bLos+AXS9QoVmOph2jVryJwyqJ6E4ZA0DwBsqYJsAah59ECWZaeEmPYeLlPL1DGSlN+/WPf9covu
gr+FT3AaTKSLewDnFmJxJLBX8+iEjnizTXEIH3spcrcHi375mpAIaWMVjleXWKkq6I/i87s2fq0i
MNtYDVN5B/kQjBxZqYRD+Evr0lb68B36fLjq+2Z4/D0PMk4KeUxpOOGMKLJdcdSwhStXYqNvxuem
uofwDq+mwznO17ZOYEZZnGTKh0SNDGLOdbctovgh21pO7cEKXQD9Pwv6y7CYw9I7cfVF+gVKU2ts
bexXhh4IgSNByKBTkZE0lznl/jNgN6csAL3k4jisIDoynstvgasB1dqYFR1YakrUtVu4td4Ze1IC
GLbOHKokhjeelHFvNT4UC6JW9XXBXUOX6uUf3gMp0/tkqGuraQLfahKQV7dZqfFDKDR2V+petchS
FgWMgWhByRQmfykC75O920PmM/jE/4J56hwF6nJYPqp4Va3mYiB7dkgFgHK4mJUPGxe4PdBpnnrb
Xf3fy2HFuOlpXc4L08A7P5r8LzgWCqGN7mF9QJmtaa6fWF7JtUVBELajD6IncJTgPUf7S+U4W5De
ghPGmb1TeKFqdTkQP1pBUe+WSopI2Ndz3DFa+1gV2cYonZ4uzFGSP2mjwqty1s9nZu9VOGml0gF/
/OpvsujCyAc0IC/er4p7IibNbwWHXyFDyVnCmqjaqN3NUJLqlK5y/v60otk66SCPX6/+PeM5OMHr
MJRa/9EqJZ+s6ZaQxFocwopRAPkkSgDr7NHrtGR5UVROd+r2BUO1/1lbJkuJ1kdJElcHfzO65sNJ
be9VGrl2Yo1Vkx2zi6bGBmTe5jkQ2nhJXhz3CMwgDFZ/aBQVA6luiSurAdBUtZTjy6qIYYolexYE
Wc2Z+2Giw0F6s9yXUFktv6hSPWMj9LiAoarqKCOIJnk3WmyqcF9ABCgNh2oB85rpTfpK4xDBzevU
CpKCt73dBVNtUQ6ude0pHX3rZ0ZXp3JW9DQzJjBLYnxfHYJxOevs7raYsEzbnsXVDDbOGlJ1xQvX
BuASpQtMK0wljs1ZMjfW9OU5ievZKrloc/VPY0siK6YfnkfE1DYRhYIxu85EasE3VljhGKRh770d
p6Bp9MjTp9qLrktSP8OpQfPV93m5zokMOoupqXkDjjlDCYEMTB+zlVXqs9vbQsDdZ7A3di28OVS3
sVGX1uyLhCy56p7NKU7oSZ4zrk4ps6G8W3tsFy080J8HWTY3ZwPXnsnoqUbtzKo8JZxUBthVLib6
NRoFf/zZ/Yzu9UK8fKdlttNA7RhcZgtyEjXlJYj4UknEuZcZKiSjGf6hywrpW1whP2u6Jeg/5MMd
tKJ+NVUclEibEhI3BXQqSKOx9SEoVkRKZRMjetDWW2lgWSR7gEU0iWmWbradaV1Dg4EiI6dOdCCo
7TANG+3bXeIWo1n+WcwXVtykwxrtugX7z6Sh/RuZCGVad9UzujFSgfI3qaivxzaaarCbcg5wCl+A
YzIdgYA+mHY7QDd4Q9iGouOwvsJr6b9Iq+Vb+MNzb4olkEgmVw/4qMh9d3l2wx88y/RkWUNMwnmg
a4G76/bmDTcSklJkHlFIuTp7j6EdtmYk6D2HH25C0BAwFSFUchTOVaIn89e28f/B5IT/urB4Nzic
vqJ8u/71kcO4xV03E+Rv4blWwIvzpF7zT0yaGrKLZMeytursB9h5vURYEvnts55b9wE9LEYmn53Z
4Al0FA6WjmeDggyNxw1ecqEDKn528GEzjgSqDTAd8lft0SefIv/Uae2di9cpDVFtsApYqLTbCDm8
M9i9H6lhXONDC6GG+ByR19icYTIwxfd+0UzjZV7L5R4hijgL/S6rXcyVrTA3pQeVNjBce+6g7tWO
9J0cSaBPPpq/o86b93QnL9Bm7ZtXKS9I9wjujNb7ScB06/+0yV+ptEJ5k45Y8fHQEm4uxfVjlKgS
RTCccfKmTv1fqNa4g8oovyEOraAtZrk4jksOn2jVZQK4ydrY+j4qpM9PpzSdL70VijK7PTXRsY2y
CwI248gR6bKTsLN9gU4NTN+Onflrs0ZZC5DmJr16xkrR8rBkUbQHUnZjp8aie4+oF0bby7LmQb5x
eAfZGi1kx4U73yQtNOOlpbpQkgZe56MgqpSMgU4F273lqM3wZ6mb4Oz8Tn319/sZSSJRq31JGstj
ssyevOWUJAuMJEkxEWoNLTnSTbUTZpl04LvJfCBvYilAKk90F9eBt29S6pbw+ccjiB5hoT+1x9AR
hG9y59SKXr6lDoWZq0rNs9eAABreVN3WMpf98TwmmjpsevmBJXhljVqt9wwWL5ZZQSXa/AJL+k75
EDAyBFCsI48WZ8wAPH/cFcVG0W9CvE4kxt/s4GCNd2lGuar/UV62ZNMGkFYQoI4flPQRF35ocIew
gmQJY5uWM3My4ym1FC8wOLHO/QRHuuWLaFJXcRJWpZDKf5UOShTsGXZbd+v4GTbzWIZY/FNGQb2R
plLypVOFdp50MzU414yyLEti+vHvAJ5PP1iSezNoVW+CC2te48+MotrOj2gm5zDdfDkTKGb+EJdf
p02z3PiVQC+z2IqRhR4kru5uzaT7dt8pLWrfSOBV4H9ZXj7PS+kdw8xOncv8p/FzFBt4B3iQOKNY
q4OLOXmRHEvyXqRgDoakPsM3T0PLjltVrWoooARQIJEUJVvx6aqoXYUz1rIwAREU296BjmAGwZl9
/Zl6U4iu7Kw07HUCoaF7+U2Ld1DimUIMfjFdoOdLut5ZdT96fR+5LcMkbjnA7+d+Q6yiM49xazSl
iI57aF9eAvtpZoCA/OQ+xN9tcU7w/xk6OABVENOl58BMZoUcLiOjRtyyyeC71ewUlS+r/o7LeiHK
mqrp53jfXQkU2XhbvdJe+BafdNDPZO3lF/RRYWkyjpwiE/RwlU6MVr2FqwzoWOi6cUcBd+QMQZQI
inQ8k/Miz3xBw3jKEUPhZMjDI/bJ+FISKKdN1CAWxso2iSpAWa6Z5fN3UJDwoj8wJEx/4mMSXdA+
zyUVWvHTzvaOeDyTbaCVnoiRvK5eNIWDeNzTr0ssYwfi5MtXyiV2vZgKA73AefpDnTc+vnAcRabQ
xPrjUqFeIWjIk694mlJv7BwLMOlGHeQ7ItrRr3PQgQuTzspN1bHc4wUtcKeL5xXizT+/lqV2VMS1
6p8QuP3gBB7+DeO2ETYHMftEM0Bibu/IEWvKk6aFAhv1AUBmf3R5gTcyXKCrteST+TEZABcrnlUm
OdtDzz4gksCwkL/TFDuHYAo669h2noKEW0Uf5TQzKvkiVzQ/9IJ+B5Khh/hb+Dpled2/JGltGcqW
nTv0pCGwDhUf59wenoW3fu3PUOCHythqWfGx6Rau0R/Oq9Uk3/4zO4v6JSv6fdkXFKnV6mO2eXeO
roFM83tg01/uz7dfvJn2agC820xPIe7enbzipoy1Z7jy+MqCm1mMWPGWWpNmHBjLVnB2eVFDtuwq
3DSoRZmcJJdymoLM8C/4i3gUkqwwV+uR/26nk0rf3oOCfHFqhXZo+Gm/mCmQpP0nTRSHj/WWkB0t
elojh/TvIoqm+VrCXvJ7dK2Ok1LT41XG1BSLmw94jMUHYvqkuvxKHxbRd6+DHsBoSRK607wkoGrl
GUZIXzvocbcKzIByHbUnkNkEhmoWmFJ5GM8VDFQ2nwZOMj4X2ZPzGBKCZwSZ18xjk8cpX8OrQ1bp
facSqW6qR8lSJ8bGmT92+eggNj+os6SclakCDuquPly82Wq4ujpw9S9cady7AK+NPJ61LeCdZdra
c+if+1hqpqbxFIzMGkKv/EnKfsyJekZlTHUhzV0oriL/F/BeiIYE/AKMtoc3kcaGgoOS7+U5xa+b
D8e0p8mK1ks/HEK7n202iS200b0D5WKQVL7giWpKk9z5tGfA/H7UxXfNLGre0XfyTEcD268mSJrO
jWPgi/Ddr/ijfcfC6DIqg2QfHLgetQ5bnvdK5gYfX05WuzITgoZhYE0XtYidLvIdKinlcjHLcgZG
8IcF+qwK83fv8yzfJk6kriR6p03X5e2L609Uz3Muh0Fz8zG4iud1Io8RmTSHuWpCoufxdV0cGeOm
s2N9a7nlAuK3LM+7Zb6po1bSdukgBs0pFKulSyzt9pxFrkDUxSGvGxl2iAqIF4x2glWcN7hB+zjc
EOfgrvIOi9hgNJdYQOC2FRtfiBrhAh6xl+AdEQc8lXJj9PCbqSID+SIZWf+Hh5Vr2zrN7P9PZBrd
aIO2qOpanmraFvnuSCnCXbpMsi9PxUDlq0qHPfOSO+3SHBbhsDky15hiJHMJX+EsI26zA0gKVGB4
qK/cldvoXkWOf92cTn+JEoJFX8Dbi9F5W9iBsC9qQAMVkP99VIddI3BQ2uEvuI3R8ZkrYxv0clTI
RbDGiDvS2BzaW8sCk2GE17/FIitw+1ntaXsTGLtlL6/qT00EUDV0uErF2GK06msCm1S1s6v0jBgX
yvc+SpalsYtsxgSZbDirpKQi8do+dAuiU/O+1hm0z2o0KEoYvrMNI72fjluXK90lxjSPRF5Ab44y
saFO9ssp75/YV/j/HBA+1QGgzPydsvLjVOcy6ThCRTkvFAdJhm22fjGZwuQaj/nArPowkX+8vhRV
tsGTq1+fH81100vDCKQh+gGTaK75GfDdKrq4dPyCTQx1GgQoZWvj2ygk/t8lm8ZY6wIg27mXXuud
/UbdRJibnVfHn7NMHPGInRV5Z9dAHpB6VqJ8io+pEMY/wQ/2FMzS3EDdl82hKKJnu7OohAeAgi0s
WeR4cVSYgkBzCndNooATX3tOqtsk7rs4/jHn91H4oTaKDzP+XlO/Rbnzo383ct7ES2Ee31pKQsBY
yDdTGdlSezWo+t5Tz5ZdDJHk4KFYxv4qkU59nqUbLzcprUn9Vu+Fq1bBGlrU6sL2DubNJaSuxQs1
q5VPtIuLJNrJMAgPk/8M+Bqq1Kii3Rt8UcCrTTLj4X45f9+3hZjloXDyYDdbV09x3wzIvhAZatGh
xabXyXeX4f+bvAY713cOa0xhYtHdwLQXivFf+VExQTPZ2dP7ugkjQQg9IE4HrgMDBmzcvpP1cY9D
cBrvFDpNUpeQus4yhQVFQ6/sMbk4Z2h7kwe6niPhI7cJS5iWGgBIoHGoCSRWkHry7gFgevSpME0v
RRsGc8iofKdGhsFVlcUZNlm5DUHH+bvXz9GA1ThTvLeATZJ2KPXyhqBhedGZqjG7pVWCMXXrX1Cz
UjbCTXM41crsc2QmFyWInNHki7Haqt3LHheVWjHCaTeV6AsF2A9ddE9RtuAz29BhsrLTHTcQvPtM
nW9a0a/5KPEXU8Ji81icF+jQwf5qdRTzaD7eeloh7cORUalnlZgfEy/ICQWsZsEYBxQHntfnzQXv
B7ikFotQsWxnDTzXHTBqkm5kuhgBq2h25gDavBAMV+xkp0kMEOXe53378LBPy/whlNsdrFmj3Wbl
5EfZUJDByk0XEbmKyUvO5sCWt/Ax0Bw80enSR9RbO2sBi+zFdB2dRBZ+/68m8NbnIJys3OxvIgMi
4OPaIR0wyNYZMJgX8fBOPwhwNNz4d3jZu/g5rv5ek07qQxRqMfXE39lfBl08TIVgyVt9VM/ZsMVf
8wuhwWZ+QeViiopkqo88O3uTzi51HmnJ7dk+Dw6BvQJJSHt1MCWH5tz2jxj48xqpFe7AjyCJpk2U
CnEbtnubeCDSYZfsP3qBGGSGhfEAF/ixTt7LBrWRnGbxkq1k9TigI+ccl1psztfnpjGJr1/hb57p
uIqOM+eDUcHXRI8MH70NPdFsOCGscT1zUJygqm1+nLcn/mIlZNyVahWfG9Nb/vXkeqlDv6CxXSpk
TE2YNjhMFHuOaj/2uCUqglw9vZaBu/iPHoF5sUzMy85K8DCOBob0rb2yu4irw96/4YArjvShLlv5
j76ma6+iM6c5LJfUsMVECnylS5wENrvWYG8hbksSN7jfs3kOkTbpdK4EEs6EMdu23R8OcKEHtUz0
aXtJAfRoFMDOhjJPDe7b1Jxk9AZzgTrWblfC1iD4ze/UUnUcic9c+pU7nZ4q8ybd1tJn+cuk3wCG
KVO7R68md8o3RvP+zz3aAm4a76O+Mx7U/Hj9h0Zsa/Zxr9jJ5iUEpe9PO79XC5eHT1sW4Jt1sy5C
JyzWeSOQQ/FESw335V2gU4MDFJ8On4KhT8l74BXnGzW+nTUWqsdEF7ibeBZgDvfRWkKqIKRyMsNN
vNc1NN2KT401thjUpwKtcrSANi3iiWB66mUj0QiLDKIWtSwWsg8lhGtbNJblcpnn2sSb431GtvSw
/Owvruon4R1ZfjnboOq841fUzC0r25+bmwbu+N/aBv0q0n3T524W3y8BtlFLS52BI+hLkYb+ynLm
Okl4VjQGF8WUAb47xoq4VPRnsPUoEYvnxWU9VXMBuORLcLE+YhwhV1Lgfw8euOulVRB3iREP9W10
8CGuH0Yfp31kTSE2cFS89GS3Q1KIAAtdTO5+vjpjYgrMyhE+WEw+XXtmQ1IPpLShwbKhxjHgVyPH
n+0y7gZ9m5ST6fSAEZv7JHzhRZ1R9GkRj4DxPTYt81nb7TI8/42eJwk80cVC6wHT5xRJlrPesUFB
nPvPpNtGq4+Xc/XuSVaofo2ZkGehhQHv9HvHvSLV4pn3qSCtg6XIS+UCRm6xJHhTd2k8M/VBTSEm
GmLlo4BUszbstBbFPMg4lQoM3JWVfpY7OrrMKKip+EZHs0fiJaAEpssayjny/73PiSi3SnUC5F8k
eXdL/qHRAb3To4/G/tjbil9rsKEo6fgdQwuTO09Sx5TCd6YAW4FIRr19Vgm43+wHox9Ck52njoYu
NcGYfXIhJKjj7i1k2vWf6Cnp5bZs22o+CLTrtuapVqLiiv8iKb8SD91HGgHX9eElps9LIW/XyfNu
LaQyAeyWw5xrZQQ7+HRI1irdwu4IG7nH6/2n78s363+4bgtoCTQK7nRxWHp6enIDyfNp89uWsJVY
8zQfU1ptRRsaf2YeVtwS5GGHxu6qo5alWMYTD/vAv1zsCi/npj/ca5/VF+k9SWqjP+VVP6MLMLil
J0OJooD82TWfqg6XcatJ03G1dn5J918Tsuf5FjZlbxIg6yrtqM1GhNT175L0q3ZLOgrQkf9BGRZ0
Th2BFyeECy/SMTfyEdwtxRqzA91uoBHjTF5k8ONOfBxlUDbVc11FzLoq3kkBoVAgeACM2JLVNnsi
lMs5y1e0FNNVFjkPLAD2ZGy9dUDVfyh+rsLk8/LCQZ01gXirbQXLaG+gDpkpQDx2aiVyJ+L+xMyp
L49lJkcZqL+pjZIszRgfuXT6qd9EN4Y9JpRp9124C2/MnnrDl/Rnzmanb8zedNMZExb1GSZoh+GZ
Je7YP/8d0kijK7loaw476yeLNen4yxJitW4MrSuOWPsyC8KDkqVI+1PszjWI7aNMy7MPD9nQc7Rt
QzwV5J8UMsmk7Han3+DWhQcMglfz1h+GeGCZaQ3ZUuiqb7YamEpkzKdV5lH+GTHezicq7pzBUUhX
8nkByhgq9EazUnvdULyS1o12S2uSlm6M5iR5QrPniYv8xuZ/CsFF+LCaDvZhrJ5c21wAQIp825FX
z1IxQJyBmLZ6Lx7ipzwLeYhwsJwmK3pv1LfGfqgj65xS40km0PFn8tK3XNfXmK1qo5rAUox3BZGy
CTJAz4cA+DvpDWoDr/j4Hd2PL0rNtABDZN0GzdMbFM2v71jP6Jzl9tN/JeWz/i/dAPnpimChVUkJ
+2y16VKRw80YlrPqaTSnU8uHpLSUegdRlIAAbImZD7WHXUDztYU35Ys8YBkG3IjnidG6BPlQZlBq
8NBJFOyArboAmo3Ur0Qcw3yYuyjQxDhVev8ETb+ScQZ68YgGvBjWYxH8jsOI7k8v8H7MhaoWJup/
YfTGfVXi5DzLFe39ChGEVHzUG2lTDZlqvLCIlJc9kS8ljcKhbZfS9vvOx0MKUXZQUn40GXmljIHG
+sPZfr7augksyuf298kEE74lopNJxih1TkEFOZNlF/M+PjzQazaTCKA1HF43ljJM0XzjpeXBcFGS
ekvU7TyAg0cpUWo8DUm3N34qwnFHiFxZggqiZMZL/WCH/83Jh+hOGA/2l5NQEZrKXynCq4YO9fJr
cg2bM8Ed5mp19uUzl4EN37bqJQS+wkrIJy9UAqKMe1me/owbWs34wc4aHMqDsMIvN/bdW7MI/StE
m74sQxGriyvrGgET+0p4/peffrzXfVOjmgjtS+6jDVDd7ruXCLxgIP6K92IwdF5nzXuUC/VUIoQX
p5EOG2t4jHWYXooqgc3asdPkQzaJcfm210vxbTeIgU5vazGmK4mWKTbfDeDVRyBQfqDhW0TcxoTD
pCoGDB4kTfsU3NKnxXHtAHNL0JBUFDFTkngEothb3iR2EdScG4Cdu8GOlbrOwxj0s6IaJgtoj+6q
QqlDXpeMI+f0SmwyLjzSKYgjAgFSksvbVh/WIGuUPN8E7uqGqN3DAhBWkbxcylD1tW0avR9mLcVq
oz1Yv8z8cR8aFwNJDrCJWMhvqUjkp+ROCjJrnOm3E8+vPtKb92eWnT99lzOn4OwDZ0yUXRcPiIk6
dgYe/foygS8bIGky7ww4LLFhFCd2gYKpuqakZvrU+YQPnaGSl4WxFxF+C6Eolo2nEFF3xu5j80/I
nRktDATqMRfwudBdhWCwCz7BMwGA7NZOPpclqcTZKNUrpnvbVlxDB06R2YER5kJX+s4M/uj+5A0+
CklMFRIM1V8n6FkTbeDBTqhyhO8xx3YrYaKtZfQCJmoOxmCoD1ugEpUIvi3nVr96rdB5efotGvCi
1tTYwzpzZnisN2yWI5EUUzEbu0KVHfIuRc9FNw9WqVvmT8CsQMWHX5G2CjGHErey1ku6uPflSlFE
dCp1pncfflsE20NW641xvvigAaJYZJrOVf/Lf9GKGjTe1XKRmrok9VU/Aac7weShnjKhrbtSkWhL
WulAeES5eTAbyPmEeo+TByH5woQv/ugDOZTiQWEExbhV4czwDSmz48XjLWA18fn97BQTEZLU0O1x
alKsp6TUOBOAgv+v8d4SJJR0WHsL0wlj2yoIk3gSzgv5E87mHg1njdI5wl3sAaCaArKGXlK7mCIG
Q3oQw6Yg47K3Y71Sr2y5OLY2KUF8STs4QwsvbRfASDoDmOcQAt1LpG2wV4hnToEUnbhi56ka1OmJ
hlau2vDAU7uObMvrcZGPO99cSnCL4ddVWPbDtT0Edw7hLtg0p+pKSARZvKHWDCAE7oSu+sYdZxNQ
ARo5LjWoWw5y6zwmpErMa1BraERQTE3qTc/Fu4LSV5xFx9hh2EFd3gyEjZQBc5j0dRwSiKyfCVHL
UV4j8DrSxEHufJwn1Z5UMDDKJQSF9PeXsyAMdCaO2lIz8gwywhlA6i5eVT64RGgAmY/Mdpfx9L7P
iY75Fs73bUFr+82G/lgNX1Z0ZsAp+e7XDjp50MIAFweTNqTYzg5t2QB4e50YDhnOOQ6eG5XIDgcM
kDqHPBkNxxpaqN8Jq4hx9o4OP3VPlCOpsSCShDtMyER8DK96Vc9vhHjdD09FMbfoJsjkOjTcpBGs
JwoYPDV9vXK9EX0bE55EkvIl8gmxkN0hrpYlTN+Nw1RkuYCS0d9DPPOPZdcWs78cUWEFeRcnGGEf
+r5wtUOpufiWcXEm+3f3D9o8HvQS8+nzj1WPkC9FcoPJivXw62e2oIT523+LGBTBaIkOeGPGW7ig
XGHccTF1VdlEkQzqAjx6wOkSi8PONiXwCcAn+9W3gsULeXwlFZVLnQ/WY3x7JKwgE6z1vTrbHtWf
GBlLCIFrJs8u/gpWWv1pRHYmsf68/hEL3GiEhQsuJeAjJ5eVjNk2jYiqkqwP9tGVUeIqAynZscIc
qZlaniNalCdmtlTM6oqe5OwiW8mt5EyOYsgou1l5izwxC6ZTGJq+X2xSn0AozahH+/N5BlS2+2nF
w9YJoycungV3deAvhfrfMHZD/lt8o1LWOPFixFhI+KehNvn6xSYEXKJ6V91NEoVkYWDI+7VSoNYU
7lnBVv1Ir012dSBo7AzzMaAs0WoTan973r43OnI5K17n6Sj3gsi/Tv7OnZ+Y3TT5XRFIMlG4YmPL
vKquE8FYRPhiLaMCdMZfSi7nilSVMV+DlfuJcIrp7gKrq3tadGRhir9M4eiQhWGU/XX6mIv+ZUXk
LerickFiZItJqngfOaOLMmF1prugw/foVafNDKjCBS9tc3o5nGgCbbwK8Dxzknucz4SRlPTbg9XY
vwfhsbSzs8lwAP61NQ+joPR3t/3w5KW3KIIqJnuxBna3sysHSG/ucr1uUemS2HZHsX4Cuycxt37V
DS83Ek+Jbpb06rg84VvvXBxZEYP1QUHlAP9yZH3mQ1rbshf7tUnGlnY3t91eZBRnTvnPIylW4wam
ksBWrfSZAu5GlC5z585TmZ4nqNaBZ38aK0NIQ2Izv7DvWaSjQgxMwegq5V86YGAwtPuNB5MLdwqF
PZG07+S8JIC0FdxeYOY5knyOrMZk1oiYPDjcNprFJyZZFRmmi3ZgC63Uq4fH8F4O6qqKurENx41+
1ua2/56MRJoKJwngGU9A8o6uIHRADVzpvgUv3i0+pLsq8eWDlLadBNpLZyZEsoZzLxLK/cROLYhw
O29/oUSDHFMVv5L/DOvPQoHUEaCZDXU/YaTCJAC9Lj7PghPe2Cvi0stQLI5JEfygmfCeMeZsxRvD
9trlDQQ6rP1hRfs7JOIgw9rz0xrgsI1lhWy1UsvnSoRWUbViUdVPi64Ne+IdnCBAcIF0lYW2N+RD
uMPCYVvAommTxELOaBODJl3kTna1oANiKwCAiHZavkwqUctLpepb6UiqG3/wUD6NKVB1sa/qYVVl
f2XQ0G1pArr5OD4/s1QLgiLxzhbvOsMnHFnnFgUc1pi3/duwr/IkH5zLPlHPAzFKBEan9Ueesu3X
X99ThAoGYNpLAZe95hm5K1kN/0Lihh5nP3Dd7YTNiImRS/rydVM6A7k2+MOYTMEVXBUGN3guF7S5
UoUaA0aPIafHA/JKfgpHI/uxsvktUJXWNqmgKhidFdGHDhfdWQFWUUIjQu+rxA9k1t9k7F8gPZdA
47dKAgMmBX4f1QqQijTI5ZAS+5xwWEaC3fF76uTN/IBa4VY+lyBfyAtqfbNxZG332ujOVOgRJPll
SuKHXEuWNEhALJPbT+k2CQXBb+C1Oo3vLhC3dxZNSWDBbJoZLO11hxMupuSFBqcr08P3JGjRHF7n
Ucr1i//duk0yj251tWsr/Tb7Wp20WiGpCXkx/Yly739B/h0To9r69nDwAva1HGbEjag1niW1UBf/
r7Z6py2df7cSN1hw6B74c3y5MGtKEonUF9vzVsRB3jLVxVk7dcORPppRgOcKN5+ILBISYLwPWfpG
Y4CXgs6iYu62qDupAvEej9fi652Wk5pjCyyRmBEU6v0E8VQEqOaqSMFGYOSfZyEQ6YrZ4O7L5DlU
pLk4Rg116m5PEuu2e0+Nz4vA1ONcJYkgl98VpWMaHccjMyGx3mDBhABfOkW2GAvQFr+6Bi3qSX2D
d5uP3P2dRWfK8TupruEbYLnLfhAjkU7IqBrQULH8iDShyUA5yoFxi4x+umpnsYwpLTtzO4vgpGSJ
6A5ouWbnPA88TcibECgsY6aPh7M8lcIKVjnLLDhqYIOq0UI1KoSc29n/lj3CeqfQJazVA5pxELO5
xuYLfykQ1QoaGdFCA67I1eBt0JqnaCzVV0exQpkX0ubyK+YgUxHlrSmkqvpJz6V9ANo+nKpYdDw/
JvfvbIHD3v0wev5xkX4HB8qRjX2ZAH1mxhYFfOt8bql7E5icWeDx0wK+5QNrDQalT5Dr2RZJgFp+
+pMRPsa1c3o5/miKoxXCNukaeW5q97YoRO0ihrn/W4D22kezbE+0edW+ss2gf+HeiPbjL1p2hQ9C
e3wPgdW/2845JOzzmbJVhNDY66bZBQiHmrQqZdTUhD92OCL6CGnxlit4HHwUVkfN0mVhdcnh1Hk4
vC8DVQsbGBqaa0pRWbctrpqjT1YPtTGUlZJUonaOLJU/2tNgcWplt1Htz+YwTsYdlql/cejmlVK3
pBJgtqmYtlFLHqK6K4I6SM4xheQ/99YzckDizvVkMwdoEuWKQV25+opQ2Eu4bc4ezFzyjKIOK+9q
2bmNdC+C3l6fijKXhjLdkRSHEdybecdUFwMu9dAeL80DwdQlp0ycsfiuiDWxe2wtJO68tEnBDeLa
23ZNCd/5Ho8XIJAj0UPK2wTAEE529S1kxUPPg01/b9jMoaryJKyeCZcLlcJYy0LebX9XCh1W7qd4
hyNViKfpi+/RwK5xv/HVdN42dfbiVsFolK8Ye6+3BPXUnvGb0jrvvzNZJTmy5fsGKWt9S854wfNC
W97XGuueINw1CkraKCoxOhMyvGYAEeYpveHwdD6w2E4wkd3dPdIGK9CrBvA4Y5doqPCPtp1R/y8h
ppBvdXDMKYnsO+KwxaSFdidzeRnbKSam01NVOuBZ44CG/JUGaP8e7EquY3+vlV1OZbh4qhSv5AgY
AvQK+amRiUpqs1SopjGFs8K0JExSV2Yh0nwH8dUPGHyUTQ0WLP1FG3HaPlgMbn+VRWS4YnxsnL+u
ozeMp4pUnVE4F8SaQHx6EAob6Zx7a6n9FyULbGz/xDrHIgFCZAbTNvLtcomvuhKAUj3azec6cwvX
NPn/f9dzZzMPqO9oIHgppX3LvsRTUj05r9kOMyc8vWSKcgkJq02Om2hCzy2wc8TbkerQf8kUmdrk
fIJc+u9+8SXy7AXN+vhl0oTAGiiqWSDPXbE83jk9lhdekkk7V5H2nQzSpFdoWPG2xHLynL4Hk474
YVZbunn8AIB1C9284O3tX4cSgrieiCLlMzfSm785aR6uEbw9tjix/O8/ZlWaj5Ic8OBlRKYEkjL3
1uvo8ofLt5ltNz6/ck8urriaLFhTD6hMgW4A4C7qH9VQRRepktT1r5jc9z98YbsJ+iwkZUZ6I4XH
s1x+PuyrL2kebILlh1xgVqhW2Xx9DJMRpB8Ot1LqeVfDtTu3n258V1+vRcig8g0L3pyYrrx/xDSc
iBO8XP0ccwmHetUEJ2AHYp4Sa4+feG9OEfTjvktv0TFHgahBs5thveEPmA5qGkr4OJRxbtEBKrSZ
G8LKvndvhWqInSZFMIxKEPEktoZ2C3sXJm6kqtUYiQ/9ZMUS5P2CZuluKByk0+H5BkJVW0SiAaEE
W0Prn9C1q0ekkiyXq+zgB70PWmETxufyTpLkoBcz7dZRdt1Z4nLectu1LbOhkFu4IIN3SRVGLIEA
EhFo5M+L3MGpodn5rAxhJXd1hwRUBfS3HaBlGOENmMamZiS2l7IIrO4gs5TDRJZkSSK9TWzzfIwN
boJtUb86GQpwxZiu1lqMy/QBWrlHB2Jkjs++8851Hr/PgxbE8i2aSBcVfzBy1THLVqhNLzBlbLAn
LgXjivVoq1vsMkktJRZpSpUrUM/4x2tYAtlK+KP7CFJmDu1B4KtyVgKB1sMmMawvo7hYIPKd2pQW
jcp2XucP2kIQPlytFsc7vEy1lNL73SWTD+AwSyR0plseqZgvyJJCHdopuxyDBK8hL5KbzBLKJC6O
RX/i3RD7ceRO1YtE97z8L3g9OOEDpFK8aj8XSZgvUXVJDocvEc3/gZmS7hnSWJ5feULuXtdtgrKL
92DseTXKhEFhuW6oTxG0CrxEFibyjQeHrseWyaIlrCbTSRPvdbPsApCHR0NYg4xgUUgHoH+aCC3B
1Ogrb9fv8ciuNdELKsKoTYzR+XOyHCYGICFLj2FescTvVnz6Z68q7kSuG1spBL4o3TaCAkDEun4e
mzX07lyYw4VIi0E+i4EzPOkoHshHnOKE+PCG1UbSj/LSJmqN4IdBowBeV2L8hWVdKWSfrYCByt/w
mvPEKEzZCgVIO666iMh2mS7PbaR+fAfimYsYNr+d8YUC+K+0xP9thu9EUvb+FNO/2GP6EBRknkpr
z2po6CEhSWxWLofgfWVhV4riOJvZc974bqdxJJ4qs9kJU+Lf1BCdHKMEsW1Xls+aY9+XBmleE2WQ
aPRgN7QoUGID5Ch++EEmziM36tXJypz56VEZqHfCnhrk1cQkwcz2XU36WLLDXyRbUYMNrvPKOkKl
dZlL6ib/yrWsGDoduq8oatiTX5wcnrYpLZpKScNzvR3GpahluYOosBeVCQgZEH0doyB8bUKU+wRm
1s7e02GEHr3QB6qC0OT/dlGw7ReyMvIW1reTlodFAv1QgrpxsYF4/HhMIgTj61RD91BXsSu1nqFb
RiwHsGUdajOY9MIT/QyxRBFPJN6w+gVN460/ezP330OPcoXzB4QwEFxKI3mIJUdGV/xWfKdW9DgP
WfpIpcbGsCdrYUAOGf23ARi6nhZgopU8EsNohTFbR290Xa5k/nfHYteRGkHw9dpxfB2hUcbb1PLQ
0UyGC0mDgknWwm9eRpBILZ+2dR+4hRRvTPwJP1k7To7WguXp8PAYd2y1nHjAchEN+UGtB0+x6Nmc
m2iA7nc/9ymoue3pVuI+/KU5ijUeM5tiHi5LGclBNnPdZI+Vs7lSkD2+EmsqJDcXWb616Njf9yqO
5SRJRbo6DHYRo+ZFue9A9YmmUunqjx+qoM+E/8HcBKAx0TTLZSPr9+bqu4W1PX+h3uCCZQj2Zaav
05c2YvTFrLEhF8A086I5xvmIDjbzheIFpQ8DeCjQSsRvOSUm1V9lHGEw9cCRhw3lKCuvxaD6EVeX
UP7/3pSI183cozMHHjCd/iymtHUpnl8vHmsIYHooRudGmsn7pzn72HcY/IpjYDJj3J1GbGNWw26/
ntZIFlR7NvQYzcsx6kBQrcst8FNesx1NkAZy98CJ6ekfETfiKo/Fcss6xUo8X6KLveqOHf0nICsW
yO3vKRW79dG+1YEX6xcT5ISeVGKW9Uj4We5UfKC60+oZ5K/0D+xY5lid09tRgrvFTPnSOxc2lx2M
8aw0aXbZXQ8EFuVnvTI4xoEiMl+MKQ31UTE1rjk6qX8vyMr9sG1W04g7L6sKENjSeUIAwlkvfp8X
V/paSBRlSGwCZtDQKNOMOehIPph/SlD1zGRVxYDUGe2OsYMDRccB86Jr+GBe4UZMcrZQa4soSeLd
cq6lThdrj6QcsEydZrq8K2WAM6GuiZAfOVGaXsnzEjh99MkmSgsXj9ouRjZ23kzwhaNvpFUKUvWA
bvm5gTo4RcVp/aeqn0Ntd1ea6nnwIs7UrSyqguta0bHCgLz2YCC0dZxAevtSvV8tbTz7QePIUMny
c+MIsTfJZ7PK4A7+v7N8qQ15qd95utzxKHHj4hW2nR1jXNgkFtxmFsQPOT5rvP3qn2Cb+wEZGS4L
ktFP+1g3GaDh7uawa4t675mk1Gw9Pcyt416dNDVpJm5sQSBRn63PW7P6+RNmLMMS3RjZ57TNQHck
dayNZrxO+fK0ATElsfOAyXz5aAEAwDcYEjQKSNTMyGc1kujHxcMfvC9a5cT7Nb8nYjT8P6URfHF7
MK1l2UQfgyIfUZ8BmFKsltFVTNqSWhPF+pVnJRg2XMsmA8m+X1r9n29luJCXeBuXhNm7WaGtosZD
YShuTE6jbKlaj7pDLwDDjP3Hi1D2cX7OyV15QIKoOms1Zf9aAQx849tkBC47MtP5qtzSV+K1gHIF
8DgVbYYhGjLGXbZKvBGrWoOkj5fFC7R8EJmAsO7cGBpqWMjPS8zcOPqqI+jppoeoSkN0gkaJRD0D
f/nGXxKrIWvIYhvgQ5yN/vbWgZry3SJK8FEet9vVA20Jdw3mVQVMP5uDzYKMF1VMQzlN2S27xa04
KsWu5AFHOENWRcwe2nCm1bECydNOXZ2oz5X52FxLDoirlIZoL7ntyVwxD9B/HJFK2fi16Pcq8d8+
Jx9JKr+nYrrvCVF/6JCitfhLLf13dOHcIKt3zAi3h1hjyDciOLeQaRyNXhsdMuvEo3XVSXvepvK0
4DpL5iFt/Qr3JIZQ3ZvA2wzJ5J4GdmKlJF80tvzEB1xyxAYfjFGiwhymkBTssKN6y9RJMuCAfwmr
Wpu1u8l+TTSmxPSTRZSYzRXjPA33whpCQTtpLcWf5mH3IjCPlTd/ZKhK/VjJrK36vU4zxYKSpQyX
84vpoe1G9Fn+twehb9cRodRWthELCUkDRg5H4mclXEIRxCLjJVIaFGs1cT/63q5vH69UNn2HApDC
KfgGUNvjFEbLIui3LjQhuOipSebJw9G8Exom4jQssxNCKOQtx/K7K7Jnlxdj/1VHyUIVYf4fW8uE
3aOPtV1D7Qt1ZywwL8hJIA2uyiDNvBz0aRhqWmeNc/qaNLGk4jxKmMtKqVgNtmrt3CJDx/Cc4ohn
9H+CqL/F/bJM0xIPX+TlEWDah7+19zYUV8HCcWaDLWtr/MxSF17VXUBYJcQZvoLF8oKemU+ncuA2
9VCt61j6MGelBEDXGtOM94Tb+7osURuo9Pl49JN2QRuNj2ROLDZLQQeMWON6+w8sHWsC/waAMYFg
RvN1o3eFBRuKwz1OByL1erMn81P0HJ1rLQ/ZU2LO+Iri+8O0SngqyFKvFw2+wLMIQ1SoQ46hVOCo
xwiCceH4MnThTLP8JH7mYepNIoOEARwthwsX0PA6gGFNou7q4umQyI9YKnTKl17gtV5pVHJARXOX
nLycMVPB8bRlzHE2nKfrqWd1+F1TSPKf1TXxiXXanlEbUExvLHgWVuOtkxm5s4HntckQGVAqHSBE
Klpyys5q60HoMSQJJMPeB9GryZUbPJpyj/LAt3ol56DYuuHaajnSl5/LGWSFa7Vh5yQ7ciQQ5jza
bkr75CFzCuqk/SghEfj4AKFJ7QDtvo9+rAuT3qk1ZciTBc0Y4o2QrmS01DMSg+fSDarxToXPQNoT
peRWmcj2Hh0f6sZub0HvWq/c6D3zSL6RfSocHkoz4QLZC0ylrkdqJXCcquAAbXV9JcKMklgobLoH
/DNhRp10zcAyPjTAN8bRaQ5b30xrr30FTEJ8aQHGkfizfMen9Uhth6HznHlv0ElVmIK3dr8W9wyS
CfgKSTMLwUgSK57BB8sKm3sruIvXc0v90hpGuyHwStuttPFEpuCAdxdV/+5NWWTrQ7bIIy/lrPlB
UpBl9xE71QESpaYS6xl77+khYnZtj+51+sMwrm0hAval7zPAC3YgCOHiuBpLl0Qp00Wl9wAR+xe1
EcyRj+1NgcjjaMxJYd/R6WJlidI4E4WzyKHlKOBvAmo6Yjuf3hZrN+8Geqd26ZwSxbrPOPNL2Cja
xkO7R66UJmt19WFwXWJAXtizBLcz1JmPrFAT326kBROgJIH+deLq4UQtech4UBFXx2GXKaRxAc5j
mkiTDJbApLozGQiKE30d4mUfAVHJkoPCG5A60niu0gCVXgU9mrgSFVl+qyh88IaQQmJrEzdPTTuo
1YsIyIzRyae8x1Q0LSSHJswUfTmyhPtyG9Cgg3PjAwyfaX+yp3QGWCWZKs6yqsjdszpLi1TKXSXx
slzF8Tet1ZsMcst1ymm6jtNRYNuNvO/h+8xjdmScOJigEPbBQLcFeQonXZAr8jlMI+AEXFX61evi
yIuVBGGJ1PPMwW1Uar1AfIK0phf1iSP3Vt1+UraUGXuiHcA8O4pjNhgVKWgpY0ncGfnNWgzQh+R9
YUWV4tTkIDxmnw2DrfrQ3iUybyjgqVQCwKIlrcSCezbVBTCxgL8l3kSruCSr2mbgGRhswSE35f5T
68Gxvi11Igr9h8sIPFpVs67DCK78tdlX4ffJg/6HGGKQmbIVXmyuOVmxXLdK/khfnxG5xe2FI9RB
t1iF8fM/qs4U3UsP/TcUStjYyE51j/6YRDs2V8wlCfwIGhz9JYpMT8sbkNPO6/fSR/Ukbdux18a7
JsbH1XbTY+0yT9UEVl4WtQGHakJDvjk/UVxFrRP7Gq99yp3A1DxaaScqWF8wcYNwpuuJNKq7uanc
e5lApMGpyHclCVjKXK0wIwvzYicuyuubum4iePsHz5U0sD0dUbOYLiBZOxQ1VE6NAEBPykAmO9FB
Pm/Sj0SvhhX5GCxgHMXusG1evH/qvlWUIgxpgkx02i09r4vbtW5hXOsHCfg8ixbSCOxhRp+qGpHE
1leE1DzxlzhE1Wo+hgSuazEU2h09zckdF2O+8Us1PrborJkFETLyOFQ2zgwXyZjZS/JzMFx+V4OM
bUnzlsrSUsPBkroRxHBvMRirwhB1lX+Ugvpc2l5gJUCG43x4skOow2/L7CfMekadHoignlqZ3iKF
rIvvzWESgIK10Dkc8slXrn0aYJ3C4V7MzI6a3alkA2mfNFxBZfNR9fuWrmZCSg9LUnYjd9f2b1nF
Yv6axNvNKNnGJYULCGwQmQQ6NCLv0wUaPeyN8lKElXBGoAcNgMj7OtHuc1qydOdnNFOQ0yDe+g8T
MriRYHwr4whRSiUTARBmLq7d3Q5p85bg/HCX4IaFMgB8hBzP7rv2FlquMaMeAc3MfVZZuBzYR7yT
sn02+2w4DIdU0PJqGOHVGnXTuBnFtu+qHT+u6kdSBcG9X633xSYwN0FRPd6lYCn5ZzkowKoEPy1S
sstFqy7VZD8akU/Ew3ZcsTKeKSLIDEc5yEPHjBkM2chcSJgPnWF/k4ImYYuDdPCZNE+jZes33Dvu
AnOsg2lSp0lPVhaGzvOCtkGuF1P6V2A9JVg077VZct6HhJv594OFDdXloZIto8aUrcysEwOuoQlb
xJl7wEUCGW9p8NkQJ+YmdLo8B4mt28KMjJymSWZkO1KsK8IBkPpc1uMYBkIae2F+tNdqoiaNdH2R
vAW/OxI/tqUld5JhG/alb5CDxu4DS0dD7+BHhhMqIlajpypVa73ZszSmb+BQlL1zM9RpC3ZQ21GK
uoXZND79JrDetHr2IsrTkm1Bc97G8rG03iouXCUpetvSr4Re2BBl9/pq8Z/cYv3Gtj0VSsS2QzcZ
IAnTjCpnhJxvgdWatV+H0BpiFj4hj6njV8iOKkCClxQHUmEPzDG8Rtwq70FmKu4uqNmQskXn5qrg
oUbg655q/dq9gJ8SO5k+33Awh3HHY4KikpmRW5emKgW1RjL0aZM61llnf/jQIeuGwlvmm4emGPb2
LbY5vrSxzJ1PG/2Kb+qkyj8Ii8+zJovlUzqH380KcOopnCLOhvL4L6JE7CJke4b4pGw3CfkbLMdB
xZOLLerLiFwwVehbSKqVAZer8FFyP3PcvTYIqdq6xO/+/GQ7R8SRPcDF/LD2j0R4ZmtWLi3dNHzH
NA5D0mO6smACYyIh6bZIw55sJRJTTmnAz+EMS/AdhC8ZHRbd1q0oUDZ5ANdnL8xpHOHSmlJLTtQ7
p6m5J18prKrykc0laC8knGx5bEDosD3qywDdM9yLPJMKEHZdFmeJPmLQ8x3jMYe0YNAjpZ8can2j
IVJ15uobrLUdj/P+bO6+tX6h8Q1ED14zlzaUv7hjXwhnINdiM2HlbXn2O8297iOsmORLS86Ip7ny
q/53mqTmiMKjQX61vgO3Xz3k+TouhzTylrGME+Yh0ZSLpT03BDBmumzuU2Ei5PNviO5EwRbQM8vR
WyufmNNIGaCjhZQRwwee4f1aT+F06ee7s6FZMl5TRgrreJ+pJlIhkm8mmu4X/FqXBQ1EFRt5mXer
5H/oSTaZEXi/S/fA4JvPHqC/rRLXsQ8MGo9IWHnsAsnjHqFKZoSnING3qK6DPgTvX0h/Gb6wDhb+
zC9RWB8yJf3luxIM1f4rSK39JBuiHSMu5IO6ztuUkWpp/pDlpu/u1cjT3XmIjmCH+1hlKUtFAiuM
a+KcaX2/1KWNsL0gTQwbr3nEYgn/vXECq4ngEudXL+lKmEUpubJEMR65ws//7dLP8WN31fXqHp1S
Q/pxqFKuPW75+lehY3yoke5lr0vplv7zO0gxo8h4xAX317poAVqEVzSxvNPie9tVXtsKrkVYUViE
3igTcAECtPlba+qQtazS8Lj79ZI8CxCedUpOCOwM90ws96E5kUk8G/ynvOtJrBKuSP2zcPVcIXW8
EKtAhfZ5IapyyP2pd0Iqg6MUXsRtZYa2pXnOWF5Ky9ayLl2h30yg32q/4c6eCN7iu1ejOTMQ8g5t
0j2SqFJKhiL1ehWne+22PuAk3nQJKZ+P1LjOFev8+PAV6/2WPl/SfQn/afxoOpHKh0ftTilsXPG+
FCyIcFZHHDxANe42viu6LGOxsYSJhJj7cRr3Bjl+rmql9jdOoV63wgQO+L7U+n2qUixowGvSXsUa
K8BvBBwCwAYeEeaNtCN+3hg7aGzcMiezNSzQzWpY86OhqS1f8p+uF0h+IG4B8XhG7AI3FhzF+Rql
70zKYAEACjhiH4y99W6yPONhocl2jSXJBnZJHhRPFX5lnlZ0fAEvAjMMwnzgN+ruYVukPWuyS3qY
gnk4nlWrt6dAkblkiP5fj+YzXCM+kom/7xOryxuGpHDZD/QIgGvWB1aZ1HqIghAeMdDwO4VACzK6
vboBrHt3PtQL50ppzBriyEvAZ+GmBQGNJFHXg3wxkowoc7ohay7xFUrP06YgnsuyEvaO9sh6Izgz
8GpRXyGDVR5Fl+q/fRzuCksM1ns0rV0z1cJdueD7ZizL9pTQZTQ78gHc/YJppsSG3kNE3Zv94bQb
so6D89BM+CYhfNQY8BH3RL3rm1+ug4URtRHXiLkH8toXDaAc7JsAqjZYJpGXyijAn5ST0hkLEwUi
uwrPoo8vBgm8w9CVEHNJfk+hjE+LwO60WaJL2QKdSrqBGUfPLdnCbYlZikE5SdhOEXfRNIgljrcI
tCf8hLnLnOVfhrgLZNwCcv4SxKs8b//lplO02DI1ml1wliRZ7y7T7NfPMX+eRQuzzcbAEuwbTqsb
LJqTPas51NZxwfTYY649dqEAU8FxzVZs4/mdc9j7t3Rm15iFc48usnb5HxlWsG9XbkuhffVi+lwr
VNlnUy5MDoVrOTFOv9qdoBMBaRwFD4KdjDUraJ8tvTrbGi4ppzK6DFcYUDtsavjOrsRfMwXNUice
hdNoJA60I+2Azye2D4aCeu6WXSp1TnlZ0zcBOJ14dWtljKjuepJY5KYG6KVJHalYVOg9wRXJOyan
7EUxv/MfhyJ0bc7Za/n/gUK1eEUW6LkzBliqg/fWvRH97k1MdgtdE2wTRnMtv+iRdy597WMa4oF3
xUdiZiOwXEdzP6BTsPfB+Vg6L69AI2l4DXmevuKDqdmNVMkkurDGyqnIAbjW3nDfgU1Qf1ka/OKp
Y3aOtDdqkhCTcnN8f5bqFvbgzAWp+UN2Vvugq5FRjKT60wH4VESspgcHicLjedCqsQUGRGDopMQm
whZEwL944YLGPCgF4EHNMfB9kdkIAfmhSZQ+4nNhDeb2kahOLk/esPsM+yZGad0nGwZ82pqgl2tJ
kQz3xen3JFTVSF9BjrBVX0WjeLnb44zjsyCmP6p43iXijXmUzf2GFalpECM7i60NLfDG6VhO0ub9
pf+OHtPRrBJ0kdM6wd/GjOAT2VIom7fhQ0+N7ilbaCk26+YyY3e1Fd3Z+UwuxcukawROdFXUnOmq
jA8gdZdIxhtlHdX8U8xywdW8QqPH7yeLp2wAawB7rrmfUDyu6Ok90eOLc1QwwlBQl9yipm0LnG7l
KTWhih5d4HRnmWV8V62vILRbp//NO4Xrc8Bd5eCqcHOhdBm/c96iZYBsPkDe3nJZznwXOEk7luLm
VJObb4DRCMRb19KHnPrYZ/src0zzOsXOnxRNLwHcfUZx3BPXmIAn5iB1OClRay5NZLxo31dDjnBS
P6HnX79SxOI9A0BKWJdbM+nWd3WqP3X4ds5QjBetaKK/4ITkM72arEjH5uCIdnhw8zQbbgEEcGbV
Cagkq2h//KbpUnzg0bfjU6V0kJ2/Dp7kQHbb7xF+6jdJBhUpM9RUIHWwc96jZkrDywBRK8VqM2tb
RYMxYjJBMzxROZ8wXtyMDFUGAV2/NuIT9HA5JeH8cnwhw/V4wN+YKHM9p0EgGO7q2ta9VMJKRGQa
NyBmAgOGxZrYDQn9oSTpSPY2vrlmPSjyeaeLHvTge+vmrGImsbOPKS6MN14Mfv5yKWLNBb5Gj2aL
THW6YyA6OhpTgXwWjrtsxiCoI9aX9r6YD9OHpUL+l8Mi1w/Ed7Ho8eifyZbcNJSGIOIriR9ueIHj
lzLqY+l0yXXBB2FWCcbXFabP2BrNOSZ3dt2hAn4CHD1M90FlEJ0iaYYaNTytki3IWCsirtNlaR0F
+gUgJQ5YsFG9JH5Pj4PVl5cuWal7IyEjxXvSLw8JWegMZ9SzVkXzJua1Zbom7MbBHhG3ZvDYIrKs
x8IAgldO/2d3T3eMZSDvdz2AkWmrBg/ANnurkBBNNzGJhmdpshGdbeP0J/dYY91zNO1oU9J317FW
fE7DX7avXytTXZs8IjSEaHLMOhgg569jtZNtz1mErimFMD4a8ACRMHGkXrPMVWV0HC+fJ5xbjLfb
/7VMpAux0Efm3X+mzr5NAP9VsmcK9kba4603zJrNhtAP9Gtm/H7TUwPe5J6339IDWHZx/DHNF+U4
obndNNGHGIt0j20yKwPVt16DrOE6JUrfAfFUAY12TrGiZeyb3wHpted94/XzN1Icl7nnoDTVsFpl
aT6UR04COXb8w60XkKZaz59eRCbHW7KBA6/kNAuK/3ra/Qc0XJjgFYIhA3jQhc/92kVx+x4Cv7zp
zxApuTYzpQwzbIqwL7aKxa7tZcGCWOxvzbXL6H8ljdL6PowlcFVrUhtMCQvEYahswCDf/vKf/+B/
lZh18kfXZLuRl4A03fYkIIe1iQjSrNS4njj6mVBNnTlxZCDuLG9MptAXiveTbyC3mHeBilN0cYqz
DxV9yDOJ8H55vBL/YxRgW9cU9S5RpissqiLD5Dd+PM5ra8lfvPVIVsJ7UVo2x1glYrcTg4dC/0t/
GPPrQlVdB9sA/Dvuyr0QKJfXq09WBugz88pQMm1Sg1b+VXNGjMV9Bzc/35eHZmpDSnEL7LEb7Fpl
OlXbuwwZVkkCMS+xBJQ3xRAjQxvGRZ3mIHPMhXzByVzSQ9kBYUydVCR8eDBfJWDYRAxNuGubAdCT
bCQ9jNgeBe37PqOUm4A0BZDGTbz9mX3RzlnyMwW77ahKamNSrdAeD/ChrZYOuGPr0V0mKqPDYT+w
fQKGCGl0Ln11kTGKA8APAwaasrhiocxXwh1hYrCFPs8ZIpydt+gw1JmoVUByt8/11xD17LWschDt
vrUH7ZkniiWgcYxL9DyUIYlr0ZKTvmL8NGT5gmFKzb1gV2uONN1HalmrhanZGayJ/QyzRg4Juet0
qk2T9OHaByqO3NQybUocnRYr0m98Fno6T1xE5jJ5iPbk6kT2tESymsW4+3lS0MFruH5Svai2bn5c
6sCDNCrJ2w1g1y/fBdd28MVrdAICqFOzlpgDQt2n6EAIIstRQvygdOVbNDPrHmwzzfkjJzIo8iZs
v7jCYGXeNxe+TnJiU5Bi6YD37uu4YYyknnDNC4OKREdugTYExJZ7YcWWfE72H1TIGnYTLtkR1/25
J7lo7+aJBJpXLGqAIJpuwqrzSSVOAydKTv7+ltkGOK1uCHB4ARCU3EeN34We3hdeMQ16CFIkj1Yp
O0Fgy18oZD/8X5AiYqEeOC6jnsI48zroTUBz5c4WGEv6pBnk6FhpS2pSYf4HSac4ur9zYOam2/A4
FG94pgXYaRNZOJF8K3XntlvfwEeDccqpL4GHKg1LZ+2G3IGVVggT0TEZ29f0kQQy40W1xfPHKSch
MczWDXXkqBcOlytgPu7IcvyKfeG5TU64oQlobD75KoyxPB2BM8EPNQKmFbrnBrVQFvnuBPvvkMV0
shYxxwEysNl3FRJ9vOHxKj0YaGA86G+j7GsP7mMkMLvZXCc8xq260SEpU1FFoRMI0nPGQy2g2a+9
/FnSJZNpQQHyxaT3xppJcvxRVH+2ieGFXKfnUJS2c2yIE64cw4H6NwiBRQOGTHVBniLCT3uJjv9W
FhVtxv7N/TM/wKoQldrZNx0GVrvRrHlPotpM3qfuvkPA7aKu4kczdF8LMC/JcrGJt2DAOm+xzNsO
Zxtfb7oxdeJvIppgF2cJZw3oBSPgEwUw26JaU4QSjbt0f85AVH4/ZXSLrJhX6hl/Xi9NnrOKvoyU
Jkjph8A+spvU8MafYHhwRewB+p16hUjsJcfZkqGlpStBUfpgvlRJY/qW6NZxKnOuwVu5si391Qt4
g60bgih12ha4fJuOTrr76J0ABBLrPpz9ssdkCX2cttzQOQYSFeuBdrcR+DJaZsNISEn3P+YEAhPD
4hIwmXz0SrSZnNbEAszDjdvOr3xwOc/FD3J1GocEsQTP25Qp4RMkfotgamy/xtHUnaMxBDBrvH2m
OzlPxrzLSDrKbAkTLUB+sfDkpVrimTFHPy6Q5nN1Gtm/m0oNSKwXZ5/vCA+1rVb8S6h3BZTcpw+B
42dX6g7CoF8J0BhmQyUwMwHi5aE0vvkY71UyltI3H87PGINRVsXBRlY/UrWidMHakvXzQKS+R4XG
E11cFej3tPNu4m6zYsPctqYXEBPxlx/r9eXtJ768EKn15Lvsvq9dAydorCgzKuPMN23J+Cie82Xt
HR4bw5TAgUARdEIAf4oNoGMYS14bD3rQnVRSEXoil8Xw/XyhjgRbfhB36NvGhgj3D4+MijP8Kt07
TE/BP/i+gwhOaUV79mfhQbYPVrVCm9m+KeAWG8F4qXqnQ97nTdO5Mympl++w1cr4Tb+/Tx9bAMnd
lBb5Dd+jcG6ulmOuDSBf1nW6uMDUl8zhXV4/kZfKJP84Tivf5y8FqLCTFlIe/0GiKqKCy5lDN5tD
v8E+maIjj49MQzRepELSkCfiEGrkoteVcst2BepJogMwAd1QOrWWcNOiO23aR2z8FqDL197SDYXv
24m9i+rGCpIWiDdgK1nDax0JiY5n609EdjlLIPyza5Q0wxQF9AxpeK2M5jcyfJbtr/yejpz2Rg3n
3ya40jijan8T1FJmyUwvqiXBW2dQyIhFajm4ZN5oVg12yGDhomZN1fUogMJ0cv5XfYeJKhABe5n2
YQaSboKqcEjefScZ+/UfopUzAXZXaoz8b5Pm2GI4iddZtv45jqqfIPRBgXYE/yAHn+FQPzHVp/Df
s4jLKXZviYFX94mhXhNtn2CWiSH9B/rvRY/ZcevuGqbWThdVJtWvE6T4kDcvT98yq0s8l/nFTt0F
opMp3aiD4drY9xgtsVRwmC6jmb1Tdq8+rcZYbqCVZ8QqQmk7RPPNKiip7InJU9nJZnHcfLshHYxh
L+U3SrMtb1tk9XgtgRg8aYS0nyC67oSLfIrDN+dfSbM7yyLsfbTb9aeIjtde21rW5G5qx9ohPKQ4
UX1B/3mT5kKEnRCOH7/9YHYt1adihJh/ETeHys/azIh5tNgYSfy9fqHJqssr7wI251/PJy9hmUfp
aY+VWbYfcDVKMRUgOkFvIKjaQPyLYGOkmBEnASpE9D2kyn6VJsjTkxUBADJ0JuKXjf2PJeh2vLOe
Rc2DCgIwOqqh/IhKlVJKa5MpWYIwo1249ZPDlJEH5Hi2E9TW+mFf5Uv66HP8D6aIvzTYu4SBBe6P
OD6/MxJ+vCnnaliDp9dO5uN4POqDDrVDed0RLasa7oa/g96Ud2Nx1bylbod8NVCI5dad8aFIsyam
JRcPW4DPBr4bJXB1IA7FKovjR1E/fmEltFRcEeMRBGYXea+c8QasZMuFNjHtjQrDPlft6oVfm9gH
4P5/VylqzZ7UFYEr6HH8fRBjUZa7s6ldiVhFo78ebXZoMlD3D0uPEhYd9gNgwQEVQXxPpuLVonux
4X05FIvnVKFPvTH28zHpyM+J7aQHIYs9totVHK7/dFS0m2OhZwdMCtU5yGxwU50zynw09Fbv+L8d
U4Yeq0Vl04RPVXsjPwGm4Z279qIQUygjJydPv267t+LF9/yFwT3ge9ogwDx3wFxt3aSB7rPyckMJ
mcYX8Poevo7RjlBX/t1OTZ9j0UF9UxTSkAdR3su2jJB5AObdKWI235ombVI1Ey/6sq1TuOGPltdp
tbDgiGTOg7TJdfj7MiOrh48FC6yR0VqeN7X36y+xHzHNf4i9x2dnaRTc7r87fkneA5airxVRqo81
ijtHP0S/8l/v+aAJazQyhDWPkVb3n1aKNAntOhRoArBXo8TqGEzEEexoztdtlXvgCZyOeRsN9o2A
CGKHzsTNg6Fi9dVnaF770ajoFijRhf8Dt2JiDNI2aZFwxH04pTOrh70+WdtAtzG37s8ZMvA4IfDc
oN58zX0qW/hGzZiHk99T7FO9kCUlyljKspr3wk/S86R50af/vB0reYZEZQdVooW1AX0JPkHTfQdA
c5LrYx/2ubKmEqQAakIqWeV2+z7jGPjdKEQaVbvDmBxOp8UEcH0Uo+fUFx9GXSnY7c76rZgk94+S
lsdWOCZadEYFATBrOSvTWdXcyoROJa980l8br9p9tMCxEK6qGOb+FBDkwF80ophNjQBA9XK7oho8
s9PtFNLvarZEtlptfgg+bS7/Rpsci9ZBu/F5IRMwDgsvsPTZDpN5djzScwcoRYpDqEz5Tl2zNFaV
c/dYJPemS2T+hjj/GpERZpsjJQkSIZAczREt4tlWugXkp4QijzbpRd22rM46ZzaNiBOVwI2YKg+8
R+6wZ8fA5WDCYOtKYsRfPaPmaEIPQ20+P7uLiKaWDjvPfiMYhYcmHcxcnxQDXyDu4n+nLMtRjXCm
tX82Xz9tdu6DCtxo1uqJu2tP9lf8RyiL0SuMFjTJYZqxKiaoNEJz+chRNKxEuvnOql/wM20fg3mn
TAiFs0fPbpbETSHW+ETmQ+FJCFq8JtiI98a3KPQbUFy1mmV9HV5xqQ3MtfASCM2fQDa/nK1kCgsa
iWWZZ5nsIBJv2+jRWpYUxiN5jYYnJcFVSK2qccRMb4eUeHOTU3DLg6WgwRapvciciaOtZ/S5O8Ep
3VGDcHvlygKlv6gyr6WDbtpG+WPvWVcRatqLy/WnpS6DR/cd5GUWlogCGRxzqe2TGvgUdwfzVAtp
xZ7q2qZFlKQL64rVWvN0zu41bSkyg7JqHB1/QiJnGPZRugAs6sGkgvtBSn2Aq4kuBjq8stu8FCIB
lBBZMTQEvQMwxf3hb4pdax5ZpcTL4QbIbCCuGGIl46UvQY4+hxC3JprsNZawWRR7G8Oc12sywAMg
v+ThyDfqjNHbN2SgxcOV7nZAt8daIoN3PPifHjH+/TfwbjKPysvq46a8uoe4Ge1pJLN5pjUrPZcE
ao89mVOTZpCsa58ssxzvAnGFyRcOnS11OALBhoh9Smq+Sgdvsq4buWJn8vRxyoSTimDxb+RT+TGp
UmEDwq+0T/p4h9Y0fk7dcYY0ncWYX2uOuA5YoLTqSpu61sDk6N+pqO0u6GycOy53DkUUJOddLsEa
8IITLQeOItZljJ9gErBWa5v7Xn+lbyIBkwGvdvO9zOtK9+ml7NL1iIZq2l+wnPm7zBTVTd8VSa7b
ttSOKglc0hBQ3viceX/szsKba2TksTXyPM3tOPw8GQ8MxVLVYoEbBBCSqizbI/FvlL0GtQZ1F+0c
5Y38SF9jilAHb1irwjw8twKzfK52uXfvfAoe14SvND1RO0KpC3As4GPjhltTjHkSgiuXZ6xw9b3j
89G52TFZ/j5NoVSMlOJuhhoQe+HT/or49X3B6auWgkWRXr1uGEX+vFp0aj+VZYNSWYT24TnjDqXB
XQlio6fY4f4Hi21/kjKQTFWr2arNnmh6u5KumauRmx13LQvwHmEbR5f7Lnr5tF5txDWSny/kDQc0
g3O5/RrDWMVkx6Be5dcAOmOs1Z5e6luI1Ag0X++XXfpetfTYpvOdYXqzkY9dQwClBquxPVxGyvX2
yjG17fT7q+dRo70MK0mPh2E4GAlOy7lW+Fe4i5uuKIL2F1r+y8+wtwzN0Q402/BakMwX3a6d01Nt
+CeV2Y4T9k6O3d+D8eqM5Wklem2d7prxBFKyfiB/HCVcO9tP3k2BQcJY2o7bXlVF90mB0yfZy/6D
zfmQ+NALMqSpF126o2+unAeGsVvTn5njTASxzePFzYg3Cetm7MrH8qGR+rFyWD/JG3ktqPHP675b
WonZhxEK+enz86ywd+te7NLEU0c83NRTAB7LfMCtQJepMX6RUYwfAVCbQVM29yjYw23nZMrNkhWH
JmXsSKx5KT9ttI0m/9Ta6qpQT0DbYRTWfaPvBnh33i6JOyjAuRuv6exBWZTs49uBCK5JXT3dUYAO
0Qy89aU3rrblALcwRDhvpTuVx14iorDj6M4Q4wEgoi5bzfUf2TgxvJfSuVzOQdXROpc06R1VPKkf
sqoAjFnvdTmmgvL4FxPQBhObEmQrrmXz4T9kJODyeltQt/8x85Cj5/Psr1d3xSTLDS73j0idHjWj
OWPbyz+VZ/s2XtjuclFwKf4bhrwjKbcbyItqXslg9nYKTkewcG0/9prorf4nIew6TpE05V6zHXKo
gDXa3aw2XnUElmBZX1hqD8VMnfCBx8gW2yBDdLalvdoQqtoHaFzMFLJugRThyk+g9YsA8RmKp64A
R2cqhtEYb/GED3aL15UEQcjm+5WnF54z8G/vQvvTzQ0suLMYYW8dF8fEaoWsE/0/kmK8JR80C59K
BbQ/+kdd8R8faVWrAxOvIBI1hGSOSlPAdZVBtQlC3tF0TD62y89nnB1nLR+XoEWYn5AGyOA6DWUM
kg9HoVvcD1cMg9quF3xd3D8XH+cQhqnvKGZYpnW/qiYEsxQoR0cYKWt2EBOZ483xXR/s9y9jPua4
LAZPTFBGNO9ZlAN8RDwrnR0MnDIDWTDnISp+o3vlRtue2cKhlxozuPBONDVWfSVTrskH/aZNfZ7L
U+k36Or0S2HyUZrS+6cvN744ewHA6tHv8ijofHkHsddO2OljH/bzaj3QRUsuEq7LKBW4tU2VQ+R1
kN27p+sh0TWfN1QGCXEMimBWOugTlJqdBg+ObNipDRxVkcL7evEuMoKHN09j/JaxhBA51AYjIh7k
Bgsct49HlB1xP+9nmWW7jjudblxKKm+wMjxU7GYP+5m4K1J9l8eAMW3cC37kj0+HRsrb83F9swvo
0CvXPX22reIA+anXoPuP/nrdAbgY6UYTQYPCbGnNDxr646zaEKc71BNHtRdQ+hhGhNdf0tXS69Vl
5FBJHAuPbSuq8Wj5FlahXqSGZq0t5Pm8mTHuXENa3bgov1sQgqjaiU4sjiJ19FHMnSL6/0p0eJlD
Y5W3ws7p9qlbWvKedrLnwxGQM+7YK0Ld7wPj2BotQ/iAUbZq2YMgnzcOAf8VWR1+eTrwyfQTiqdi
nQC50CsbqfMX5sCbqiD0iuePuJgh7dDs+ALzgCRS2hrPCBk7ha5nKgV5qK15nQE0to9/ayDAtBfC
S/8CxGDqxaul20zd1Ybx13370Xxy1CEe6x4BK3srwExVtuNkM1LZbmyevY+WFYGx0o7S+8FGMsEv
cq5NonaWqby7aUUNu+/TvRnLwdHlYZqmgsJO24rxIKbMsJPnkraLIaulfHT7IEn2YjHr5KMKXjpp
iCDR2c+BYm3iUafr+0qUMDIithHL5IoMiMrq5En5hE8epT9+Udgex45yFB1Hc4dWwfik3UsJZdpI
mIrmXmAmQXobz3xBQnZd8yzwcseqkiM0jqs0AzdMkE3DrGfElpWn9XwuYpdRhz9rV5YvVFwY/kO9
ZfpMZXhU4P6TkEDQTDesIsWkLfVIon7pX+cjvqbyp2D44LQJQPEOsGziNXI2+AbCVmOSRSuiFwDq
5KtRiC1P5n8MGWv+gif74cCQPEMkZDjNcBPZKg/MtzDirW7U9Pcp2du0E7UcrS5Y2OR5TrlwmgWX
i+L0PdbvQ+96f36kHA7nj0f0C4KdcQ3fh9SXIHc64Rhfqlysiy3L8Z/GDlZjaRpyb3DzB0y/c1c5
9v9LxEEdcDyupeTrzE37bmP9I7nu7D8P8BSTFJXm9xwiOv4dfL8v93LH9jEJidMhxJbj9zB+iaMD
eM50kLbLMkRYJT+hY3WgaSA3VLE32hleb8Dzuydjwm1rW8nUd3xWtDy7H3vTxionYhTHLFoW9qBb
zz/HGyKLJdy5v5LqLASiocshZuvC2xAgHj9fNaHN1gT7hu01P4jKgM+3jVydW3NqUWyIjWXAGTU8
xcuIC2cZMBPSJgonuavWX5R3oQhCuuTZ64IAJX1uW1rw0aodaGMMayILK0RC0PF7qnEQeTno6Rrn
yvOFEM8g95hab1HTBIeBGZySJF+NVqsWpMvKai9coBx8lHrSjOQOD3Q6snEtlLZWwUpRtHBgsQCl
pjDFvn/9Y/O6xv8IMjJPRvJN1XQU6t1VcYl94Q7tHvwOAQTT448GDDBRTyLesn22cXemsrtwGiX1
AKnNlFpnfcbPrmQMK5OIF2EX56cjLE5pg8ZKLWQQq44msuJSlDvxQk7hS73O16Ry91SnUDb+Nakf
Xmk073lJWkwt3NwGZESxbIEb3l/ahU+yg03LdPZYcBJL7HF6yMfr1gGKRB76sWzZen13yuFMded7
JjlQ1yWFqCFhxO1ZgG1yysxKn8gmCSOODPr81yrSBiH773vcVtSWfOzu/wUUPNvkAZVQKxIiY2Rt
dLyND9OJ4ZeWG5tjQURWNmlp9CMoHaGKkiXmwHsXbW+V9BDQR9NMit7J1FFwoXx1BdY+dRtLBj9Q
bt4IrKsZ7O9iZJ0GQxyxn6Xd62T42uKLtdaBCfo9yXy4/qJxn4G4IFtobO7ZX9VStOLOHhT+Rpti
mk6Il/EeFl0jL4R93qj4XT+dED7CocnJFLgHk2PttN3xDaUdLgu6DuG4EovhtXYP5WNebjHO/dP5
JeKgp+9wkUopkHQaGlCUw/s5vrdhoY22U78h3BsS0V3pxRuUFAb+FjKI8oeOHdwORVyXUQ3HEP9q
+++A8bvo3HItdwSGi7v2mhZHIbGlRClqwSA+lNrMsfIT6uEr8CFBwI2ZF+TcT+me/5rKx09gHrYi
hxoaj6hBphnk18A14rUTv0Tuq2wxZGixDadHmewuwb8Q/fyNUBDII/NcnTX2NHAggfnUcKe/h3+0
YbV7lJrhMs2EUvEAaEmDw0yBlLj5DzRCXL+crlGV+nbVJA+U7nIYzHsI8g5a1z35fQ8Fc4+7Nu1N
397IkxD+VHmTSvFfeYZ8cFVUr6yAJCHABKD+Mr2XL3LEE331075z9NLvG+DqPQRweFcWu/80HXbo
rTQwY2WVM29l0tK6XjSwuM0RgNn4aTzd2wL/x95ez2KMzDsAu96qyFIZhFtvarckkIDZKKUnNs8b
pU+ZIoQ3JHj6Kw3u47Rd2WHJ3Vu0aOpPPjN+Zupb9urfIlPJpWWwVf4R+pNv4C21UA6JgyBsSl7K
QxhrAgGGQVzb3G5A3W3qiRaXgzKskS25JQXHNTZvPqJ+AkFRRBcLKZNS4Kh6ZAVR8SVpicFINQeo
qlvpCwD8BIBbFE2fAtmjly3Y/WE9ulOCq9wkt+BZ7uPiwwnu0Eym0qTu6gCrq9nyLmAjNHLll+xS
8sRoRLsfRMDbadVSCpoejatdeAIYeM4f2dEg907Na4jy3kxD0yOlHvAMh7JozWsGq9MwbGJA8hmG
5GdmtKAUXGtgNvHqkpfH3mPEGOLhny3TKjoQb+pdKsNuvXbQoGBP7Fmmt2XH1GqKBWNsLQqUDZ6R
uvUskUX3jxgqF/h+SEhEWXutffVuN8Ko/ttH1ePS5oFKgsOXUncd/OT7gnEWCiOSkjEjEv/wglCK
LHoR3dbjz1/ypTNpDtk+UWB189zI9vKyfYtfHOmhNrlbkpAP5DFkCQE/PCghm5oOROYH8yIwqEjo
8g6CYgactvIxeQkWsrLRrWZh2G9q0LEW5kRwIb+8w8ocKCCsuWH9JI9JgdPSBMyEcAjno79j+CWR
b3CIAP6nXbmZQaY4ozXStJxlL0QC+RsLhVkVSbsx4OSk8hr23fvAxUZEC2IfEQPUjzuNaH4aBuVB
w/WR9PhnvO1Jb8Skyn7b3lgrsz0c3OqbMZkzBLSr1D9uFnf07TDzUCd2fwy1sVNY3oPFPsRC7yWJ
Wx9TGncMSknzfhq5FKeO3q32H9hQau7OM0EMjUcgqxwh622rmNYrZPlvP9GiBPhkRweidi7V67Be
vhgilRHax+dIqQONVeYusCHVEnWCqKU8dhKfQSwxsPBm5R0Uhd//FAfeztFHUdvHlaRh2HBfgoZh
XhfUL5VxXJEMV5dngEPMtCA2FZBGFjlHkmxSxJgJUZBTcm+xd+mYqsRjeGMSqdsgC6mFhLtCXhbd
sZe/Io391/9312gxvzkLGK7038VAhZrGReTpZG94RVS4R/i/TMXuhrQhl6Siz4JCaelR/xYluA6m
6sqqq8B9xPBkJKTH3NvYSXx6JvVg09s0sd+LgT8Ro2U+QlapHlIvVCYCle/nIAF+Il/Kzaf5Wg/S
sZoEZ50htgcT5t0PbU6iI9Y+N0xLhV72xz2BbfzQmSwX/S3HsAa61c6Qmk1feA2I3D+FfqWVF4Sz
ohMfAia4nd/6C0kzmhwFqJs4NusxWWDgWGpvMUVy0y+MakslEfxj4bYE70tdEM/ycCX1hOQTt8J3
086HVTjBpeE2AyuTulIdqy02RH8mMV7LNR/7e1WzHOg7KohE8RH5GO/xZbe9rEPeFEvI0ap0vvB7
7H484BIioApp7IQA8MJU4RYePbzlLrWmKgODWoFdvwgwEMAzJm4c16Cv0/T5Y/fhY7vEes11zQP9
ubj+IaFcr0AFIfDiSSvycKfSF5zoGeU2SKJXLaWG7WlLWHahbz4lZXjpC7Zbk5Lh+1rF2FCHMfvc
t4Sx3m0VaNgo7aPrWl0D12z4ej3lodJYzRBSpCpuYKaEvD95gKj/SRaUZUnFWjRBD+Tw/4Rbikgn
uBmjnh+AF0OfSoQ+lZzdG1RvgWe+hWFNy7l2ppUfVkxpoD6BM0joaXfbytCXijntcIHxvqcLiDRh
DuntVE252Q8DQTz5b7JO0TsMMtVbv4HpbHh4U0mKI98G5uvpVDQkQ02//N7pG06S6PvsRpdYbwcd
fijh1ytyqACJmIp//vRntVvpetE6/Zr1NvFcn0BWA1WxudS9C/SyN1HWTaPu001LWcqaBLyMf9OV
HzR3C3u3TpNcPL1zkqhQphFxb5SEHb9Q9jWiOqIsZO8JpiD6g93ZWtd0EN9XaQZA1Ig2ZTxQLUzv
bFJhIo5lp1sE+L3jOcfdBxJ1uuzv583do6x629NCAzlcpZ4dnak4LSP3xff5ibiJz8S4qx0wUHXC
JhC/+K1Suytu2nSfguE0tI85oDvzeFgbyl4QaAHMJ5RK+81xHXUJ90dsQ8CRxKmszk3NaxlIiqR8
YPZpW/KtHPaUGm6YWZ0tHotYGE3+yRghLJzcXd3Ps+Jq5bzEb61Hs/9JfFuY9fGSsq5BpAvOgnjT
MaUnEqHds8x5cbgmTFAyHeEeVWpcSMZMnRYFxsOrvT4dy9b6uKm1wBgVqkq6yUjn34spNSUDwkGd
9r93uKJfmjNO9AKgMSDd2gCFfSBPkG7NkF8k2LFjqTJR31d99IjS/3wczYJbU5kVklXtpGKSB2aV
h8XkL2eswuSkrD2Sw+IXxjI4GnPw/385LNXj6Aa4+nFJLLaQDJg9JSz20hPkfTyw/3yIxk6N/WWQ
1/HihawKhGOIDITxPP9Amh+k1rFTRQ1HmZfoIIsh0uxNgIDYp1IEwg3Elu7ATJnLqIs11Db/VIPC
c4btvDeb9HEUm2rT/Vgx+HBM+BLLSuDWXBuNR59MXdg5RmmN3v5ifjZ1+VAgmEyd2cb57Uu5/W6j
7l6BpAGuYgNrvKQRUgCyNr/IYuILzt/ZqlA9SkUydc0MrAUfHzn8HIluXnAZ69AvCNLirjE9CaN9
cnKbuoBjcTwveFyH1TqjNtPQ/dJcWZp0asLbp8CQoeoOfI1c+FavKtBYnAXCD4tk0IYiB0dBM1fA
tl0/5Te5f6tchKZA5m2F0nR4BGokl7cRQ/p0qPPF1vKj+ep6BvMA11if7S5OPASTKDYsNxXPlDIM
JBIX1RiIMfZz9pUh7AupZR6nsDTzvxlXBjdzrKq+yO+IfJoGHYyFBFSNEjyMHhybHQuogumgGJfV
/yskz9xtJA/PbCyztvp64LGTMD7bKgX7mZH1bxyIaEnI1Q8Q3sDZaT9kQ3blRHxNMmeJQjVIiHQa
8wzs7ZzcH8jFcOYCPmRVTkAHq34x1nNV6nVL7lmnRY1PiARmMbebOE5C0O7QGacpTDG5wJ5xHDAL
CtWH77SG2YywYFbjDsTu45BelbPg1pF4CtTefvDAB1pwTd73UERMcrEYgkoboigXbUg/lGbrolpW
8y7Xs6JywzGOBh8axNqu5WNGwkQxt3qF43bNNa3yD5jfdWmzJkvq0h5BmFVSU05Ja0/aWEQAj5RI
4EktupHbPcE97xtftiFGPBhbnDZHxsLFs2Cj7mnQb/Qs9jWBAgPmoTGYTMnzgRYSbRbc/9Q+16dZ
BF32rCdkFZfOOWwwnmkloowHIGLlkTF37cuWTY0++qUmxDSPMkN/BVXdMEcukRAHguKWaPE6N0GA
2aq6a0AlMBYjw/qIHtBkgdee2BFXNrteskjlmddNp80hFt+SJFsPQsW2daYkzuCO3mzJsFWz2fEY
cDWb9sIc2iin1RipKactiLckcmsloXDSt+dxzybY+rvzT0Md8bkPwktUj+zgGiE9mGgL6nR480RA
NLrZzGMtbgCVbQqPWgAA/3WBYQbAGYUlvaEIyX2ekwnqfnoXtWbzEUJzhfTNxkqu/coGxLArUf/l
K8+7bRi8fiJstvKmYqeJq1Jd4J/utvPIUVUUnBloIAmGW/mkF9uAxNZnF+BrTYy0VjxbAAvB7/6t
/Ii7LBZvvPqT9CkDQ6+Ozygq/NWV671o7JtfYLHxqamgdx650qx8kE6sS+zoROqLfLL1JTiVngvx
dzcxfRGYsuVYQSswigybSnfnSJvgQscwTGY1ntDqg0cUgB16c4SfIKXP96YTJyxQM4vIyh1q+U7s
UbSmA9aqsEqUUlB7mVus0OcDbTwWv1lHMRK4XdTZ4SvGODpjRMT0xSiL+pfZBsoenUF9b18mJuD0
eZBOyKs53D7VtnPY6hEBopPBBKKvOHWGLklqEBpneoU5dRIIB3K2WcHoNEW5wOEa4QmWLt6dSlWW
O+JV4fkS4l0pVabo5MAt3y1zecWvANcnPWgNw07csjots3SAYltsUQFstX82uLrkMPou1qDQAVq6
b2pD2YvXw/P0KWKWCOpFdKvSZ3vtQzIIGdctC78Z8RazUl0Dj6Ej5lJRPIpzacnmZlnTOs7druVe
IC5/qkvrbDdyghpeCpGfiWEwcvzFlklQCxiCe4VREj4LzfJpdHBBEHt5ijiK1Z7Nj3RTzf6F9MuC
arbvyh4aQAVZdG7Oq7h4gDmw+0cmm/IlgnikngyH71aFC7XqkXftaB9ONxPidFoNu0rpBIO/ijU8
lRe6EiScUkeqVXfNPV8as6GcX52UV0tMGrCNjYExg7QVKXJcj+xok73XlTroE9VmMOR/idBgFArC
PoyB9i3R5Q9sTtjs6c1pu6+DxSiTo81E8JMzl66gcfiiA7UbyZ0Hz9Yi0rLX0BP3LTOyLT2Hfl56
FKxT0SHujl60dXhvcOK8BHf+TS2ur2RxTqCx12nzwshHriupAzM2qKmBgLQ9S1Vuq7ZytdEmtLcd
NWG45zoV23ikqbbQ44jGYAlxSVyaEyY4wB8gqyydsqldUGyN4ZoOai9gI1Ch3elE2EAvJtzPprc2
tSSyy84nQrxC7iZjAPtIbJuehpGT2E0Ye9pGVT6z8Q0AmHKr1ob9vQ2PIYGoon5smuRjOWTqltDi
Y7eRasDHbCMGgUcUv6Sqmk2od+T8LJd42ku3k2MnX6WU68vzNtJm12x9ab9Jst7gZMYjygypjk6n
pIJ/V/WE+19Dc46NSYk7hMZ3itVfDnw43D+mrNszDJJDj1eKqAfxvu4TEJfQTcxSMVKvsuczd9Wa
+Spvae9l5U5+a38/zqxzrGn4FmQFK0mSW2xRJmAsqo9p2lngS177SU5RH5kPAsNy44/0a8iSw+t+
9Tdjo5VXCweJIEsi0sc9sSGOsShMexthdaQidwqZ4s4OfiekdN8Qi0umSsSNmU1leTlu2GSFXTLT
57zPtppqP7KJX4mEPVx1vMHgq1jYcL/BjSdtPBoycA/NVvHuGskO/FwXQFsdLS2LFjBdswn6BCJl
6YvGNF8m8BWkqYQkiyd4JKBsjIPMXAB469ShUT216gjJSKff/PfQ8JwMimezYu1KSyKfcPD1uKd5
l6HitRBT8t+DexC9IGT2NsO44kF8PVf+HjP1jWq1MLpVg9Lnfji0RPhuM64Sf3+KyBKvWcJkE5rH
Qb3fOkmO9+nCbUKmAadAZc60smAtyhPSmz9uGv3xMKmF7HPlD24B7C9+UTTBD5jnI9y2ObVj1TL6
tHxTmeXBdWu+UCDagqYzJmnfmK8bm4vRhsoSjWID0wBddD6l3OYL278O1RviN7jYtWFI2yNkk/XY
ZGlYbSRhxNhvenODtr4pkd6zHar7NpA7BQ3bdULXju38P3dK62qsJdLUyIa/oOFVsUtA9qU9024N
purinLG1UjMz8NqazyHh516pNyFSfqagsUPXx0p0bcowast48FLksRZ4mQ7uCR0Kmg+MQxNeA2ov
pFYOyaIDmKQAqysU6vIb0DnoJf0rdWzThy3joDtf3lQqVY3emMoBlT9WUCayx2cqXAI8UPXebcGh
H6ZSXL7/XUM/ufBxjai/SM37Z+w/Q+uw6vgbL+HTdIFfzyswC2GdMdHQ1HAldwyBcxkk18Ir3hMM
FRamf3Qe7aRu1Z+pKGIVEkln53H9qx0JeBgwoiH+D8abmeuMEu9EX4ozGDbkv52bEy7XmeRmZDlG
ZRgbSSllEw1AXgw/AfKZBYWv9xqWIKFVaq67kzalDhsHqEHAMfxkgSpnWH5i9xJRDRGQLP/v2uHW
7pyMNvGx9xl8MkI83SIC7go8ZDCC9qmLQ/PfGO8G7FsYBCoHyb5UxQMI2crsDOOoZZYLii0EQo7j
onPQSWZxVJquGXrrf3vzkBY6tJDQ9NOifFmrd0DYgU31h9l3RHftDF0AIMEWWAFAhhzh0+9NXH5b
WXwIF4tarIJja59nVWmtW7HqnqzlvjU8eSLDHVh4TKfFUHUQQrfH6zvcJBopaCWR/QhJU412oOkS
Umsiy595LIkxguaWtH9nq5PAI7MnuS2/rZoTrHvuyXs9+WKdAQTDfg5S7egPBKGA7oF7ZjAXfVcv
EJfvvMB4A9pQBSNUweigge22tIMuHjIaFT5txQBUHhqvrxLP6foQOcH9K0pyxHCYhCgF6YNNl6TE
+I2q/E5DDiT+qy/ZdpNFmcLhe6SqGBkRVDsGA5gbV6OUSa3wFrt6qWX/A0SpxU8qdAEpjsS0Dspa
iMFVx5QIzLbj+f1nQON1mLLh7oVqEyKm78/NT6ghK+IottUhya0MvmsIioHaahHvRomXvKGRgo90
oXB1NEGA245wzopiSw38hJ+PxRBUEqPWf1vbubYFUc2eBk1Dv5/dVrn+PECuuWpO8Ks8u4vdH6xQ
2lsYAQjHImQOMS3Gs3rY4NVbYYHHM/8VadUKl8iHccG0U+EYowEkGeb7RTAAXbdrIU335Emg7O6e
gsl0VaizRBOwnGeUbhXSeiNqI2Yoi+uG/E5RSqMA0uy3MN9rRqz5tM4gz7qUbf5D8yD1vD3npDPK
uVGwn9fixqUhl1iDONMWbkLUaTTJIiHIM5lj5TS4CcTv5ydaYKK/mdJVAWy9FgbqCxVAS/WT6V9p
RjHgh5J9gNCFFKgWzo2ZZqFU3RQYwJ2BvH9SwOwFFVbg3Lo25phYcVoZB8K7ck3JToD3DxqobeFs
1QoH+GIQg1rBN+a1p28ilENj6YqGarroWQw+Ae16q4unXR04/pvIGC3gHQ8d2zFjgwSpjk8prVqG
43igBvZAS94PHJnXNfHfTCQEYQD5MHvxFO7zus2cjhFBvozhGgk3ORs3IqNksey69jNFuL9unpZi
NKlVd1t/yaGwef1+HSm/F2af7Ye4FTjXlL1OvI6EOn6In7j/3gLra+IUPrbqUDCU95aTXEFG60In
TANc/RB6Da+Lg6de1/yzxaBQpZktHgr/vhKIbR22UUdfymdPs3jFVWbWbh5Cpx/HVyUZnjEa1iOH
lskV9AgiJNNVYTRnK3vWYEjkWXvRGoILdtK2/i+A9t9XVzsb0CeOoGRb59kFHC6ZVZYKjdY/m0Np
u86N+tM4RrNVM+qRkWiXkVbssNGXPbnAJi4yZSzjLlrxJLQ5kcIMdIMr3zX7YRZrGym1pFrCmBDR
J0wgO/6DO2il2+hu1Er8TTbuszfceP8UcbOUSIg7Dq1sLyouIqOc8fEr+RHDcs4ZzPqJqtL/LDTh
RGvWmDRCsUJlk/oCaiLr+YeiJjxQHkPRGRiMtoLDFifYpM1ES0fCsOsc8aONSQx6uTO2mH8q/mjM
o4xs2JQk8rI8ipYYhkmiqtr4rFxDaw0yZano+AG34GSM1MTNbxzFiu4UmE9xUbmBgQZKDJ/wW+h9
KZz/IwWmZgf6Y6GHYPHFBLBomUgjZDxg9crEJtWOJjbhOIU0GvM48u6BQwXagf2AE+hfWy6Y0G90
kqiuPCmks3fEpdHCjEipuVK/gWZZnCAay5VgdfRnfNyxop0K5XWj8NCILUbtzx1kVqtRxEMhlPWV
Axgs2xPOVKtAyyxcEsDEJ4VVZJD6IAr2V9MUasGe7vtKJ1S3AMxdPpgvym4Bwh5UKT/rMMfPJ6M9
AVzEiMGQZ44qDIWwuHXJRkGYMSPIuolAboS9/UbwfoxYEntlqvIUroAf3X+Cqcu8vqcy6l8v4fpB
Wx4pUoJGW6L649sQ3Fy8ZZ5nTeeRakcvOboPlvhfOMcHpPLpPcBNVHl5q9A7rYLTtcaYH3H5e1kC
fdhZA6NzH8KZU3btts+ctWnWI1rLB0OopWIcRdZqeLntSbDLtHckZglAT0/wk6N+IhMboioWPCJC
PG76VrAMXAd8Lr5y4+mQePtS65r3NOR4cITnNGJuQYk4NO9X5tosomEbGj/dcujeV8WM3StIcjDJ
15U7AbZuJ21oUKJc0OUx2kR8O4C/EzaZiQK+Q9UOfomOh4VVj2cRtG+CRybToz6DXQi4VVniuDQX
2OcSZ9EaOvNBE+ITJ1pWqJvYqnsL5tekLn6GX60547vJ4xc8npNLXXJpDXqltVVkFNLd5Y7aLd/H
/QsAjhPs95LkSopzjx0YjnbQISGvVIMGR/HIwtkM0/xcWqpNEiNYOvQY10R9q/txUHhH7SPAbw7f
VCxjYv8o2O0A53xwjYo6tJxfaQhZBFnffpIlQfZsOkYfwBL1+v7r0jFOKE8FAJ6keMTho6LbwTXJ
yK79IhCeyhuH/FCFKwlKGL0EIGqXUBDXwbBeQf6deQ5fdFO6iKedT4oDCQDUDsoYzveTEJy15N8w
d8ZxoTP51a8XDLaCl8BNcNGFyZJA5+QWrxUswCUAJd4Nm5W960eHJg0kzc1alUdEYZEktRVU+8Ra
M3u9XAa4goDGKcKv2bqTNQsR/hIiBnVNuihux9OAx4xQQB/Ls1fBkH6KDvYaN7xxaApgQxUY8vhT
QCbUwPI9fhLdClOqCWg5Qnx+4rG+k/ciD98lXSY9KftWWwBxCIuP60MKBcD/DxSq1+kJtH/wE2qV
+/Hu1oj/s5/FsVB7eOncn6KMuHhefQQ8i5Wm+UNyTX90cb8JGJkgxM7MM8LCxdOJEY+T2X9YcHkr
1dmENM8BUKxvzpQOwybPBX2F8LxVgUiyZRZ1OgKWeZdq9zOyTPrfD4Pv/Q/krOuGSKJemSb0pgHp
xbXPfmrZn93i6kb/7RUJi03r1rGLnA6ieT93ixxq8B4VA2yos7UqEqJXvWEteeUocJ23eZNOb3vQ
8M3+zqtVeo0D9oVo/xWAN21wdABHNrlP5jbN/aFDuSiy19EwMaj8SU9QL90zACBQZl693HoQ+Ir5
iy5hjbWMxbsAsF3aAYCaqvfKyS6pV505YHeQLVcZ/f1HT952LMhWIif2JpRhPKH8ujj6VJZEKIVT
1Ld+39EomEjDmODoLkxhIu0a5+Ul7Uld97t7KkjqLlnRqzQpoyl7s30Xjhidn5jwKD8O7lQhAI4r
HrtnXcfjvQQlXPv8q1KiuDYAegY4zF/20HL0Eg0bGb/RV02V70Jp8ZLPqOdF0rDR7RqDMBOthZoG
IZ5o742lAEV1xZAn6Rx/ppD3msEJe8uQBIa9c/TF8chx+q2Ordv1TB5HvkH5D75BpVMMbvxE/vtb
pfX7YY5XfwvXZ/I2/bA0H5DDQvdmZlhvpg3os5PJOPUbr1x11hYB6OCixXqouQeV+BNyGfoF47o+
sOayK5y/5YaS7cjAB2hyc8BsIJyX576qSWyAz01EjlzsUb2RlmYesQMhpIS/+9YtpyggyvyI1cp8
+c/Q2jdVu07W+pNidr0IxbR37oq7nnS2VpmGwp5o+8gWeZpN6I+mjuXnfOOGv5KUed89NWk1ExSf
zTT9sHjPLAvQ4HxkARjgM7qrbcvrX1WfPCkwDyalA4/FB4rTMDamQFLK3z6S9fVUY7oKJdtaEG5W
dga9Uqwv4gTVdYP4OacybJn6sklgQJgB6/vWOPlVI+dxacuSJ9DVKnUw6U2QmXMgHU2XhgN/9ujV
wqgNGCniUYuAzB1UzWaMcjI2PsKhYeLehGkiOklji+VMGqOMLD/jUb9g7o7Jgb2vMSVg07SGkMWf
GF1vu9eZ6VnSQlcQ4vSGBBfjX7osdw7GQulBs6Og6Kf/AouOlDExNUbpY/mNlHXu6o+LYAxV0Psw
GvWC7uNCkcdNdRqtLiQdFsKvXP7k6TMBLPLB5KENZZ2lGS8e/U+apfdA6BNUK5sRmR2QHMdkK/7i
W+snTb355BKcIJcuVUPo6tJMtBkzKAZQQpWHQQY4R0RmkS6VWZ1kNbh4CKLC42bFY92T4WqE3ZCu
3OUR3QhxuTr1b0DfDdqysugrL/gaYB8n/A2lyR+9rQ6fFjKghMRos22pS9KhtTylndHvIbC/oefD
qIz7OrPZ3u5MKAYjZxaQOLEB7Ods/erii+CJTf0MfdFF6Z7EUKO0zP1nrFPNsj0WHE7cK41qQ7k4
43QI3ULzfL10YLF3YnDfry499+XA+uiEKzGd2gBfPBajLHJreJZcxDC2otkIYCYD0v2wG+vSxYB0
VDtmXzDpRv11rACm8UjN+esMtDvwlCWMMlVwhwZcYnxF9QVJ2e7783lVwmybDYEnSaQrNWskonDr
aXUTHzE3JdAUFfZdqkaZYmMvH3N5BFjaa8iC6psrsfazp2wHxT4bgDbq8YxdhfBj0GnTHxy3mKQv
iCgG/hMdcG22co+mYyI1AY+0F1LHbBJ7KWiOx1SxwcDvOJtMigkXGruDcr6s69VB7fIRrbVkb03a
/3nCAs+hOpwY/etlMvul9XAadqpdXYIC4kxB5cf4mOHKIgehJqb64ouuSd4IDSitPISdmTkyNvuD
lrCJUgTj14fKdibUVtru8i7OJK/LGMqhzWcOAYLxS7ktGzSrPSQS+oLjeu/n/lrd0hYG/+8M0Dzn
Eg7rwiZmdUjLDtcKHYIiwyViEGLxEqTQYW1xK0/OVh2148E1Ud1soAgPAMMRIaR76GCf48AHwvyI
5HUERw7SoJ1RHNP5J6wk1Dc+atZUS5xihJeqWHQrtnIGKVlR3JzKSK02beD8ag+xig1ceEtsZ3GQ
P7Nd8K4rN7AHiaApm5OPDvmYH4miYAuqCVps+52HfFSXOapOUbmoR7p4cYQ4WKt4QNHESxLOfP6D
R8wTEkRmmAOOOqTuEj0Lkz1IPv9nE1mRd3hsoFCyc17JSXc+mY6g3h/xXzkj8zhBVFaNmojR8pLO
ARXsNONhp0rgB+Io+ksfDxF+YNFs8w8PRPHgD9dwpEnTUQOVNmrKQptLEM59YAhtZFj6MRWcT7aR
xj7nefoSfzYZL/ctNOIm3Qg5RflVnTNpYGz7BWW0J45foIisKe/6pKQ10tYKOuCWPY5S0Klj0UzT
/X6i22Re89Q78JsPjoOEK5Um+sXXjg2Sz0Hr4Bm3/pIzHeQP5auwrEOKS+UtNAPuIyqcIwYfmmPh
jA1vbGg1UQq3v2BaT6qCxOwFXapi1s8CsI3oqaPlcOlu1DpKB+9HjDcm9IMmIiWh1S3b89wE3gpg
E+OULEn1AJKwkCalH2Mz+9QNeCy+gJaG+spLnBFz2+hAPezEUG4m+qaBiZLiCuEwcjmKT6Dg34TF
iyaz1a4aOdR6L6Vho9kQme6/sRv6tuSxvgp27JWGsYJQ38Ikw9g2rDdyOrKQNycbrv5GwA5MHzZG
erE/M+MPuk8y3PcTVgQP4XrE7Wf5WDBcs3QrPqi0ddKfM7v92PyM6/excSkE/P4tBmuV05ox+/zd
dPvwaS9MxiqMBrk65ZnQ8dsPmM2S+VsS3h5OTLFzM1LCo6anYU9QSKvhxDTz89Ga7koDJfQnVMTQ
6lpU5puEW0GudmlOVVWjEo7eXuhqO80aANMuL7t+8TQhUhnA7If8oI5bxAz0RgmNJMVPyXrgVA/9
BsnyVvf+d9350vXYtFeepGAuURjklD3RmpD26/8Vfelpo03lXmCoXS3cyyoeXC10IRuEC0rTVU9w
8sIVxzy5p2lHwNQLQYq/yI5JVF5Q8wJ8xlyfcqpx5DuJpX4dhJBNymvfQJwMpgCybMsp0osUnZPI
v4mXECFebo35jO+uZ574gKvnVaonKimVaxLhoWyzo/PZ9Za5gP6k8euya+wgk9Y9/y0Q/lONvTQj
fz9x5mcCSFZ8kfKw7U2mx4or1exB9IL+uJfiSVC/COigWUuNpvLuRw/ip83vGycg0dq9yJ3Tf+Xm
c+ZwnFhGG9kt7S/wmivIUToQ6FeTpw2M1VGCM9Xvmme24viy0nZMHPCn3PXuZPhmnYfTKHKXs+GY
gTGsmN07PTgAgqjx11qW8bNNlv2+Hp078eGgRryYIoEYNd5uAeifyx9sgscIkYlFDsd7nfkjPO12
Pe+rsCHTQ4ds5sW7mQs83Cfmu0XtI4unYUiv0eY0UlYb6O34HLuVi/705V/efJnYyAIwCRj/S2Lv
8rviWbW8K1oZ8++dcVeemlTAfMJ8LDbswPuBuxIqfwKdo1qNZ0k3ZNxuS1c8tlxGfoT52GiJDKZq
ihT8V1AJvQcGA3xsyBDvs53IbcRJX5eJcPVsaMyC/vwV6vZUFAUFe2lU/Ifa185kyP3yKZIs0Dtb
FzdJNPCWir639pzZZIZ00tQOi0SIjdKX+IYWoTp6TZEbCL/Pc9tgRQMaiOMj0RQKnXk/xPwuv1CT
v82aMG29c2nqjeq6WMjv6V1Geyl2GxfpXIMmwP0ytQgfSTzK5J/h/WPPnwQaYrEVT8xwHBSlWIEH
ra5FU6OrOLZH6Hd2vINkB5soxGC4ezU/DmpZVF9l1YAK9eL4LOpeVc9QMbi2Qxd8lOXyo1S9P/qj
+vWirIaleuZgc74t1pJ1+hP+yOgH+Uf47BALdclDt2z1uVJ7Ka3/1VQ+2xV6Yj4TCrnIaGkSqG9/
RikQi3EgS2SaShPC1USt+qvYosJoweFLMI4gCkcetaSU5+OwfS0+/iVN1ojaf89jOimFzU5zeSmb
LQbHn87Pr9OSurePrhkrx6nMeh0CUxYP/CXTEwdya5xOLszDNCdGsB1njpoAIcSE+mxXKkpemHtq
2Nytm08+70fZLgItf2uwSLuJsIAhPy/g7eSNapPrPi9KVAWBZdapEVNHnQghRxL7g6svgYmHAA8v
Gu0G7vlyv4uFQD8FDDzzs6xXmqcfs6/vzCvmMdh0nn4a6uWS8iIi7d+OxQ3eTIBKR8xqE5l3+BXl
RI8O5ZhFX7juTbDFClmxUnuePPO7egDHzWkmZEQ8/z1Z6fkSWxAaAUNELBkRFPKD2+XzT2lt53zX
0jxWau/yo1OG9h5UwkGkeRP6ikZ5Qcs1UDppCR/ds39cPJXrYIzygKcjy8ZkzJt1bxfg/OsR4VEW
SX91QFIKJy5JZGhcwRG7fZRVMeaF1HVrNghNu85U4tIHy+/RU+zkAlr3f3J9DFAvRND8oM9zy1iJ
jnwUMJ4NwSx4NAgGrJuBU8eFQu2QzRSg/Mozy4nLmMYZoxR6jelAftEqCZj7RFlL8sJmyrhwr/uF
0ZjXsjzGQ+T+PQrbnIsnoZhvGssANz2gSUZNgLy08oEMuQdhtqD6t4g71LtGT5q6l8QSK8oY9NXM
mQMQrb5jKZW8SVvIzOC6bN3NaBQWnLTi54KKiGP3sMG90R6Xz81EaV2rtCaAHHy1872/2eKaCLdM
6aQNgPf/hmQ1+RaEj7I6scIU6SD5k7I1wmmWgms9rRg7PY6UVXaZYENzho9rJ3BXvghPGa/Kjzun
nXzF40flroYcMeWpjQNN3ZtHuqR80xRtknWJdSdc3vLP/i/ieT8TiewsUEP7jA5TGwqhaQYIhSSF
KdfQR10na0sAc7yvTrZuW/mvz1JF7Om7blVPnyPmABvCz/KqET6sJGgIRnU8UyroGAGZ4/sCKjot
XJV6nU/i6zKQJRT6CcT9rGu2jifF1ekg6tMbGQqqhgbQ1yJtOhdxql/8Brb8b3KWItbE/8nZYUhC
4VUaOuMzaWYDYnD35WDSzl6V+mWT2U1dFgI3YVdJZhrjC+zieo3DqdgVr8VFOwFAVSCCc0pML4AF
Ub+MnQmL6bhAd6JIG2QJ7Cgo6/ML74EClSguXtC363MQyeWNGgi8u9jQ4ksdIBo6uc2APEBmboKn
tpUoKJnCnzKvF5AGk5PHhPxBiLQCPOVDnISvue9Y7C9vcUKR8oWFr8ZjhOeGQ7Zd2/TLn01hpWFp
HiCUsxAmSQ/YBO0tMvcuSPFqh/umTVVdwOfPftRGfGwGKvLavT2zyyFYYCDhs7nb2Ol+CRUl/2mx
iS2Bm+UaqyA1Y5Y0wFyo2itV228UEI49e/AQ9STHcBoqYffJ6FHtLSkuXFC4bBaCJzL65/eyDqvZ
6jFSEvN9TyZuT9SLDA5DFCiyh4cONzX6SY7v3M63WHyQTuZLKrya6r+hDKfZPCEz7Gi9insmAmi3
m7aVq9yTvpg1Qrjx1L4xQSAHgTTrSzImE74d8WYp9oV15ts7w0h4wT5iTZ80qwKu9Dbq/I84iBvJ
ERSxW3J4Z2O1/WHYX07dLDPKkh//EL0vJnUWJzfeJ9LdvnbR9XUTQb80GvtlhPUJtZJfZQ44CF0t
HwFzls8ZPrfHt0naAuiOr1/BsAfu7LbxtXQBGoF18DyuK+u4rZixqm3PcIimqxbgIiQwJQe3Hh6v
IlGhvQvKKPdqeRGEOMG6F7B63bLiJKrBn5oiQOHPep6Vj2GnYd0BnvK1xrQAiPBI8az8jviyU+7f
ASZ1VYtsFRtcy1Zg6w7UDOe9WgFxSJztM9gMo0gnA6spKho0ZeNRMnMP2sb9nJN3TB/H4YCD9LAo
PaRjx3uLYrAq77mz9iiM9CQmqNUyoNb/rBzOckZtl27DGeqjKbyJV1AvkvjtCap/3CcX6X2HnRLe
2jsZ9fR0U2Yz+vNUV+niG5q7q3aU599sDYFL2D/+QrPmSZl5YkkrJeLYqK94gX29C26fcLMckWjB
Ur1NbYVAMgJtZg8RiEVZ0KylnQn8e5lck+vUgwOsjOYffu7IfhIMANahYawBdqJDQRH5PhANcA9I
am2279wsByZKXKFSs3G5Kj2WcKiVnkMKXAYu/0ip1EQz2Ln6OdRbNGAapmIbveYen2eWIKPDIyOY
bLzOksam+3BUIdoLQvZAZJTBiZBoxU75sjSKAfnF2CgGzQbs7T8QP6SVmt/WsTT/aqIt8JR+iGVC
UQevyOSlSFBu8nWrNOdpppO/3XuvPQ9U+l2pbV6hAsNMykf2OgmyszE3bOqedX46WFlhrA6vqte7
TTuib/qFjLNN4DHuLZc/SBnT1LuL+XpDK4VBtnfH7PA7LNisMW8Rha8AxnpXJ4IRGDOzPaCdbdXc
jppy+I/TMEOtiA72j9rFoummI1pJmUN3xTO9Cy1XM0YEQG1pSBcJ9SMX+cfo3Dbxz96zIW/FsZ9j
kkYpeoLP6hpXG4H4c1cqtGhHGuf+wGESxhykkL54AFXs/s6zjwdIlyFcZX7WIsmd1gmk6S+szgQ0
x6zeExCogDL+aCmrkI92WTvKz6SJ6gVh4BGA+MJtyMjCItt1yFsTIP+0spj01nAM9Jq/bQi/2rbx
5dOI+DZZHcOPnI4Wg4wI6D0Tj97GlNHQAdRxOk9O8rnFPWLR7HqqNI50+cySzZbHgXWQ9vQr3AWE
k5lp4sxnlHkR/tJncUrrD2Pa0GcUQhrgns4ZQga0CwUagqceKC8dYCuNzK+LGOD29F1cLzMPMbId
6e6zxMGeIZ58DfKM58FQNvtu/ThL0EuDp3FqZgadV7dh4KK6SMwyeBrEnfAH9YGrn5P+ihft+kMQ
B1RDU3rSOvK4xcI7L0aDss7py0MdQwXwsI9gGJlEFvAQkC5E0yuHOR4qx5Y1bmmzk91leTEli5wg
PtetBKzoVXQw78jj8+H9KKTBXHnu2vH78r6cNKmMCkE1UlCUg7LyJrztsaCX1jRtXLC5JkVdsVg8
a/5PzNsgejp7LUvsCqdhIb3XBTTUqZ60yRKOM/ZwR762ZBrEPiR6ur+9CRoKZm2G+H7uu58p/d2F
ZNdKFYV2oUXqySipthYzTuiqH2iZJyjfOnhXsc6jajsqj4SkPd4hztC8lH7POjh2kWVKrKc24d4A
rA6GsO8xAYdsejFJxwY79ufhCP8GZXV8pvGIjgCd4UAhDfFol3WJrQ42BXU5/czLymGUM4qG0D9+
TZDTWXhaXDQWfzi/z3rd0nlBqybhEtNGuqmZFWEovcGU9PVmhM+kCAojus4grtq1nsVSsJ2aRWPR
+7MV72VuEYbV57gE3AsK6vtn2z+jh7BvSMincerdyelwGUw1wEUhJoY4z71HjsmWMMtn1DTJyuSQ
fGCWHSzMxvRDL50WpH2aiDOr21HMB6uvrdFlOd/dzXMvgXtio5X9MP+DshmIJpU1NBY6CIatP8Jv
JE89dEiMO+YG+wOucmNSeHdTH5bkQMcjGzsIOVqHkCS0jNdPyUFpcsq6wyXlrUd24tTUVJf4+IG0
G+6M5IbHknhLD63TuzAvAnE47lq9bS1ae0DGC9qZa+Iyds0CQ39mpULwpCX4cHz7OAPm+0mB9f8L
iN/HH7iCth7Hjy31dXlcUyfNLuCGR6sgwJ3JmcSuBCuExBZzEKHSVeyZO7kKDHGpCK5Mdw8uam2p
qLrjBRjFlS2Cu8jtQjkQPBm79IUq8Ds4kvR+MifsZ0qOPGdIZLUAVHl3Y6dTgufTbuhW628INkfO
2BCGcONwLJjzsEhfwI1cw7G4VeFGA4bCjDATMOgOi2AJyVdPMpVoB0TRqlaQP33XGznqrKDQuMWD
lA14CEKeDez4PuN5zf3S68mc4LsFIuCNud6hqt2pCmnH50kZPGEntGKVy0fuHbo0LXzqfO6sEL1g
7sGebUQqpw12gJrKrEcTxvfAkOwz8lM8/3aRXU2OR37fs3YffreghsvNn4HdtOJ+PJ/vopDW+SAm
CxvdqJEquqRNNlSNGEfgIx4/iTQC1gDdqMXGwzPrd7XAlR8rfjpNKa78/R87fzbl61Llng/aSpa6
n9czPhY4+A9EuKL+bQT+JI4HP0x3wAF+1crJGpVqtfxxXaO5879GA+gJ29jO6hFCZwBJs4QUPo6C
pxpyjKX7rlETDrEZbtTE7GV2yOmAMqsiK9xSf1YuTSau4NFqINLQiIc6/mN1YNceUTXm6FtIlzap
Uh2OW42e3S7wcTUqYQLYNTUoMiUXnsVi519XolENv7jwpxbRxQE04fjTtA8PZaTHZe1Sl/3bhoIW
GUIHSG4io4Pno9DE8m+T26HCIH5fsJdqPkY19VHfEVbT1NvLtdTSWb/bylO3xsqzyuUFufvE6gNo
h9xkhVYbYE0Abxm2+SozdGmXkPezM7aqtlWEKkS0pJBGr9HhTdOQkQLpS+0mIW6Ns9/adzRxMfKo
tINhJnHv2sT6cJSS0CL/WkCuxsmKpnFiJFDTm2Iv+Y7JoY467gpiJ8hOIIxDkb7BwhQUD8G2Jfe5
FtxDwllpAsQkDJQwrgEauuCqaXOQgCbmo41bE0m5Lhz+dA37ij+ZBw+LRwjHs67yrUNNV6gbOQO2
DPR+pL/tPDu+WqUz/8SLeXQCloux28L+2y0PMKWBe4qMSVrFNPaPXikVhCggtm56KiRB358b69l9
jeNfIg3LIHgiNdB7yTT/SP/ljZkJMkH1O4zH1sk2JsyZvkyQyJVjjnFnZ20WVAB0WxQZJKJrzvU3
MD2mBjAx9Hro1yGqhxYTNMVpgE2WUbRqqen8OEOzOW2xbKoT0XE1KjvEOgs/0L+MkICIWr79uwBK
GG3rvvcxVGXAsWo1CeshjRqd63FeMzZrear5aF/yMeYeNGWAkAyALujlU9f5x/SNy4Dys5PCsrRL
Yahd9Zx4sUZj1ilr7e0rQuJm2CAaJjrkjQW9ghL5IEmVFJTS+KDPDW5HnFsXeQSj1oSfr3JWnjMI
9f3mEiGi3PifhfmvumPizqPt26/FWx8ftKQ3rw//A9SM5Y2lckfT00NUj85VAVzgRp1/DOIb5qjT
Ss7+mbAOSfTIfJpW8ol4UMKG26v74au0Eessz1Lv2U07E7VsPy5cJkldSsr3P9Av8GV5AlpjA8pB
2XKmxk+8Mr65NCWfKiAWLnmWLLr7BQZj3D05w/jeADPWPlQbvrzx5uztS8PKUXFd2O/kKfUn+QVJ
8K0RkP1QyhLEOAXiQwRwSwvu0W9lWLbw6y20pOvbQWuXFXQzXOSwLrSecdj8Y+vLACHorMfrDgoS
LgAt2NZsiZ7wPzBls2f5Vic1Rqs0qXzejc5nQgqvwTZva1BzH8aW8D2Z1/396CDuYo8hoiO6qPrs
ylfjn+SywC3dY7T0Akqnc6uV8wqRKWguHrnwzdCo9/aKnRIa8ZKzIhYmTLIy/KME3cLbme8M3gnj
mtJARHMmsVJfhNin0xg6GAJfRluCdHqWigd5+6aAb8PxJ/wskHOeHv0uivGGCqTWDf4nSxPn/RUy
OMX9j+aXcK9CPhtsoNzp7KYKN6kO6ORA9FpDgimS5/y9kwD3ZdB1JDVQOCtKOakmbNcl4rZV0zSB
Q/i45MD+nziULSHNQhJaa92gGiZ9rznYe9zQQ8e9GgHLDf8arbNF2BmypsFIVr/GBiFHfbxinqbs
KbjOv5H1lnF6P7X7NhkkFnT8I5zXqpisI+W0TGqejjUjXqMIrSVml1yeQsapd2359cg258bJp7LR
8p6CyJU18GChLpBgfhBmG4plDKlktzTeRF1Hx0WrRfnfPuEFUyx24D7G9MrHhHgx+3Sa9nPOFO1D
NUCzYty6XwExWdGYlub7vN69Z26ynZJmL0L93laMHn1eUKfK0tGFU4gEofyl7H2cwrggGRPpuPDe
72sSOtmNyp1z24AzA+RLxst5TLj2e4isQEhRb8pW4csspaAKczgYiI5lBxucNEXOC4CcvmozENPS
7QpZ2Mw2ZDSW/vLeQzOdcbYhX5SvjXQ4sCcBQXK4jQj6/6ofcaWE1GLfYcuRUhNrSpZrrMuLXgfr
/iAUfhDI2ZdA8CWkfckFEC8M/pKAIcZgfhIdoqJZAbx4gInBPoUyKIPB2rSa1MRumLhGAtdfwmI8
Xt+8eA6ngRMgd0BhqChu/LD3BDTps+8HTHp2IQUIZj80dAdNrpDNkB/1NikwDQuDCw2EsvIg7he8
4N+WOtido/kxPMOtdwQTnwOPSuez+Z54ve0AhInld667HRWFaE+EQJs691G3rv1QK47gh4jCFpMq
amrdcQ6I0IBtJj5V3MlwZOyQinD27NNxv/E498bk9GExTL3L+Tc2gSMioa0nkg5MUXp2u5B0VoUs
kHnR8gGZQLkantwedbbuujQcBlbP/YZ5lLOAX67O7ZOki8K67awOENwpyw6MIhev4bJ1XkH4YrVb
r6GWQe0YjXipKyCc4RgXIw2gOMlWvuAeQfsw/DPCugbxC/xt6rrwFh5wjBBh6Z0TpbeJupAmTw3h
yzymvTx+OPumIne0+2ZTLcOvXWmpQqu+qnPRVXw6m1RCRGg3Fu63rjGVM/O+SDHwBXqhi1Tkgl5k
EueZwhGTR0fkuK8Y8PPdamEOm52EI2sgkKL/A3tePoBRG9xsqQouA/cShqSP5RGLo60Ry5ZbtVi5
HjPVd0drf4iuWTPGm8gJnhXSo7dDmKiw9xHOFlKsA1jnq/DLjiWHGnpDPyEKNT+uU/Tl79e9W32B
3oyZBd4Qc39+xpwP/5RwNaiuQV12Bawu6PLGmwiGVcrzIjvOI457Ypj9TkJa66UBuWFmi/s5Q05D
IBvZv2pU1wwOdRsaZF5FetCKL0DYMN6QSiDq/nbEya0k9u90WlL5EG9dcfjZoy5KRpghOFO6dKTP
g+jKV/TEiwHE5Kl5f+JOgujucDIgUYWnPNGPbVZFh8n/TRsaA3ydbZTo85aL0AVz23Shp8uowg4w
XP4dzSrq/qnBQBrxTj48fz1xTUn9cyAx/DSAsSnLKMfcR31dMZKxzsanEa3lg/8KJifCG8HxCHbx
sIjAA9M0c52fZXHdxzclUeo+Bc3jwxQPU60si8sC6uFZLFOQBCtXgPrmE0lz+Wkr2gh6IUZJqIkc
YxGkK9w0HFu0UcAKvBPGi4+wVzCe4mrYKAjXjL7MCZ2f6l4p8P01fJtSRmf+C4UrRWwXcyN24NNS
r0WM2FmCleuFhI0xBW0Ev2s4F03ZZP+vkP41uPyWuUTGFcIpeTjuxbblVR8KYbMkP+jeLmPJgeIU
pDxUb2hOJOrwdpQc5AEp2XsWNNS+io5rakRNKHg1Q3NQ2ks2oJMw/i8SJ4iyUmina+l6TKdnIRdV
mMTvABh21TXG4CWMh2IWcu9EHADanSeRg3QXvFX2QP1X2ecOhxMQvlXwj/Bc5P7GoZVorfr1gbK3
EHIej1aMobpEuW6N9DCB5PUskrgGa3xtLgFuaDbzTmgjJ2miUpABjqJNEXmhha5JylAhQyrAjAyK
Abv1gPVSnsBTtCXm7RMkoQZWDDXfhLvPqIJVJBkVBYYyU0Sz9hRYQhsJp7CtaXgU2bocr1BU/C3i
YG5+yY1Xq6gCMpOUG6OC/5iBMxVlXmxv55O2GWKvBin8p8EPb4+gvlFJaZABwQ1OwqYkqP9HRh9X
rPA7vABXlW+UNZklhbWNXoPpd/ccwXCAz22gmuKqE65e6VchHBTPohNcrP1+S0KAMTAU98KVXVaK
TEq2SvKM0Mh8j8rCk2wPSYhVIBQygXOrNrmf6TPxCI7YNqwNcp3mn08uEZT809qRZ9YTJhbmHuOb
YD/CdHwfV0OQhlO8Xj4u+Aub7+fMR4kVn4JU1T1woIhLkO9ps2hZCxON4uQOIzhHAN+p9rbJRmNM
Wj0XqLvz/GMWqQ3D5Yh1SFsGdpSYW34qo+70aQXu8+K3wHJmeg0CILay4ah8W9fvT86ofJuR6OIb
7+OMljaQUh4BxQId0BIhGTnYrJexvVOb58+fqOTKTfr4jP1sHAVcNM9XRYtsXBD163R5Jq4dbYYm
NL0F0u2c8W7OUNbMtVE7CukcOZ8C6Qy4hrRWSbKKDYOFO9LSExk8hgUrK5NgPV7ZMtHVmkUJDkF1
pb5aqIETmKUYl3T/dEAr9Xp+7DiuvkyEHIkdBZqN7jfPjKL13CLqy1ylIMmGXBlxh3ImclS9GK+3
f9KI/ccREGAR48o0GB8xbN8s5J2Lz5PBh/jF93JKgNiw8eoQ8SsdRwSuYhri8BVP/51g7s+UoQZQ
j0MhxQgVEiXhy3XzT01rjUdEepmiWutMeWUx2FUj+4EGCyQ3kIvlkbg8aRRF9Bql9xO5KGgyJ2Nz
W8AKj+4ix9hhFnwdoSpUIlywGd3n9UDLqmFvsjvj0IEg6tSYkwvsGjkGLGkYlU03qYh6FNKVTrdv
cOlqHIw+Ny2MVp85TRGJrHTfihG7Vdpr9yoo3LJzHhJ0w0n+Z15NwCEqfwkk6zDiCsjrfUxC5Jhg
PxaI5OrmDdXtfAlD5D/RLzzPUhki7IEoBBWsjQc1T/MvrgvTqVkack2+FVWfebbrtMi4jSx9oCCO
XTXu/7mLJ859jbPd/FsXgbX3yW2Y2ugnESvB/nqTRrADfzeO+c7g5lSa/YB3tWjHFUl/QQaIQ+LQ
kKC2pzQGGHJnQzYZy9j7LgNzRVYBTFcsRRJAwu+uQ2xcshpLx3sTF0W/H0BA71qWZKM0sQ5uk0W5
YIEPRqRrcQHYR/dtX4JdMCG7YvgudiRaxsAI8o9/nx5Q+FmiyDm+IyyvRwupEUDP4cDon5TszBe3
b0kEmHlQKiFBV4LVnHT/HCfdi4JtrAj99SDGVV5FTrEeSwB36Y8/vjwS152DapUqMc3x5KaJ50g2
8QPpYZcYJDXaqW0Gdf7pjmpVjhhYPkxOp/rNP8fT96YyDzssZwttqMtegfeX1NNX53qPspq9UIU5
RYNhAEVtfo3XXY8k8ovvwk5PO51iWlse2TRO8aa/4HU++8M4PBCpxwgSXdjH6VVCJVHeaOH57WPX
udIN09rHTaqPJGc+QBXltpGBpVm079mrcz5pPJmL+i3KFzToHHBQs8YFGmvBKxYExcNDho9liHno
+U86SRwjPSwlkjJQWYrjBgJO/MEP+PvjF46j/HEuWxVtlxuf3COVpttU0FZLx8e0BVLDU1N8ZjjY
rm00eJthrHkkt4Yc19/RhIqpaoDshjx9pQB0F4jGd7i/jwqnV+UGuSyTVXuDfXPMd45zEspHV/A+
dGbFTvk9tO/n6oT0AUbqK40KKByZzhux2L79f0DUedoMyUw6NYB8PWJ+JHi/GR70NUpeoptdbOo4
ijAjGQLwV9E4Unp4444MOaQAKnueQ19FhEMQl8WPObonN3ezUyDGJ69IRKNyAThZuSuTq0ALTU7r
kVysIHvsMhSDMAQqfqWgq55aiSJhZoSh3ivxkTfpKl04iJc2baXYm7FhhoBn/NHrQgoS8X/EhydE
hBTC6CV8IPpMunbH0J5v9Bdho+wTOuySvrfwEdcerI371/6bzfW8qWaINPnq7OZJ3FXEeryZlsuP
swQazkYDY7sfm8VpgMmyCbYbrUUvTOZX799AZULf77a3xWRgQi01keibkUOvhlpF2zwvpEY1vUyf
CZTvplQWiHx3JxE86Oh4CLqT3jKE8o7QW7YWDjzYOQ5IVrOXvXizGc0vwww0XQZ2XVDYjXX9yGCy
oR5bXfM4xKSNyCOrs/mVM6Q55c0IQSfkv1giNaKT5w7237hE7ZHF5GGwfDO48HRcekCAZNYFA8d+
m8fx/JezRspsSbE3iN3cCLYV2zy/1IPMEFCL96gOODB6hhlk39uZVw+ELTZ6IG4u822o+OcIXqBD
tTJIPFjfVP0/fOHTsgG3nrtt82Lg2Kt+FIyCV7UIZuHupkemsH7lPEepuIPFhK0ZDC58yTtQ3Z2z
cK3jDi7d0sshH1VWEVOA7YAiVmSdeZE93YZHQ3ajLGzxxgz+0A0JrqxjKXnEsq7te8/vmAFm9CpX
hnlO9Fn7RLZum+kfdhwaTlUt5cQFFckCucbsmHT4r2+su1nifB13vqYuJZcSsd+GALjw3sT8WxL6
Y1vWOB51wkWAI2gFR9EZoISkpxz6IRIL1WNSArsgfARKZ7cWSNM8j/CL6usAuzg/behS99O/CwgE
bAeDZZ4n17F+fKk+DXc/V+NHuf01LSbZcdIl65YPsFigaNTuTEZBYbQ7UJ2NSSIdvj1PH1XT3X25
sLxC7WhLDDbYNghgx6a7wU7Upyxlyuq0IQGy+HWnG7XEXmMF431eXo3V6mpdRytLGFjdho0JSqhd
Ed9AJeSpRSXPnF9op9+wXzDsPd5zOiSS5zDFj/g9G+LXyNLHtEC8y7W8scJflbivQZgmOu8m0inr
iuciSe/qh7NBNStRZhV2KngPeFTn2PzG/ryzjmB/6SFg9ngmVUaZm+NDvmnVMSZ3RclgfWbIZVAR
ynd5IV8Y2YbQXh6rFUvEC/krN1h9kA2OUXsUPBGTd1uS1DEufTQ+5H2plfjoE/4f0ofBeUhKZ1eY
DLohkdaT+OYpVYRf6Ol2pX2UhclaC0yOqDPqd3psDrei60aQNoYtFZ8Sa8w0ad8coOWpOgGeHGOH
c+3Efd7aymyo8npM/b8TfL8xfLmadHYd8oBOVwnxWBud4ki1jxv9QWxr5Y2YaxW36Laa1XRo5eo4
pdXrELMD4r/x411bvEUAm8IiOwyCE6uwXkmQ/Id8MAmh8uDgAhKLrpqpzVWBd7Bf1/wQz9JSt7bM
dcJX70qCUl5XtW7HfSwNcjMiVdfL3d1nc9YFd1NTZnebs1LqnSJa/to6q3dQ5FWXNcEc5nxxRIFn
ExCRUUBr5cChDlVKwovG71NePSO8cuRs13EfAPvALzPaxD34jqBRohxVwoHQNx3cL8FER1CJ+4Vq
5u94zdbXgnDlw87rdlJPx6KXXOmHRbts3ELmhAotufYSHato7XiXqeshiW0F1jhDyUQrK9wXkKhr
AMem/KDknxK1+UrtqCdQnszxeKBPOzjfT4lgesHa4sgIbpaxUk/H4gDnewhDn7Ry6tJlvBeIyMJM
okdG3j45OyVQVBAqiy56lS3kMZU2ZvSiYvrrBQIL6RSy6odzzrEzw1xGRyHIrENwgtFVlfR4hjUR
f6M85f92BQ/ZmQDS6AY9NmVLfi9NhuQPfYkyUk2ZQgJGh6x3zlwUGHEaek7jrGDJyajBlc8U8hOZ
LwML/HybFoZPpxEakJJx2NFLwhDcB4037zwNOXuBkLDaF5RKQfCOtbHiZM4HkIkls+SqoajLu/ve
PUcFrpZi5ndwUkcniHK3nf+mFYST7YGQYUTR3TGzT0K2lAU4dddXVIRiS8+5mWWUrTRx21uCSms8
y9ILE6B7MiiEAzuVeLqfdaJ0Mv6gAo8mlPglaiVfgCGZWpoAYKuKsPi1KAPrhYSCpGzCECh6jVQt
QRFvByuuvexPLpOGqHP1YP/vp/HWoF2A2r4RIZZGEfBuyqc9Hhheebh5JeajFUPpQSkWjMRg6EVF
yLDp8FbozDYvGlvUEx4E7lbWClJ722LRQfAYLJde48Zeb8G1BL8ZRkO0BXG7Jv9fpUY/g2rBXnXE
XlFza1+l92ACzdkm8bO97rT+0a5ofO+xm2VJ0Bco8/wgPXw/E6M9m9qEqxif5BgEYyfcbSX5ZWqh
iCAwDNizRADM3ijiKRmP/0sj2uM+PHXy8Xrmhf4x0Gh6o6Q/wwcoOmCPfc0398bka+wdUDoL6Qxa
toOEct6Gvom7rH3eF6oMYIMB8SyReliydsdRfXJayEx0raOiAqSKeK1wEIOnjJIoQMAvFvYx5/C4
CPJ9mh0RDOGbLlKliIQ/MB9qVAmt5Kt0aoW5dv0Xo3kcvzlLmx5NmSrt7nC7gQYUCJAbKj/jtNqr
yjAI0plO8SWcjG9TiHelcvl5OqlMuiLKHP45/SgA8yN5wuY7Sdv+xIRRAUWAJwCMb7zm9DbVZmXn
i2sn1ALo1Rxgkjhef0KQzZuhvp2/PzOuBmRrhblQuzSUCXK8zE9uA6M3teUB07z8tlRSsp+xAbO/
PcXfOhfix6tJXD31axIroyAkqcwj6Ul29cQ0Btj4V7N37xmYV7DpKTo9eIctv8KfEYr+15/Evh2i
uhRF/uWxzIqM/DFvAwO93rMUMcnqOv6wczwy7TfaRRhXmEVFRZ9RIK9YAo4A+rTiSjOKJa5wMOUL
qiHuNV8Y/NMt427Nkd8fPO+0P4nTIEc6csobk/bIUFCkQNFJaEVNjWx2XgEV21GZyHgf/kygSwTM
sEqKlkdR0o2CDk3BtcZYfVGLPwzowWph1bMAYEma3M2tm0okPZoiaGSk3DsSnnorEg9Qp9yy0Icz
orHovHFueAa5wyiDlNdf1/FLDshx9TsJ+ioWg8lTMaHo/wd/0kMHJ80ixxL16GvkLTQJ34bueiFS
OOAwTw6T7yV45cqwHbVbL/9sn+7lThfJ2NL3H2eF6rDLe/2jsoE72UaChNjJMmy/reV5zdRWd7Gs
0nx4HxdK2HJMuWRxdy9L7ZZ9MMOS0P7hE3EtSn9WpyAkstO18U3matqPJu0DtVsAzmPecnhsT7yE
FifxuljAhluzRmpqmI4/CJAglEwirQ7ITvXk9VzG3FBUAFjr2PPy12EkuYMJ1Sd3le4NiXxrRbmF
cHFsAeFFyI5wd1O+vvTrH/aKkMLV/Gz1FvTSi15Q4z+dM3iD2M2kCJUoqoKAsiO+kDFlU85gm4q4
TpG+jsmxbC36rL60Fmiq2pzb06JR2ZcLR/fyGQXozMlob8PQpQlWZbbGANJovSNDp8FMt/Ywj/7u
CdWVKnqK8PQtD8J2wOCo/AWoP1LY+0yLFCd7U+DNogLy6C96U0jgWv1btHiQl+8ubpWI0iOu1GPS
9NgjWbEnVVrChfM0pW/pQYDLlrxlZreThYR7IXtHL84wYtHrvMg6kE5l0ny9gHP0G0aVwOFhnM3d
LEMKM/0gC+xvyNUta5NXZvCv+uvZvHEPBE7BuxMUvX/J1RMI7nDtbGgSEXE8MQx5+GjogGknZSfP
kseTbeqsaxWKFc4kE+UVrswUmCRWfucLG6TBDIqa1/m+N2ICxbJNbi6ZpUAJqbNe8hef8cwdJF+i
yP6n2t/2+5thKstpqmauDuKRQmjFgL5K9hk8aB218aOyHDsRE5vLVXW7xPyXfRobxMUiLPxWJZ4e
uUtp92pJZg/6aGwqozpVZTqno9dniFJNnwfQIEcq41EsEwa4VXnLWFa7HcGmnSIQAZAMbj2e00XV
ohAOy4DDVV5az7DFaOXeMNSLXkMC9jFGNrg3T/RdfnlQb2/CDaF/L0Ne/gnSABOtNX8kXcL7fHMC
hGkQB+ToFF43cS/ZB4r9KmMGADM3epsgjpzkdMBcEoIOLiwgKMyHwDD3DsZfwjJJezVkbkOHKQMd
wUxNieRo0WOzCNaro6agQahGEZtTPtb5M3sRR7g2ySCe2szYzxOyWpEGOl6HCbuRe8j2Mp6xUgWG
zbEh5DeKyOY/yPq3uknK3gqzPh3jMiI51kTKoKBqTB2FClp0RNr9WrQAFZ6bnzIrJLuJGuXH2X9R
Du/G/tNZ50bBdOmwWBMDX3xYTDxxIivE06EYzQp/A3zjr1GkzPk9OPB5UY572jewILgKpmKrsqwZ
XDUiZHf56qx3FPACVtt9eRsXIjYQpleU3Zt1mI1ghg/AmNdQj7//zrBpFrro7oXSvfXzzO18JZJQ
Xh/x/lwbjO2qA1gi5dTDh+94R6bXbMQlpi3JV8fvbyOg499Al0tFGDexJAANXmv/P1Bl9r5OgeJV
QM1UILyhZntSRZOTxk1Gnv7nyLd+HR5S+DK/tsrzZAvWTJR4hLvufAmAAN+nu+U7HFSRuFjcnLB9
T9/VVelTjfWCQd/0Aac4Y5k08qKNrq/nPVnGxOXucpmxCmE0QVASnutpAIWmAaKE7wgV8jtYe/87
DkTLR0CisRg1a4agB2h+a8oYJ2dPiJx/EYl9eaKv9CylKwNrsZM9IUNkRkV2q9dSJvRZez77GAj1
9OLsvIwAhwsnb2u/Ncoofttns3t1hr3k1JrWxWS/0I7NqthjfLfuqAs99uZ0PwwhazVsdJSXKItT
QmutBXwNnBVzZoxTOS/HXFgJfTTnt+DUX/RtN0GdisiCOuQFMIUAESEbvIvuT4Ghm3Bxp+65koTg
Ld0QvVnP6Ihpk3Hyz9LUSsjPoZ2QSaKT2DfPztYsn1jdja8bih6TKssY616YHWqAyphCJ/BCBpl7
dLaUSWlyQnmEPj94Ralt09N5BI8SZZ986MoHv4v+JxBRLndt5jSuNANLCMh55j2yL3I1S3oIJChi
MFWZxhFfMorSujlfmLLULK6qtS7odtaSMDu+aAZdGmVI4iIXwgeb2YATbI3mHks5dWMtCuw9tCfA
q0dKW82BiUoiLlFUAVb1k/VU/a32gN2F17We2U14VoreYd+RVP+kGI1ibT53JHpR0++N7q4QGjm4
TRnuk5eS4YsEmONvGsLk2lvwc4POQDvVHnl6dAzxcVB443JHZAGkF5vWVOVqwlkzT67ApL0YN+0N
hS7U0dKxtz5dVJzYi23ztCRcK8Sfn4dODPnLJ2k+CcI+884lYyiSZQRf1PpcORkdRz8/QOWwwnbj
FQTlbCqfM6BEHaymi/ChwRN+LLg96Zq8hBsfyUvx28JoFD917+b7WnUcgOQ9Cu0uApayjv98vZmU
oF50Z5s9BmSbPpizrco/p7UAZcOsbOuXNXAH7BDr8nqAgRlBpNFUUloz2gYL4kp2X7cpx2B5BLMZ
AgaHm746Dq1fxRiFtM1LtwWOQH6ctQwLJ/x7JRoIxePcUQyLMu8nixkPTZkRZAYwKIPKIAUj29jg
9rTxZe4XdjWMtliGYJvNZAlYC3MyvAccnURIAWiXx0HOeiB7/LGHXFGw4VVYSBzgdGcDOM/M+0dM
wFXnY8Rh0JAnJcRusiNUeiq0QIXTpr5g1P7/AP/rJO5tX0XJmdxiZirs41Sq0vwM0FR341A8UA+8
I5zx36CBI9VvNIq1QJqRwomNriIbHQdohJucGjIY+CvMEKfsFvKbCJK4z5rhW/iEnC/XMA6o0oBO
RkKuDWeDZWuZLxyPt5B+N6WURCQc+BdcEZh4WeWqXtzK9tBhyQ1w4sZGC0CO7gq/oleG5yCSDIWw
ZLiRjTEBlyybyHaJAf3vOCIHpbJ9NJNa9un0aosoH8fciQfLxI10LYraqx5LtL/fTptjM8eircMJ
I0TO5F0daX99WC0d5ThKStddljd226+b7pV/fJs+p916wTbY/i3UuHuGlm6NpBGgQw8qWLnA+9DP
XY+7uwWn7E+yChYrVAIIMEy44eJqhGWSDMSEa2g1EhZliFwugYtv6W86M4O0A85F9xGLhJMRLgMq
d2WDGjuO3wbPVTnffuzlrG0rgwiPyRcjeXpvxVcq3rnG85aoI8fboYMDGw6crhYUur9CpIAr9lHx
aiyWFCFBO0lKlyksLreUo5hshVV3XJc62veGkjGz+C7PXC6aQb7s6PcOFQGSs2dbHOKrmN8RncRG
4RtAzwa3Aa3IzPvHBY2WA8SOkNMFxPG8XYIzZCdSLcu/2o5n+0s1Lc7u2K7CQ/2q6572muKcKQ7x
u3GXHPPLa5L2MzJYffU62oWXBp9eImCaPzPnqWuvlInGcAOScBspo97jBcU4QscFJAZVkUzNzb2t
3tULzL08UDgSGzbkllHP818bpWgnpVPzRQm9ZR0MslyNgyNFXLnPpnufHxImpj60jN0rX6KoWiXr
r/mIQdQrTrLJmBgyBj6uue3fDKqbrah5kqYcfgonKY1wTu7aSdrOu++38hw2naPHriVMEPorQSYi
NN1Tz0qAJg+lXeBn0WLB0J+EsG14mNJiKQY1i78A7EQfgP10pnyT4fXKKizGTObcCRQ0rgTEmp4b
ESR7cUFZ2caChGdCGQPYF86ixBxpVgVJ+QBjP/T+cwKiwovNhJTrQYnrNO5KyPHxo9PXcqpUjd4Z
UhJRXGNZO62V/jVyRg/FRvM4L/8vf5g6L3DZcrmltnAAASqg5lUOoxP4zNnLrLZ7u0PzP7W7CQp9
j5mOBjYnlOk2MSbfbTQjbGuWfU9k029ztKuIM1KA9nnrImf2YR1rFVnuV7Ya0FQiFmpe5KV7Ukno
UXOHHrxeIYcnz/IWn15Zd1WY7qJlgz7vZIaMKLyT/Z/eM9BfO3lD+DVolK+MPkpYOS3MNU3yUSzE
JBDBbR8+9i5dNMALRtPQJPE3L6zIVlJeoeOLmISkq3h2FEKMBs1DOi6CO+KmRhkUq2k9sL89NNcu
ObUVEdUNB7v6sbzfFmPfcGkbwcp6WBFBLhx8q6GQP1TfvXv1JLHiXGPJY88EEabMxfooEqKw3U4Z
EbSWtrBSBbeslEl7ZkcaiHDydulR5/zn6Rx9CF0/AtECr4L4zJgcxz3N4jKfzs8A2qYV22dV8J1l
RdnFYeO4XChT4IxPSFC6ACpmL2MfMULqhRaPgywgRAjRTF8hzMonLNUzRV4RSp1/FH/tQsYY9orE
6SIJ9Vf09U/MvdKhMKXMwYDPdAWwen5B1E9sPb7upcPVo5FH69DF2zWuDQL+03W14XG5GlGHGlzf
jBT80AVLmjLqG4xhMh4akccE5wQz0f1j4aDOEWTsAn37fsonzeMHprhjcdtJ9vLFqxi4mgPnXgeV
8lrBmpFYC1v2GC1qb5dHNkMPsXc0eZIVeRmNNcFKOpMFvLxDVmH1GTayzrTXRjgwSFfvflDnI27T
DsUFps0GTe83kUeAWCnfbnyTZ25ricjxqv36wDvYKMYzW77fUuErznNYCxXPEPouX4POSEEh0M4r
EEg0sDLiAvtE4fdLtw/Zxrxq01KkUFu8qZcNHAS7jRjQ6Da3FTJ+YygndbzZVFdi/SFW/ZkiROqC
7W/5raBixkITeRQrLg5WJT31ZNGO86W+ILruM2xpXpOhAhaUFHU0xg/+uFe06zQ5n5NjKlGw3Dlp
kMapnjYV/3v1z+nnkUQ8atVph0V3pt24G8OzfhCQ9Gy2gz8aARQ7r5CYbnSRfnsfoV9tatqNfrSL
6SVA2uUpFpErKWVg44kaWVwwh9wTNqWWZWTsUZ9kocq8T2kBAhEsAZPXiULzOHHYqe0BpH+YZxEU
hXY6NK4EE5A1yYFFjboMPXlLa+SVdn2DN1Bz2xptCUSGI8NF3kPKwNE3MNOlLH5zJyFkoUfgwcee
EB7B4oeHTvBCfB670u7KomopCHvvg37Yi4ie0WYsDCfn0NWrS9CLRbR/UnF7qcX475nA02oMHJFZ
UtNK0TpjvQDszxl7lEODCgweF8SuW4cL9g4Q21xvgrGx9f1nOaHsG5Ip99GLFpjEeIM3Ua0gLJiS
j/QlnxoKc4llxSfW91yxlEQCf9/1m+aRIlYb8r1ks1w32VfhoLrFcnYzLnZBG/LmyESlrKd7KeJT
ir1BzDKA/Z58ASWB0w0HtDfMBvcpbqbGajePvRs5KXjqUPi62Q1hRDefdnRDziTiFNcc/uDiz1Ca
RzT3ESnioqYQ+eV80CN4o9cYKCtTsyTwL6XJff3EU8erT3uEPaiN0RLwQKPdYkWBpqrDkymzytby
Z1yKZyVRiwEl/2gGGn0eKSy0JytiZNyNhf6118Pa/GYP9wx6c2ya3Q9ciI+Eg0vqsgISnlhViYjW
xhP5psqse5D/gYcCtowcZRfb/VQOi/VIH88k4GJmmvQmCt2vr1FAm4RjRnswlUiKJ/qLkNGV2W+z
pE+wwawBIcXjGn3uZxqGcS3KCGuGF83oPYCVPkWJOr0Qbt26NieefE7TqqmsvFThSiQ0sUPOIbXI
UnItoJxlqTtMhx/vVR2saJAevEzxEoFDEsl2P5ZgxqKJmxMfIpzWwu2z9bdZ8dJYFEfdWbFVMbph
MxuBhJqJ/dsIzFmA68do2iQ8APc9pLr7LMuaqsuSAf9ByRGTj9n8Qs0bKV4rKtvx3qbiOUfuV6H1
TWdsYv+jvbMA3NFJtHmVQy/PCbRySIOZAkZPROFjQtpvBZhx9UUlElvuOxgHKEWaSmqSUOagX5Fd
qGtuw4TVHqKVx8+rMyPVGwOCuBfzIEH3zrvtTd8hxwcxi5wu5S2szHJ60ofA347KfLO5scx/x/dn
OzzrEkcYa6giYB8IfDBM8+Z2H0swoReW+5RMOF5UV+5KyB7Y4L50Oguhq85sbqdgZCXpkRR1ognU
p2n5T4b6qmpZSUu+xnouWFCvFhHf4K/t+EKc1qbD6aB2UKw8xVF9/PHIPhQ3Lue80L00V5TXbx0r
/p9gz51S/xS6R53Cm2fy6H6Or8VGT3aiNqbz/F+nKa4GLtrgCMItviiN76jORHGfjK8Gk26B0/dG
zVLXZKgkNW3vNKHkQROCTFAJqrzLo5GsAsaHjpTqepTI1rQ3okpA8wGyxCRwYrFqOGaN6H2Iq4Bl
lVssVuTWjXhehWs3XR/JQX4LGugFQ01u5PzkZJ+R4yc6826ojYemqnHj/sFUWfwla1zNZN9hQ4zl
azbJNtQ/wzQu2JK4YeTeF5GwoxunxPj/IN+gxSVC6Ek1oDPuN2PbpoZuImbYmtYYUvIku/l0LNSy
vuBmlHAvj6qSZmYxyQC9HqpS8VC2tGzUOavcdrYeJf+LCR1eG/TRw4MIeOqCxSqwcRfqtikCUe7f
OlQcEKT7hAoxRNwtFkSYg9usTwGsr2+z1CTv7+hvGOgK0kCiW+qYXjvbVkgj5NZnxPiSBA9WRmDk
pa7dIJECiT00nn/W27J9tNmHLBsao1nIh1p7S4lhW1+cUOnQixEuFUjnJAjdXyKf9PWhBhVDcZyZ
aQdo4WLK1HCp/UFB1e/V3WUVN0zEgtIQzxexbkinQOTHWJQdXcf6nMAIhhoc+PXg5o7xa8fCzf3v
vjrxhbJOjm5V+huwaqg9su9dBcnn5eTRQcIvzH7Z+hpxOPSgCePjjHNsI1bs8+1y9Zvc7UevEpgN
wXh+2zMnjRgU0ejV01HzkxYbnSpfuPzvMb1Cgvr5rD4X607NyZcpIrFJJQhqFoWjjymdQvi6ni1D
Z2Ca4mjPKB9N6BoQzTCNyHadxlKs7CVFjwXIKQ8tsJ1YBjKAhhuPsziig+BxjhlpPkBbRnVVhNj8
aGFPhTPRaF5gLy7KFpXGuwJNAKAYBziUaHD5jnmBtSu9xIRLStVxgwX4Qnn2gOwtRcEkKt1ZKeKi
ZNV2bvFkue+jjAuqi32o3+hcEK1TVGcL3VoUpvsfMTsAUw4XRGiBGl4d3j7sVbU2bQVPk46NKadU
jyFRhvii1fRMKzv1TNFF6cX+uwRBfsNClh5g945HIYf9rW1ehb0wD8kZhrAoGJ3Ql+FArpW4HnBR
fgzcFu7IUqC8w+KiG6e/KTvqKZiRgDr78Y9hQcd6yhU7KsFZ4wabqUD8/zHQstmWsnZ+nD+/6QfX
vtB306tpx0El0hZ+S5WLmiRpZrCGbVzfYcnFQvY6VufzilQidh4ZnVVWc9uCa++akN1hDWEF0iWg
u3VlrnDIOw8d2f6fChohKcF3R/btWeAIMPujXYK6GiEEp0wAp4D2gWFBdC6C+nrelJCCLSMLwcPY
cCQUwsECc8VwLQfZIB2doZI2UtGwdh9M9ylDMXWNuamdaD2b0xi0rrtr//3Ypoo35HJMks+SHFRf
lkxS9OmLuKyX7Hqs4FTTIQWj26HSgk5I8pL448QWOg0IcWkOKBRYRuHg/T/VsSn1iV1D6EVYKmbD
gLnkYt0G63DY1VA9ZssQi4MfxTfSqDrvtQwHxsHffpkLZVb+rpVHhiv2/fMDyssc7xwbBpPGNi3O
X/RBVlqew7rrwSWHCXFTwGWMavmJsAszahE8mZZPLNk7+B8Bnf8RqHbMd7fifXgiEs7y0Zf1kjB7
ZblJs95fGRCz9vgtDjP/pswkrTs5MsDyYdWOH2XT8fAEP0o96d2uueJ+om61vwatoYWrOSA3CTAe
rwjUIIJ8IrNBkKttVktQaiWeKJUgP7A/RpFq7ja5duNRGwyizX6eWGYJhmsuEYcMaMP2N0A4YcPC
II/6/8lE2Elt4ZGFZQNSstbx2qXccJmlwyt9ypc7dFuygKJytDQZM8SJOLLS5zmZvJSsoLMFzos7
V1of2BXSpt1AsF6fnup241M+C4liEZWhllPmiiGc/hsMLDHev+2wpTohSEkj0oFPvSHJs1sKhWTe
CFYYG2h7mMPRPDx/moB0ldM1jaz0a2dlghnAfuJOo1/QSyloqC7E1uI+N6x4wZt5Tlg7bgeT3z+z
3tgQDiGLSQSyYM67owPNgLNHiKojCer9te9wFFGWvXTWAlv5upYwefsuSm1d/zM6XYPAoPuBYSm1
ZMC5Eh41YGPTp1Glm9HzTn5Fq14dThnigs6/VXu0CwMRakVPPpojY0ZaY4Z2Y1L/nEapeevsczFq
fpuUDu0oUcPNSRa5mbeivPsanQkR1Sy4Y12HINPgtkOh++rgIJiWtZrutkYcsptTInKXw8NFHY4p
P2jeTh09uRj/Va76SW10zYlkp0WD66qU8HrLpw6Xb+SBX+E1XrY7jfuTCzCqmZTUfUx7LwTF5vaM
YNwV/Iyxt9N3NIKwdGNv3mxRc8AvUGTjTgAseKAjnaPknujiM0SOb53BE+aDxhoqF2OkN5Nai55i
YVSrzbt09NFh1kdnb0so214HQSC8j898GuLpMCrcc7yND1WAz1Udi6PzGBK+M3aYQ+rGCOsNaFDf
dMAN09McD6KQQD6hzWb1TUkEBWBi0PTZCV/OT0QaNYI0iBqjqHa3vOWXCKlICrOG8HHTSTAHzgrq
QRfNL5XMGMUJ0tjOeUzJGVXthrCslzc3Ugi4kEwWL69/pXOQuPqSu6r0NSGJMc21j6Ca2CznhlnN
KCRZNcAS+DGI7tUJ2V8GQOWDjpevlG+0b01FiEmXco8ky1i8436zenlEjZIXmi5/9z/tnKzlvwHO
bGM+/o8HZNwd/re4m3GIrWQlHApvtM09zoo1gR3oGT2klxIcdqomn6Iy8LZke4eqE+YOqOJ+muvU
5G2XW9crdNqMyxo5IXKEKVZzS0lISUErH2by8fRysW19lh81YTG+Hy2YJYm2leKHnE2Y8ZD+FQC/
3SmKDG+yPqWZOaAByVShbgqK9olIMnk88w70cXMb91jeLG9W2aZy3KJAl4oiLCRRI6dt9h4BE/DA
YVGOSz3ENxN2GKDvF9zTrRi5FQq6up6U/uYTWyOcScOOt45RkeaQLgxL9TUHT9uEzm7TViIR0oZe
+erXQD9zQ0YNg85pf6OQW1RvN4fNrBM1vvH1FB45pvvMJmo0GHJJ5UEj2QMmRrn+Y4Mbv6Ll3nW0
lXHEGblN2EIjbgg5ClFTiE8X90U8nnDTaAexZGW0zc0caNfqCumcqZh1AZWJMPAuWrB/7F+w1crW
tp5t6Cblt+rRf9NzKfyVP9yroRPp23ebZ8sNf3Ezz/+TdDUwXzv+uG/WRmc9yA0lYxJ+ac4U6oOT
G0x6Ae5ySKbO38DznXTWdzQj03J8dbcOCJ6a+S7YD7rudBTSO+MElI0XuCklfKuP4igUP4EE1RhQ
QCrd4n5TnlfumqfVUWNaMXSTTRua5G9D5NMkXmEvjUHRZEwa9LWckHFlv74AmsauHLp+0NaV4kEV
IUtpMkGMTtYoOOD5dFk+CS5ZFMyCLvAiyq9H6wB9IT1WqyztIx6uOWGylOggLjCn/9H9Z7WMHFeq
acNuPJADRoRTlsKj4LgtuKyoaVNOETdxCYAl/1J3G+rowFlPugJKeBCYyFq9ciuuPwbXMaTUQfOh
IPovA3SceZHwNCiVZwyzMW+UIap85BaUejII1/qECeNAxNgcNRe30eGp8jJfT8RX1eS3VRYE5myD
q9xqSYVnRy0E5UuZbkA3YS+pOfYUa6EkhHuRU8ZrXCU2gTR9PSVrBN/70ipifvKJ3Rd++y3fU+W6
yL//1fHnFcWYPnqhHMmLOz1HonpUFn3m00AtDkKIozYsxVQalB2qzeuCj25fr25H7+iHpopWFy/Z
tCckt1QxA5HBfsHhy4MTzATvk78Ut+cycHpjW2Dy6Bqgr2BYJvNlZokAzZBBDXAv7IGg70FTuu2i
kB38TcW0tWfHu/ws3KHGSZcuVtdNLvYwefBbUGlNnNZSBiAY3g5f2Cr2cMk5QJ+nkmCo6S1uNlKS
v0WSFSbf8vIAg7XrOEPinemQkAM+XC2eP9+aV0FgC4x1pZWWXjXl7sAWorGE0/EGe0W9a3opqJ4M
/eNZqG2tq8TjQyM/Yp1x1v20ZlgtDbaGcts2JDU6cUlsdMNuUYwOCNbUnWDxgmRBobo9zKD5vrPD
gRfWnL8oz2cAyZdUq1zZdKoY51YDv9uEIuLt3CCqxxiZugnTKvhOgiBTzz2HyOEs5sz5nHTN7t2x
+rlPNWwiltwh8mmo8UW/3zcfk5lVrfsRqbGDeLLz7AxlPdlfz7MuVbW0qEXlgT3T/iRMWwEVgLz1
P9dKzNZZQAQIVFQZsl3LaoHOZDFeHaEwsbxp5S9sneCf8jrJS4HJt3i2jA3O39NKnIEx5gwrVlxP
gFJvZLhIom1gG8jnH0/Q7yQqqkkTiApVTOi/9UWOBrE/gWgFxsyGzEaR9XBYSQhaUvDz/PSA9vuz
v5Hk+Ky8Ch0tMjexNCFOkhm19CXRMqckPPmocLSavTwVJAT42Wa5N53LjqWl2qawzWCGb6umzFdK
q/FuGRLwyUAGVZ4JWXg1IGvJ0P5y1cNDMgqfcpmbufZe3ieHW3AFgTTe/txlLq8YnX9vDUc+IE/L
7NjAntlhCqBvM+pQKdiZtmiPNmAM9ozjVFxho2D5kQqCcHr6+ioHkAff9ZXh0mM9ciDpGG3RISeU
7EYB5czXapRlEv82YFC5F+WaWU4i70v4zPrO79aFQkOvTKeNQRi0NDd/Nysubm1nszVTFaGLaWEY
9G7tbg76qww0wI1yKLnODGeofsKLshj+Ag/ywqdVD1YPygsGYWu/7SGSDAV1Gwv3u67vYaVSIY9Z
fqpVHd2MhTnuMV7a9auLVovAsccJkX6xeapIh4Cl9hgolImO24Z2kH7xM9RkKGskKRfV6iK12jws
HdABivYo4j5DZR9/geMTePkduLT0R1v23RtLiQdtJ9fbHEMPafT08BivPWxKBaRuBK2qbHNycQhe
l0iwa7Gnp+b9dQ4FPgX0Y5unQ9nT4pQp5eckP4xa/cQq7L8u6J9V1EVuUJUH+npL3jP4qPEJoQH9
pfGnYhTO+UCWQhEXjozixW1IoLgzepxrRMfZotW66V4AF4kQyCNMo7b7OeEo7E+No/XIDV8Zn9Eh
NfaUk5ADcf1512iczLtR2spPiYgUQezfEGenhd4Q71iPAlxFBOnQN5YJChuS8geIfc9xV6CnaZwC
DsG2xI91jKagHOHcM7UO10VaQUtDRIzKD3AQ5Bb3K+io36sIAvMEfTvNlnOxwqbfVvI1zbbx6tYg
QjtRxMqy5WUlaUdbmTkP+oJdEFmtCUTAzhYTtljC3C3esIyxxkUF3aE4Ks3apGQTV6Anx5Pab3ZV
72Y3NyxkmKcWGNZouA9aafRDPP5Qcr4q7QxXdiF/+B5dM0AlbxK57jRZpRwr7EvqFjJvYIwUU2rR
tIH/16QUHJMsTo3craKadTf+JCdqicEM5j6LW1KNOW5iXnr5+3MIrNh+gh3G9rqHKCAyg1Pba/ZH
Rs5mSlzumJ6JMb4+Iokzk6CZVgEBppZPwFFynCOyCKHTbnYn6ITnxQfR0Yd5QKvIucrUPr0pp/5w
A+fYVhUNiLLsAbYE8LjF/cbEBzgueCvV8F/2anIX/v8ia7qTUtPqIT7RY7paWWKPkMVXekTtsfbr
sQeEVlLqo9ktblbu9vRePIWtg6FKvqlYh/p+epn0PRgEcSQxwYLnjIO65NuHSJcRRZ9GvtfXQNyF
FB6BoY3xpjeNwR7o0tRacWH4NTPiwtS014rQA9YH1sk3GE/VNa1xaQ2HKjeHAuuRd9m60go6FnP3
fN0ZH7KZ/Zpb4MQeKaoBW8YOAr4n4qJF7TugGDTZ14wmDDxy8uBdCtb4+lpvCAk3SE4baIQ6vW8m
dIJ2NDoxTyAUqYQMepYyYFT0OefKy+iuxYBMYOAHKQ7RA4u7P62vVjVMdBMyvYlLlGuzBQbBU4if
QMYxiJ7liH5fgfQjSuTEUULxj4SsfBQH+5fkRxfji1TrZNBWVUjaqyo4gonB/Az3CCzkvD/BeKU4
+D5Sdov6QPmFbobo09Ujs58wK+zduidHuQJ6uiPREFCz50O77Q7OUEQYiB+y/y4RZqq1Pw372nR1
GnvA2LLFozimqPL/GoEYyKVuzt2ddFrd2qLl5s9Jmr3+dXD/zVXtHo5LLkxECCNNoCFHG+3z3kmN
ihXeL5q+8cAW8+JR6A+1ZU6MRcuq7YZqlIg/4PPl/77Y6jGvaK6h4pCrARwSOqbRA29eKzVvf5vk
psJUjY6Hhwvz/TiFnFC9V1wAoaKY2ejvz3dXRWnR6LiE9JbjbphLDzGUe7YAIKg6xdemfZAXduRv
tGC1mizabv3aChweg0jvkWvtfMrldwkzm4nSuiLUy7IvxniKqVNLVaGXRk/jw8DLRDgk4qqYVNDa
TcsnPCmO4KHq4SnTooVP5VJ/hNCgQ3/YSPMN5+J+HPPG80J/zlWvJ8/NbnVPnStTnVDr6rqlZrCh
Uxx+5i1PvTtLTFjVoaP3kigUEy3ab9TzUEFoeF8eAECLtIAsJHJYDo+DaV50gCvbKkzl5IL/gd7i
XuU+f+wqeczorqbJ2DYgnD/OJbKkatpph7mEF2op3NV+7efL9yW//xBRiG/D9m7wHzX/ITtpxOll
gYWrmpNPB9a12dpDlxOsjs5IqV/BwwgFZcWHMOX03yl/gVwrad0YR2rcuPMiRge1wx3/HfOwqQqO
BixkGSVW72Hl/iT3GKyai3cRbSZWCCCHdsYpOVjIOeLzXygUrHfY4lvXRhlMM+XHIT2Y2SJHvaLi
LkoYY9tH0JCeupf76vzis6H865vD9ayZ7FSua1u2Z6xEYH7UdYBveG5toUNvMk0nOxkxr6l7AsOM
3IydGYlCCaamInd3qsNpm/18CGI+Dk66UWG9znUbtyxf3J4jcOPZ2ueEcKTH9+/qZGz0Wttp488M
HGDzXR6gnB0wYknEPOX9FSLi2/3XghiVhjBzdenccczM0KwfLAhgA8ABNZJ11TVYw9YPBpftccAV
XS4/V0otrFZouv8KU8QvgyA7rWmrSTswgRd0ngDosKPQJ1sRiSNan6Uc2chM2HnHbvB3zNpkTzwS
K0H8RxGwbpJdlwKN1z+VDzUwvlI4ryuoB0Ao0rxNdVV0CNcBfGeDwaGrU8C8r7nqamAma+1OLjnn
PQFmlWSl6rPWlz8I6eoPE4UQtYiLTDz6Czz98a00c/f5BjL5iXofuxXmUdmyPPmQD0hdllo4tG20
qeDcQ+KQuomyzrj7usryKa2vI93xzOc3wDXjRrwnmj0ozigMRk9v6u6a25NEduSKD3re3nKbj53h
txuuXpgBneMiGnDSJ6GJHhB/BOfQeMTdzOniwaF4Ueg5sytF8GYqmp/ccPFD+jh4fq0n1L+VbxJh
wAQ2m/v08z0jpIrZe1CVe8hEz0qcJiSbOXvZ5qi0HkTJXJLB+9Z2RnujnAeEQ+F0AMVclZDUlyGW
cXyRJkTu+qbjNdTLYNlataK1Ik9EPOAqlxrQpOvTnMLxSxTtpqJ0VoX2fxRa59dDobgb6ho9Q4GV
Y8wZqWrEllM75CyfzNr9SSQ/ANxhoaMw5yrrCT5rpe2CDWKvIN1EwZQBlYjgELTuJPbkas2HlzUy
1tkFf+SLl+S9fvpFi7lXUeELQqu2M9oa8Z9ZT+JwL7O7chKgVQXUOyS3M719kDBfgZ3xMSWIRBO7
GDlTtr91NeHrc+/h9YGd1YZMWzeDElT2IWiKkd5t5IFBEYnZ0Y2E4TFUILFwa7sbJ8hlKGlzuEjm
2J7X+5RyVhfbZXymHMYcmWdf/fKf5moqxJk675JTWBF3OdDiqBa4ngUjwvpKJVCgvRQEhYobz8XO
/5X7/SyT23qp0LsmgsMb5zgKwbH9G9qbucWxsJ9OEfL0+z1vmjOCK1UKqEuQ/709X78oNfxHalF4
ye4GKsKlg/vo33ORZPqi9tZ33pT9ax6R/iZO7THsLwwTDPD3hl/pjkZcacRJFNva32ECM8WnOJcb
qM6+9+jS+CbNHLBazD+ROkqYdRZi0+fZbVf6qGw/qomqj4tzKOlugr9RPdJd5hdbMDkrgk/p+kwB
wRx+sBQECnb22GST3LIUFflzJJZBhH51qVOk3mboDsaHJEXEm077BhEwkRbJ5xxFC9LmmZEIbrv9
xrUv5ywXVtExXt0FRtwWCwu2AMvd83r8lvPzwPu/UZCaLeymq5kIHlI1X60w5yTmhiPEohyzhGd6
UZdUGt5/oYV9tEAVVHYEj5TondNFhExZGcfGpLnP4dhpRaqCP1gp/uphHdhS6xzzTxGrduOg5lpx
xxa8WeYqqK+VpbM7mshan+tzKoJ2em4fuj3DuGZRt4dWVRYf6xCBrNBUERIXRY2W564V1aCoKdve
DCtnlzK1Ys6pNDT+Fgd4Z1VWLp41bdqmMsw/hY/XVm2Jk/b1Z7QbRoOvSM6z69KQDU93L6Rq5rUt
thC0aNvUlMHgcsYxXp7n7wJMlIhw+nBRt4PBq8klAhtFU7UyntzztNohbSDPpiMn/KUVKZRIaZHt
KMz70KgTLoeaX0JFnoWS2fmNkg4zLzuyr7B75vrGplTPA+yNOaHqRv3kpCrKLiEDiXVIpJD1XSmS
oeBPWgwXljxyPhwyVqQ+/PbjF2IW3YKGFqbCdGpRhzcSEhXwL++mI6jFpkhtCLxj6YXh7hdKYq+T
eeXDCtlXv1PI7xXYb2iXieddpleD15fFfcbdpxUJ91LI0FVPVrWoXGoa4Mx1xsbObFkjVF5tIzun
djRb6aVd19D57I5Dky3M80OLZPxHiht/m8s2awGOY93VV8tT92kocILTWQLviuLwJWMxB2TbdHg5
93wh1scE22Dow4Rjc2v9CnDEtJJhgBbcQ35sjwaFduFL0ZxzaDsvxVOl7lSJxpyvrtvMGV54hg1u
FeiBzkvjeXegJyGxw4/oSClMETT0jmPRr78COGzONecjK9lTvaK4VhAqIdvKFQWeZoKgTB/rArfm
4JX0ibF0UBS3LorURf3n6O9h05uJXnltpzGI+/rnZdL9E5LAWlT/J3nerqQwGNTDoVNz87sO4baN
oHHcAXTeZ+7PQMLkOUIQQ30s/lBZONBQPHxZviVAOFGEkV8lg+wGdlzJqngDmxRjR2jlH21xzdRO
C0sHWOW7Dtnq6c7Vmy1wqyzncX6jM4tRefaOdLcMzujx3IGZWCcVBnEJahoeHKhCSE9309sftUa2
kmoeM2w6Y7bluzhEeBD1p9ChMrRITiYXIlBS3IEFavZyiLOFo+RYvNY1XNLwxFQhOh0oLpQkSGFI
uOTcU8n7hm8FFpADHX027PhjBg2RtE5as5iA0xe5oqemd1Fc/dGEhUqTfKdyoAmjnL5O08BeBnmJ
qtbwlEP62pdaNyL64N3VrbFiQK65s+JlVXd4hSRLF4hNuU1IIqJlC3UcinHhZhgBu4MKsSaK/wzL
DTztidr04QQ8G5mjbQKCohpJPxY80wMkJjZSLdZMX+WRdgDs2oVz//ePo5QeRky1NOGh324KVjUI
9Wt8hXhmRH+me0KRCAGu+LJ/dQg2d2HT5DnI0TpZqWNsHxmSFMYH5b8EtciATBIuPW3T1JZL0Dn8
wOz9zUXErlirN5jWRRfM1Qk1OE8IuzFyK1Lr2aaobk5VEPJbfVBRKxPXuzHUXRlyeiu05GOJ3FQf
+x2WugD7Dx8SF5TrvaxTyveF3s82VElEvUorMrk3XhI9htWcFLgsARtQPXKKtopm92LLzGSsne7b
GQrltWRYRuHapsx5pS/vQwcm3kDVJRcTYddxXuebFawXXuaLwMD4W/IQ6g1/8qtelSrsU67g3QJO
QwFemvEzQ6wqZPjq3jnhl6yNbKYWcEiwoTp5NGWe+Ozpnwe80YpUpcNkr1qa7xD5nlwx+jCV1ekC
Oy5duFqZrWe+PhaE6Fu4RhSCkkKpLZRIIgRmgZ6qCFE9/WFvsPf7waU9PwbBcLl4YjMjZVNb9z2k
U1zSM5h1q/Nha5sKapIomUYFJoF0GlS4nNxnOei3wTHlDGFr8pkmyD1hi+202K4EvzXpD5WIHT7x
d4IXLpmXdVwKC53GeAEybrFo9mjqDCYPAU6YWydBJzo0f2detfC8boVH02ssSx44KUjsKeRoxvTH
MZxp8SAOy5zBXVAczDOsA/9KmE4ZvxfeIB7kFryup7R8PhmSpzqCb0ZnNr25TthlJY6WIZWUoG+e
jy1egt3ItBVMQIu/6pAjRIkAVNwGPT0ckTMFO9DltxVOoZntFqUvp3rcY16kuhiPaGj+cUxlP/iM
IbzeNO14h3cu39yyG8hlMW0/5vEigq2DEhQobe3G08kubnUP1Q09vF9NfAieGcqsn+haJzCfHNls
jOqAKciUm/jOm7GcWMsoFKqkivWuEPzxWBack2BKwX1KaEk35W/pKi9ZOOFJtXzEy+du+YgCXvbr
2JaJWKm2JDBx3a9YPfMMa0qyAsmMt61nMDiNLh0HEhKSlK4gvDURzcZIIgvG6yYhqcjv9gMB2UUA
Me+g5Rtt3DSCTHLnejB2MNcMxEOI9ZVKguB9MEMycurKY0m8cGFNOK5UCX36GZt6q0e04BkX5H6U
G3ASP5tIBTwZGgEvQvhNRQqeb55eWuM29KkDXPdq49t9BK3jvN4CSu/sM6eoVrwdYXnNX9Kk7zPM
ISlAW8nPyvJZqWDrG/8wk/zeiEx0I9Gr63ZaA2My5kyFJlGII3UQ0ha+RtvO3o0ocel/4ieF57gc
j2Xdi1xzxN80aYy6DyBxQeX7OcUcsTyWnjAKtUKmcevtiYnJG9ZOrfn0SbgLy6090toFo4ohVSN/
NNkM2W/jjX0YTS1Bydf50dZiERNgOdPQ0HSb0fzKRj9jwqYN7MM42VIB7T5oWGnoJwcZQR698Ro7
464AA01uok0h/wIgiTvvSBC0s7ExVMVNWKvnw83BOh2PNbfKedbVzTcJqNhUTlZZuLxzgy+J2Elb
HR0YouTAKwHcsIp2jWEol/ZxkgOjfYKq7kGG2oAMEtyKsKLjycFBRLZdnb5hug3keEnXYx5+Hc+y
DQQpxN0gNZt7Fkeq4Jsj47AiJxOeBxtUcO5XA7pehCvO18inzTQurpww8Nt+Do1SxEqzJgDfNAed
x99yKMllQ84YgOZB/+S0GaE2lF/NTaaM8TuxuNBrCsOU5VoDc3VesPxqwV0c0OpeAeP8adgHTo7X
h2nwHABWV4w3CxuXCp62zr/c/1d1OPMUtkqbmu3RAbxvEMZXCyo9BzDi0MZ13EpgW5PgV4KIIpL1
5OHqmljU5sbwpKhQpSyhK4xsn8dmvV/FHZ+3dnbh+NsLbbwUbqmhgv9hgmWhjn+6iTJHFCQx4dY7
yeo113THormbNG2626Z72piQsC1qBfFfu+9QI6ZCkr4IjmjwQ7qTSn0GChNzAdI/48+3fsVTcOik
8MGtnKiSH7rLKBHhmt8q4iIHDoZ6vX9XXV7OLrJ73FK/l9tYtQnLk+xOfLtspORUoWGEcEfHZ/6b
iuqTygl/7RacQNzTCVuAs27/5cMq68fjTL+wB4GzpAzawhG/d9yhsympf+8bhhcatdK1bhl8vQHI
pLOUcDu2LyvB43IrpG13Rblv9qthe7ZaPOcR+NhLO7Ykxh9/sJxCc5/vCjHKKe9oT5K8kPj+6kQw
jKDuaOsxcG3K/mA2nRtIwKVM/ji6p2VJaawMugWyzm3f62yP7zQzslbvtwnGHewoSZptHg53O+Fr
QpxVa0AAtf0ZXcrgJ+zpgMWNHzhXFjWrTOZ85dAvtk8vmbTNwz2dXuFdEPxeGybjb3xm3sqceOEb
SFkUjhvhsgZ2zJ+883rpUb5b0yrEfLCUG6/9/eLzMt5uGw3262d3deg5rpUdCRCBSsv76geNN0bI
hzvzqnT3Q1PKCn5FXuQa0c6BBlrsjUoy8jf5EY93hta3OZHH5iUMGbG2h48jLIouRumHYqoyTHsm
6orkdmv7uDMiY/ggrusQd5uwmHtiT4ToiofkXRzAXnutikQEm6rAosLP0EsqnZloWHJp1IuVe4lV
yAiUJZrYlCD3lwZ6KwGv6WkRreY0wtYJ78URg//R4PXaWfYPBEVPDRvwD+bQHfCt1o+TBSJyv76R
n+3LL6QB5mLSz2A0bu9GreRYEztwhltwMW7w2TkkX2mNTUxVC3qCamOFsIc0bLYq4ucKZT7ldWtm
jtqdIaATwCiungBplqNFz7zIp0AbAUonz2j6mC6fZyoKVh0yH5qgggYY6KLH3KqwgKzS4f+TjSPU
hqGkqbX47WyJHaiPbUhiwALs/kvLlCbNcouIODwfgAITeSBtJGcY4VtUKt+qk1e28tLixdtRDZxu
N4ED7WzhwaYuzJ7YwjYg44A7A3KgzH70foK03asdTfsv1/X5/SWYyk0I9bKYl1siuCupEQ4fL8fh
NNBv2/x8IxY55azBlFmr43cP+KqKOtI76EOCWjLrKDN+5nMaQ3bRxXZiaKt9A5err1/zOuJBz1rI
JT3OkuIPJ5OjfM3DMV4bmTbR24TRbE5leGmgFB+qqTczOUNQr8gupoYlKONFXLknbn7pgNGEwHry
GWfHANieF1vcka6YXixf6quHvd5QrCT3zCsyWXGjagk+SLHvFYqrgBIu/9I0vMLmeGwlt8zvXmTT
RUH/LXWgf6P5SkgzcLaRKX1RtjoA81cyg+HNGfeMeTu/iAUA3HWnUYwgIfWKe8WedoR46Wul4Zie
2QoaBX52gq2K56BuyDVu2jlHP1rgPJ47j5S4X4jhsoUSdFMqsQAt7hQIXntUZcTkIJzYYhRZbChs
RUK6KLbUfVDJAZg7aDvMIdPADCR5PEGwF+R9oPmMzI+P7HulmR4/5EHYlwFRFR4rJdxo3f6Mh8PK
A5nuWbgNtfQDSYgDww/UWAJj3e3qeu7ziVLCYEE47kf4dHetY7hom9FEgMLhE/qE4S70GUcqEE4i
WIsRXQcKHuFSP+BHfwNtN2PJR0yS1nyf4e/4a76DCzLMr7UUwSND4CLbgds2tMMPw2JFwE1cLEHd
oNUtrrmgP+Wt1+x0B7Pe/PvrzmhM4ff65dSUKGcF+uJeh8A2mCoJRhl9S1mJT7EvKeOVmV040QzZ
mmWAfHaHuqtTpCNZAEvKMyqvxLRuEpzlUI3BGiu3Z1YY59W3WLCHCXgF69TQJOIrtBNyoM6h64v7
go44p9Q0gMLstUfgk0uRL1H64A1R3wqLoJ66t+Y7JfFUXiw6q4obvErDm7kqQ8jTFnvObW3JRelH
AWJmA/ZStnwqCjQC3dZRA+RKHm4ia62sgKVX1Pqqr+4ORgPFjhW7sUGZUQh8n6s/UpMRtLZAdDZU
vpPvbzLdnHZh+zYYbwIQkVWlyLnrURWOSZsWBqudu1rNhD42+2R5W1Vf39B96hdg5rgAKhDs6/M2
QfHjE72NVhpZ89PCUqz/mh4wpP9G8MX+tyENkn3BRBDaX9dOpTGrwOHRq2dBRKC4He1BlmHadyKp
a8woj1FK6iuw6VlBtlDNAy4Ft4SZ4nTKwA/Mm2KEincBt/tY/u9GqIk7JzuudtBwjH/+3H6SUocN
b9SyNB/5Oa1CQ5Kl8XfZl/Zk3YnkcBvj/cbgiHkv14k5RjsZDfDUNpMEqU4Dr0qJXx5B1Gfmrnvd
M5B65Mfj/jNK/6tpiJJ4wAO2o/F+5SwZqKQHeARzp5pZ0iTWrcDiXYF0Qn7/YGuhQdUXzxX5ffdI
klD2zgh4UnEzAK1Brnz479O/8XWqRng6DQgbVH4KbxhX9a/xS6XSZLlFt8kbAIide2Gtx2W2vj70
Py6jv5sVbDtNpkgfBG4m7dgaPPhp6VztZ6ujyOY2QSPjCnF3pkGVv5S381YppZ3cFu3Fu9Q5Jzz/
cTe9QHlMxmwh+u3fu3CYBYIltSG3axtg7aS05h2X/qc82n7YMVCr1WyvjLHgPxZEW2x0CTEPMbXv
thPx1BGpqToq/t78zbcCBlKQCB6x+o/ptZjUzE+SZAZYPsqx/6VpnDEobHXwLlmhZSOzgoYso4Pv
Do3ARZbKN5WmS51s6zFgNymvIwAjAv0DDuU7AnROebKj3SK9qJnGVHFLMKrQ4fn5zZBPsvZhhwF4
2mFHiRyLxOx6n42RiOsYStApe9b7jBb/OfpSPkxKAQ1kQDZESh2CsjVs5ETqgRxD2RhpQzHPkIm8
stelx/nvIogHZYXEODoG/szfyqkRmm2fOkBxP/XS31WQKNAWuKMR+Pu3gptdgJE0qQn10nf5t6pH
wXMyrzGd6VYTZH8SYCoMEnNojnRdDmQ5jNAxa2AOxhwB6sHG/WZqBDY8V2aHzM0EAv4BTzSPEB0l
0cXnSzl4jwMZlUELmpTXc9u49rbY0tSZJdurVq1vqbCfuYR3yaTo0O53x+6q41aF3sr1w7uz0ZI5
NUiosDsEFI0KoC8ZtR4JiOytwhgi/z21r9OwBRHwq22Kd02makDhTDAizZAiPIGkJIdJwPZoD/Dh
FH7sTygxqrXdGkD0dU1rYESc24sAc9EkUds5IBfUDsGHg2cNSuYlDSEGoruONa3Z7l1QpoupiZek
0O/nSALtcWQ/UYLfx4Fu5u3dbRw1NGl/LwCiSDVnTjbPFT3nou7q66umVGkkIbaL4jmQr6tutDsM
cRmaoFJ3ukHr0gmvCctX55szlNVta+abTfrT0FlHqPE3FKr0LPWdnyCzYuES16k49NhvrvuUP+ss
BcX6ou2gWDyWMqTAyFvptPdDALRvmlJsS1IToD/tUd+6D3OXxjXmhuMv1yuZoJIA/zpZNtInKBHH
X9bZdCjCYb5m2Pfw59HX5izfotswYUszi/1tetpFeI3Qy9dfDeDf0/J3OCFd80DK+TcHaWzCGoZy
BZ9UG7R1ZEpnAqeYLUyWWd0uTL9dGbeZp0Wk9lV3Jib2sS3sGWAkXx3FhUJ7pf9enDf8bKzks0jl
GlAMKkauaNykcecI6DpooxjCBsbbReMTAI5klKdU45AeEYiF6tcc0410xxbSSTktOrtHuLbmPZ7C
pVpt8rqzHC5LUQAlO/UZ4WRxxpr8gfxMqtsEAWXnMkVgcVUN83KOiUol1vOrq1BUsNJfd/ouiBLE
pK/7HQ+lEISh5ZUEbSumQhY92Mz2X8m39fitHVOX/133IDLrTPmUURN8nWv6N7+gD8IwtU1kixBh
b5OT0mfxk7YIngo/8nHjuS+r3q2qnHNqkWeG+ovzO97p8FAmixdN9dNuPnbBmgsUXMcKy4SynwOL
zLyfet8q/V7Mf31jaXs7kcCs89XrEjTb2qMp9TCJ4omVka6b9KyteOJAGpqfuL/TdEw4nIAXjIB6
A8mn6TH/65hbU3eFufEJiKB82yH7HCRrJZedbZq+46PQBbXuAM3+w0VgqJ0w6s7MIUJbME+zsa2C
fZuEhkGoqPvXtAoitUUunIqiBY8Qo/q/aUa10d4SDXGOdflp6csvPdo4VxNpk3wdibmzGdY6ryyl
Skg1Ey2+icLRAHMXdFXqvG289nvgfSWMLAVCtaSVkL9d/EsdaTTnnbeJd+J2tl0bpKkqZ5bxzPkB
UJRmlJBr3hSq8MJ/o6HArD8BnQ4pP123TT+tVweARgTHKTo04bAKqRKUi8jEj9wUuSQ1mzOck8R8
mQF6++7ZM7pWM3XhKQ/vV0bMRtm3TvY6MPxFJyKeCNiPeZAQyGk9MFlQWIynYOteCxMis8PP6oMj
e2+Cce8mkoDac8/gpfItBo9g7C4hYBP6sbPVFcyrVnuvqEyi8AfvonCvSAGv2tmjkptyN1NeNesH
HTPho7tPKVkCzFwx/xkXAS5GCOXEUjdXOFDlzfvqbpfcOyLPV4g/eLLR2WW7syq06ACryng9WoK2
Btlxn+9H9ei/vowsCqzXZ/gCyiaFFFTnDXZSCBoDvXQNtS5yvTuNUr6sJogxk3j7a5uJEzNFyOBz
hZEW5eVkdEtCyRnQKFwD2NubHt97jjnbHXTqa16LN/9rTXJqixGra3kDp2/8LPz8bNMNF13mlDAK
LLSzVGAoBmCFw04SrZ1tpGO4tsXN3nL3IuzXr2WZjc/dRfZ73ImyKaHs90sKQ/aB01UvDXE994Yq
bQjo9fiXL+dDEZvtNDlFI20H6Y56WfvURKngW8LIQgDTVzQZixWeGM6GIih8RahA181+WanRtcS5
8iQiB4XEX/VmHgTKZ3toWccN6rmfvP/iI42nta9PeXnPHf3bognYwPlUa56wy2pISEtMMgBaO6Dn
6j2deyUBXGwE7QDC1tsYPsTvTeF7/0xPmOHyPOSQbZmOfMStV9G33L9nJzJmLV//dAQGj2I80i4q
Bp8fIyxcgrgcyX92RTSBjY49/TMozvKeiH9wvLdIWltJOzrOK6lfovDhJaqtZzuw77ZldGR/xJu/
xuH/4pwMKbEsickPr7ejdKO7AufhmfjxIUiDu0RwucV7cm3N041hqnJ2IXVvEaxs+ClLvnbx+V8r
D+lIHshaeJn95HJn5dC9gMDEVUQzml5fQGhP3pp9tGlZkLADLSqVsdRgqoNRY5YoKMs7bquGu7t3
BucI21ejcINIc7zUfv8uxvNBlAsG27T3y/wqRy6cKYNqUvWQbbuh5GcJ7IanRanRdFsqA7WkHY88
LDtcv9k8PHGzqtgECeAOwa/4nykefp94MFeco95LkNAeC4t0R2AeyBNh/zFl6pwsQuyRnjt/aCNv
G5BYiA+/lDbE7edMjidTwg7vC674WDwg5QeKLEN4O5jqDgeLOP1RFWBcnJlRfEdg5ol4LS2krNKk
xQD+Ew3Zx1lSbdGIxufZY6ST8WiaUgbEhC9eikfzaGfJd15aKtonYaBQQfb+YSU2Q9BgRZUO50mN
9F8uZL/sUMCmEcR5KvgALVnRoXbfBez+T9NnPRqeOusKsy/ppCjB/Ga5AtSr3fx2bbxH8C9FspLf
oX8ke5jeZv90zCpnOFUNNqvkFc17q7rBv0YeXXf7EyBllWVoATHstyDGTKTRPAcxip0OFKtjpoGN
L80A9mzpUFfsKWyZF8G15CKveI0gnZY+T0tbV98SQyvH2PvxJXvNb2vjwRj9jTynjMo1MSSCFTiQ
mM+DygBPT8HnA6+bMjfIV+AVyCIEU+0nyqoZZKcmvpaM9fu5BTmX+hgraiIad9uBJOGfZ4WJKagB
4okd5/FYUI5uzhKHBz0m5nEXU1vkUDNAAWt4vDoDDuagOO6Dwc8MSQWf6aEPV6XccslHexIPr6zq
UGdo932TZtIHdX2T/l8xYTkw8iUhYyHRFZR6pC3OQMMiCkcA6uTMshxtQGM7omiFJMTYy9UaQ+b1
qGxDfUj1jnL6OzbjcJpaCwTk+eCDObusNREEmacz9zlKNjueiUVsWzJ/wfC8nwGmZG9QD67SWj0z
i041ese5FX0aDf8xPKd6Aw/6jccWzkU2TZfLn6TPN+CCOjJUuGVmD9VTKXqC60zeaU/EsYKaPWIJ
XdlqQUQp9UgkHSnjf8VeAeuTtbiubNWK2dsk4hji6aVC2v3X4GMQDMm2tz1E9GVV8LW1XCKD0RqG
vrEjBHUIILLlsDH6OVCnE+kj2OEKjQphQ8UFPInxU4anogQj0mK2/6bWIlyxiA4rzRIKbMxspyY9
jGsrd15oyYQt6B4MSfxg23qVRp0id+UrT/O1WYVpfFBwS0IwDrtXyGFIovDeo7XTdvrAkrsLY8Cr
83V0r1Lj3p23Z/uLC/yUtYT/MPiAchmr8n37dm/KiK8hBBjr6HJ4bJhezDk4HZoxj2SgUvbjvC50
Y02aXsHUeZav6P9hW3MCp8O9Y9c0hJbr8ubIzRRm+HOHhBI4n0Bo39je0zUfuffZxSbtNpnmAzlO
TN1H7ihcCWHcAkfqWUs39cTzxCkFlycAjaVQCjL/zEodcdtgIQWr3ztEoV42rhNTRTxQWlvApv0T
JwVVG4nQW78L8lwvFlRxOX1OMyfQgbNsEfSNejMpCoSK11YJF4oKcKldXU7Byzdh1sa9XvYcbuk5
qP8pW5peiIJnbDgwByNC/ZtliMxc4PPx66zG8Mq9kE25jp7sVM92JL2Fj6UtCJeakmfJ+blAm/LB
HljxKgexgaYPfUqraviHqrXDjliN5XN0AVwkXcQNs4TGEQdf5g+xO9/nXyWq7btbCCuY2UAR/ET9
Qzxn4ulE+2fnVRJIHQHK/IFO8PCmiiGDSPIGxeo2LvBUYfy4Tj2JCkZz6ToRWcsyp1N8VGymWzTr
xc+F/lThaGZ70Y+soktpW6KGSgsUXUqjF44IweNnE8VW8+95nROFXqVqfmNvENrfpL6UdBB7yhQf
qMpN8V3Fgf7KA4rCnvS51Rf0tEjS9XvQhkIsHsNMtNWF28ipdSwbtO6MGkpFkSEiQa3NzK761X4D
9FD+uWrZ4MS6G5VX9fI6fnWgaeUO/SqQTMFkDSKsSx/Bqbebgy59nG0TRT8pXylnQYontcSxQKSl
4+oSnHt73c9jQ+KrvcdTJzA5WQU7mE6UNvA+IgNgvLM4dFxyERKmqJp7QhFg57+vdRqtf35fpChQ
XWgbDS0yidOJ0P4zo5j3v+YWWZ1KaNA3f3mxAjrxtDpeEZAdBP7Fr6v/4i9NdWtz7N1UaTQCijHo
CCQ2Rvh6QTMMruvjTFgfokKx/34umbziBZxq9CsgOdGCSZA91y+ByC5DNbJLJne+Krjh9D4GAkid
fCDr/szMTtpoOV0EdPB7/vVtQEOWQqL+36XPZxtUmpgrG/v+FjhQI/roy6FafbuXVNrPBL3tfr+u
h+6RTpfckqh8eBJxDmHKmlAdm+iCPqxoBMLrWryCc0n7WyRzHzzTlR1VZwHdwlCKeriEAyp5F6H+
SmjcsI04s9qOrZUmOCSVBDNX1iVNJz72jVLhOk1L1TT6uYVCSEOYr1Fm0LPLhdzgJFqYDnlpH8S3
ug5pDyyTXBBshQEJwCPztXqgFZOoQugbWjhjegC0A32aTTmwz71ZZdNul8c4+bf0xwp3xtukz1GK
lo1u8f+VWt5dZoldFcYY9uaseRS8geKIW42I2jG2B2+5o3rlwfPWY2u2DJfYY+DN463cTsObw50B
/CWb1FkyPVjaSyAIx9hCxXmgAuSWNmqlByigEyn1GJf/BW2AKr1spie/h4laCd0BBaDYqKFb3D9/
dDaqjj7qCqaclQEjpSBGBOaAm6dnKGBeKtFcvI+1C1nTQB5OHZwSGEp2qTuM1syV7VOQe5nNaesF
4waGc0fLb9Wfogfdnsdy7vaGAtaEc92KSXO+bt4j80vqDtrm8STJd3gLhdScQ9oAXTboMgqtR2X4
XfjS9+8QBpX9BA0C5R9D09TH+pS300eOkCCT7QVkrk3ARiLako0CDqMtfKGI9wyyRi2W2XzIhLBs
1DmQMI5q5gMiHT7IEqu9XbKjYN9rQsuHmCZ8uFd1x2Qa9JN1575GDWUNVqcPKAiAZL7AvEcBq8hz
Z53L0UMjVFwF8ib69+OiN1bk0PQnx6LbOVQnNtmA9AZJlt3OzBOpOBMbOS45w29++gKvN+h2jOs9
U43d2R363/S2VgI6wnjcWwQAEJ1QY9u4bZS7bIv2oXGhJJCtuVodWfm0i4XIM6s+2i5AMhz6U415
R0+zCCzm3dvVGK37jX2DebiB+M+JuJHsjfAbrugky6peeG6h/mvUIY27NfKDE8jr+kcUEXJte5ky
WKXYVVjNUz7kAkiZtvx9vtU1BmXnzUXT83kTtSyK6p2QaWg2PGtrJhclATnxdz7ibxiAktUaWOQV
BNyOt+xX/7JmASiHtGgrZByj5epvR9jO84Yf+sbbTTqMeZX/Oo4EIHT3eV3VVB1C/LLIVklbJto5
xIET7oXpstZGR1CO1VJXOzB3vacynsMlJO6bdlr9ThOOiJj89tdWutiyOhkfACsiV+VD6YMgGCv0
iUih/n1iWSIz4Ly9ydfNAuv6zao1dVU1PNvJH7v9NyqD+a3DJppxyWr8NTAjmLWY1nvp6mn+qZJx
ydWSbCIUc/gAWjaIevCph4AE5WJXalR+WLxENi6jkTM0PrvFtNRcAjdh6gVlm+l46dGPQ65+jjM2
pkysTnyN5TNecAEjXRljz9O21e3J51AH3N9LDO6aVOlZGxpMP0ckDelWNIJCEfz9HYQ3G/ziwUs0
IHN9Hxk6mCxM6rf7QWfdqlLmENHoZ7N1KR7TEahLKfbBEswp8hYSIDbx2WNSufZtm8zqeNkQr2qY
871VM/RJ6OPbmdNONgkzgP1JYdpM8KeFGrUXRdjP9AdlI4zwfopE1aQ3aLO+6viJ29VXf8kSc3HN
5yp899EArDCC1lJkmUVWa2ShsOApoxyyrEAFKehsNMhTB8nC+AXGNVcUEGTDFmLiSxO9+9FsyrPo
yAgjrUE5jigaHhlz6fHcJMLt99PIpLAk03IGRaf5/XukkaNjdghFLQ5JzmELjxOxufW5ir+Grd5T
3H/GStOahZEKBbpdH+AqpWeKrGqkRC84vFPppxbaXWrzHeHZ3bt58mhAJsazECfSVWPKWQCkdLP8
lMYJH7E2Mv7gb+s5MUYsVHNZqKQUTx0IHHJ3+rqT5MH95XiXbFfuxMYXOtfhes3IoA7R0/KcPdCY
0U4hgpgrNd7E8i0291d1aNxPwq65uO9Ynd1tmp2qV7Bu/IHzjHaMDqOoD2cn2xpTmBGJcxgSj4u9
zmzcUAOFSaUtIIm2qH81CMAZ5Cd1Ceu3IPCz9NwSl3rjuTVCqIbZrXVwHhD4Xs46Cng/OhMm6tJq
wxuFYRrDz/MiSarJfJHde2T5q3D0IySKWG+w3i1hx7Xevv6a9Q3gQPeczIUILQ7dRNEfUOVzIPjW
BgR/9+EMQCLFFy222bPaKMR4NWWYvIHzvvX6t93G+/rQS/kUKVxZVOYi94aa2R71aevpZZPeB1Hh
upIN87w+T5eDqqtjgzdQyEd5u7nYhekjoIeo5x7ekfx+zrt7UevDyZeWB8ZIdLQ9KMyldkEGONzQ
lIWpKyb2R+6/2T3bwT6s3nNeOIf71m2m9hAu/RFgZWhde0TSHg04+fDPb2Y6fNBLVWoXwuJBdSFz
3EnaGd2pciI7ztIBb8LIsyAkzbN/hPS01/PwPUV/UwyKTivKrAvVOvGAVg6gqxo1+GH2joobOHTq
cu6pQg+3lky+rzcIL965X57wMFfuLM7pNiqTk0Hj6yaqQOT8XP6ehfLli0qJwE345RtRWUR/EPOa
ckfrehy0SFsc2h+bHgzVHRl7VdTW17bMPRFz5IbKa03uzNhi6VM6FVHtSml/TfdQfgg3u6scMdL/
DFpqfmi7vc6OdtLi5LhpBH/cN33rwR6qvVcb2GHNGpguEXkZKyG0Lev8/NvpURmXSnSHmeBRyUK9
JZEt8BJz37ZYRfOBzohqkj2pTEx9/uoIXaoN3ZpQBCM2Wh6p9LTDWYEtx/FBP1HijFrPb84qd8yl
BGXhOOF09u/75vSK1/qZqqu7ssuIb71+liF0Qwhogi16hZ3jlUSafFt2YitssD+51lGkjBTZRhqx
zVD0C/Q1uIcVZQFt89KzTJ6/wEQhs6Wu2lw6y9kC2KrDPmBjBRRNYufdwinz72CYFV6SGieowwDt
+84cVZ1t90LOdB3wAj34ZXWM3v8Y5FIvZaornBG9ygx/RtIgBWk8/jnVN2XHpObqLu3SnskWdhoN
oCdUHUfUI3km6bnHk3tTe4KV7t8CyLdUMqUDX+VdCvH1dnkKZ03U6/ZuIY4c+xKY3RpULRRIj22f
Ekp/G7j5phZz95OgmbTE+2AChyTx1C4wjdB8JslOyP2qsGicYKvr0fmcKUlzB/z2ZX/L7t7037pK
OwFu1qvhA6ZSCTQfrZbY7sExnX0lHDG/EOFdPtXYIibs5AyShTf3ZOUSM/m1l5ExTHUAujKv6FDx
sPNHz4rgpEiRllSpZVhGyZS0g8IFJKk8QjCnTJjG1FwbO6Qz/zhBSmswN1jS/je95z0/BtD3M6QN
/epxUXDJz5GqY8GZUItnxkutu6UVgCWXoTrp8fWY+1S8TNkaBF2auxR7suuF2oCpafBBEoPxPxfd
X3CiLyrnW7cI/nQ4vrCef1A6b4wmkcXBmB88QJMOHN4LbNAIe1+JCs6jLy7FV8wZ5JhUS4mToyFL
ZxNmeoROKPJGOWfMs2tuJ7bJOE9e8FWass6dVUyRig3vWT+jwDC1yKIQ2X6VIkfAH97PHlS3ZviU
g/V5WBSceAvqvOmMRjDb+OkKPsU7SfhKL3sxdM0quto2cqPzfZBVyDehtZLNmapttZIl8RXIlosC
xIKJvF2gzK1M/q3QvA6aB3UHMN/O4LcicsymHE9KK64pTbnFOGv4v6AbWW8diRHcVQzpcKKEiNuu
c7r3eshZhENDAiaUInLklqg1TPV4YkWGvMZa5qBgCjeqQZcGmhith4XZrG/JVXKhe6iQ6fn3wA0q
PUl+7sV5A76CwoSKHIsJZMyd4foX27w3/XUN0PDECrwqEjeLpLh884XxG3O7vvS2nqFH+VYqnJp6
yFg6KagifbLww0+iYnPfey+SY7oSLWikMzlBEja+Q8Zifbf+8fOU8t2Hko0/NJ+T+rG6ElmmhYvU
gy50R3+TYuwd/95ZLosWcpTsEuyOMF0BM8SUTH0APbdNy1OR3HUnlenzYirLeeDSxBw0ye40hJ5M
HZIAlzO5rJD3pBFcdCh1V1y/WGRW9AU81CHkGZ58u7uh2hNS3L6MbJjyJdWt3fuurDGfztrYPmC1
IJ7hbW8ZcSz/fAQXWNikNZI4AtZlzlGri6+XaLkUjiZCWA1KBbMpEVMy6t4AsKeXaqwwUG19Ud4D
eGtFnQnH6btk9O/fFVtAR5eoJ3WyfAwlBHW8zP0KWwXHFAj5UfbgMthBZS52GDKmVaaUDO+hYYO5
mgi6rHDq8xOSJy7Dcxq4uqdIWH6a92ytJHjon/Zi5meeQ6jdnBktvxjjd4XpxgZ47mxRxe6omD3+
f9VzX1LILpsP5Z77/+VZVvNKJ7gVImmUtL/f9/qILtYRqCnqAj9NdjSt82nWRcIO9tmb87sio80I
Y1xcLI46uj4tAjWwj/bFhNyzlsNS0dv0iRraGAA3upUXPKoFcKT/4ha3haUy9l2ulcR8oNHBpTlF
H2rLy8On1We0u79GHkY/UXdwpDe9epSvssUD4Lr99+jcIbdVfD4FurEyigTTp/cpKcWaJQCqcfLI
N43qzefLDdQLL+1cYkhuCsNEZ2hDJV9HytLR4T6Ky4+ylfqr7x2pHF+DB4UH33gG+KnZvY76LuIU
kIRAGB0q4xI+nrgH4EXBkEmx/eOq9577OPeiPx3sexGSptouTX3M+x2Ygd1bO7L+u9QPBjnAVzQv
DxxjxRTduDhH2IGkWU3eQ54FW6crQDqaBNgW70utNjhQ7WhcGO+7rdyjJpop5BlKOToH8odXVnVe
CzEXcHr6xSOJu0vMSfnML7kK098HrXQxwNt3/1iFaHVqswPj9/nYQHyWcvD8EH/N8HvLXi4bWnWW
I+QT/Ss7o8XC7kfau5O/Dh9IrSv0e1lKUDwqVK5PXxJXyhJJ4Z62o2prWqE+GA2AQuMDlQaMJlNE
1lAWU6O+cYySHGLEs5xsZJKlTR9/vw3zfAR6TFROCLAM501Sw2LE3m5ekwcgupu6NM3A5OiMCmBR
5ydfzU1+9TdSyczjEE9xc64Th0hpvWXKW/xXBAfwlieLzYVzcFcWV+Gwse7YjpEd8lxbUbVXXCxz
eHVvZFAeCklemiKxOGWzyLZ4qS0TUxo+wB/JEmGjPhEDGwd6zybTfR1/Mbj7IN00ODXTqCnXTI1T
CNkG6IOnNiPOcTYdHETLrS/zPBLWE75U9QZCSObP/ULl4np2BcUgEZaFsiuLgWfOxrMUEqb7v+tu
11ErGPGwLgnvBD5dMsTG2dKWsA6WHh4LQFOEAz4OBBgdFzwlirrdRr/P6dpHr8EPcMQbSWL+ZMPI
MBE1Wxvrhqrs/HnhIQ7jNKeiRJYsvDnwUe4ZwwsT47S7/hnac6jkhln+BrkN2p7umUw3BKB0/6RR
vHpXziwURj/H90++1v+Ir7FQX6X6atpsuajIi5e6+BS/YGa/dFuKGctYHAp5B6JAW+TI71NWbDwS
Gg3M2BzttyDIZEWxu2Ztasv7yz+hTlsff3AUzpj5AEJyROjVfGVpZylRDo7Yzwoo+B4yRuufgCnP
6hf+7le3L7KZqEYQ/5V3jSZw6YOCgv8Xt2FxC0ZYdH34xJbP6Wkjt7NRmXBjPOZYylaLIZWlfTL0
0NXZtpEE4dKwCD9Kc2cr+vx2/KNQ9rAUfROmdxh3OCgyfhEiasBU4ABgBjFTD/JJoLBgQLbIC3Be
IfR6/8vr7Tgwe6m04pbel9kmENrYtF7jXslJuMsRhT0wC/jpXJa/YwfGWnsO+lrJPwjm3qw8S2lf
TYS3bCibhH/RrhgZujVDIIFZqgSzMx6lCJnh1eN7AsyK+8L6fbRAsmjqQ0Ac4eUiCrEq9mdPm6no
GaQMMx6MN+s4SdFYgfW8Na6hdBVFivGXNQasKV96ZENTWgbXA8aYBEXaW4zmYLz/y8k4tMXOkGiu
07vt95dHHXeoGZTO2aaVoxdZc0kfUPyMfnMBYudCQYFoiWXn5ng0veR68g0oesmUeAFXqAzBUH2i
ZuLal8Qlyreik6In+fIFfWQGNI0iGHHAKjR/Y9gQAsfCmrrcaVzXbYi/yrNkP6vSlNUgA7sKIScO
QQqRVh47QufJYkC3jzee+nVxV/1+Ky2bgoULPkzEZnPs73trgHzgrGvj/V/yXt23W3tQX3h0Brf+
xesWUtd2PpSPIjcrpH1R7E6P4Xh3Xfp6T8jF15cw5vZ4SeYpRKlY6ksaNEh3nQsqWrakP0lJ/Hjj
nPBTNv2bMEp9sWusOPj2GDO4+oM55IrF/rkaIqPB64NviTX3QSfgfW00S/L0osQhP07uUcYiw5Bo
kAj0or33LhuCq0etdGY5kDCJF7xUghS2+Df7m7ok/iuFFt6Er/Y/uUVfu0n9Tr1vyO2QMUxtR4xd
OMXwzIEYsoSH+Srirs4exkjqeORtkqxwIVhleNvgPBgTwRQjtr1ILRWd3SmOYNw/rWmo1sCYtCUT
abdwyZf0Z8q06h93wf3Yu7m145Bk6Gmz43VLbqxJgq0gqSLh4wkn1dRR6qG9bI16Zl7dYRBIYmKc
iyAIpDofLh8tuWMlBFwyZY/is3dIIuY0V8+Qf4eGeqCmtxzD2GPHM3U1CdnHq085md3tbBItwY4y
w1YKHhE5H1GtgiWgscjTsr/Lj2oA08Vl9nkIVYF0BfBJaIZ8pDj55ijybY7GvqepnSPPUJ+ufFTI
pniWyTryeFoYjf3t3DI7V1IQLH39+ovKS3lfxdK2/9YALkL8GuczbAH00NUeq4cLPb/u3Upzy9m/
na6kLttF8fUjiodm1Yi5L+l+WwMkU91VJswYt0D6oxQcqaqZVDOXp+9hbVfeIl28au7igd+Nl+L+
wyW1EN4sxBdX47ojfk+4SPflU3dGMMVKflDcXtCis/zMmmPLXXczXCPfDg5e7K3/A7O1f8+zDnU/
8pB8r3wBdTPigYJ+I92gi7z+hUj50hPp2yiw8w2U1cyrRkBFGGxlMIIBuIDWyin8cxgfbQ/UYgGi
HvC4Y0lGDaxEW3B+cnVTBJqAW24ZZmH2sYadwNhi0y1756kYCzka+jv7oRZKUmd91GZXgkkFaJdq
A8TLqgNGrTECMhgO2qn3oh7OzR+3ozUWQ2iROpYXc0mHwlSBgjhiuhPzqmt2UrIBYohW/4Dkxq48
SXvwIunBQY1nC5HgCrE/bQrWKlDLzJyp0xk0f4t+/0cz0XExreYg63rOkBw78+fXs4l0I0Pi1+29
w35ioo/1vmSd5pZ3BqN6cc9WqBoD7zj2SBVuI5pMxESHp2bldOp4ZZ2iqf/o3ULThC8oeIGZAY92
AVNHEtrEkR5J6DIKXUIX6VESrJ9ZREZfeHBc/LUVAazaxcKQqsSvEt54NfmSzs0gfG9B5L3F+Zb0
Gi4p22dqWNfYSCnPM+4s7K2nyWcShYQQx4tjgBFg799buURhYbzjnGvWvMaLfYQVKt9DK3Vfur+1
rFpDkpdN+C5h3xbeQiWl795ZcmK5tUjff9nXDysctWn2/zIHwf2ovw5eH5ZV871aDpg9Hdfa6b3c
VdWpviMH5Z75OeKOvT5PM5Toe5QmUPlW1CVcTelFgitk+rufN83ga3DJIMXXwlyKIma3wKYGNtBF
zkYiOu6yjqv7O9uXt1VPGJ7bMMP6PT2s9OHRKC2Z6wjnYWb7RGLAy15LEaV4E2k3i1BZJNuvx9tF
UXz/TcwYufUwGVLAprn51efs0UCJnxtb6i1PGzTLyl8DJagcw9HOIPasI90dD8EG0pf8A6lswjTT
bpABwcUHw+NvG9ra/TwR3deMn/SZ9AdAfE8OiDPGN7C0fMob4RV/tJwmCrdQ0ZWSJICeBFDT3fbQ
A5Z1d/lBmteQztV2K/W5xLMO/QgCFOphWB3igfwlSoPbd5p8HtRNRpWerS0UT6Xt9t0XGEy9ATPn
4jOaHk0ZornEHkG9NRrZ/Yj+6bWhG9J+D4b5FssA/PBxoGLVNgp/ARH9MTbh+GgaXEeccK9i0m2B
hWliSZ8KwZs9vYBMUL74+UEbuPZfF0R9gocqYDwLHAJipvRJRzXdMmFDlp+9l2ZdXfLy6BMZKObG
8R4rJpcYBPp2b/asuXLNyAvnFIa44VfwHLRIqDe4kxQJvG4A/v2ChWimvWF9f1dRju/etRMb70OP
3KoAkXdEzxE4ByPIFrOqHqk0bw/BbMY6QprGOOyRuyeNBVZf2sNAqqyRsNYL+Tlr71m8mp/WjoWT
yn///+wTYzQRjCSN0hnTBk/XXsdOkrKZBXfJLtBB2fz5e5il9G8i4ukWvz8gXNRVo+bucyKUE1A8
tFZPXE0ZpQdF0i6UR8pEEcY9ja0djbB9VFqQoUKMT8tAjooOW4zXhiWqfTm+M5N65HORAEjU4IgD
CKjHASyDCEJcjNLbZHeudzDp4+9LVnnVAV2XGP0B0x7M9CLkPo/KkVBwNhCWXj3ANwHU6jmBL47q
iElMP15avsaAlfh+z+aMitSYXkrrHQ52xBmDmRcQ6WgNjounPdGm4gPyTob1wR6WVbjjnVVOZax3
nfBssI8eXIziONxE/MFYGqf+4q4E7T1AML3fqVuWT4GJZo2mQrytsocM9pKeBQWHegOhYkrSbHZn
GKgY9LkUHtPosl8rnwuVlJgpIHLeqJVkZoofpArJzi63JARsxxao41YZ5CpJmkBQJIfumouWpbmL
gcsW0UT3FM0CfSEEMiDMcyy0Omplm27O/+jycJeO5vjTaKPF4UQesyIJxgHrwl19DsdcI9E9EhIr
2oQsKHraRu5vGYUo/wilfWAN2eLnqYVkJ0k0jT6cqwdz2ZqIO+xrFWOYROmq45Fs+9JrxNcq9u1k
EvAMbNXbU+rln5m6sEg+2oDJbyAp4Aromo8wS3Ysp5+HgTD2cKDA02/yz9tj4RWeZAptAHK2CSFy
nMwkNBJnsYG0AP2V0OZR+2njWO5lbCxptkvHP7qcZ0GmPDuzOZiiKGsOhcuhKlpPjHU8pBsjCcpx
7twqDHZ6a8Z+Yk206FJVo7NSV40ESHha6M1E9Ufh42BJi4FPo2C/ZwHrik94rdDwxENJ4V5PrPMr
9XjC3BK5z307wMwGifvfvcnL0YAyipuVxGhKeTzgchQMzJSBZeG0YMzlWcpKF6lQdUNWQ+nzF+Ct
0sYOQafTHO6jkoaaqX8+ZG6e6aqvgJ1ACuX07VryV5qJMVOVJwV0fjbGV2U5EqTsrX0/6CquU//z
LChIqGtlPESdCvuw5f/9iyMpbqo5IRB1Ob99MA8klklFQNcm+zcNEvnYRZT2B1EEBY75/jvH6+cB
gNNBzdNQVrh5ZtkRLacMKdh9zTvqDCKPSWXTsGWWZ+2Dc/7dU/j/CxFcPiJyoEHOzWo1j7lYKIpt
vgkEOqUOt2DtjS1M6M+guUNdYIeIMUF3xoOS7XVXBdlH2wHp7sHHzlCinJRUwHPLD5i4VxkzTI5U
MA7XgqtUeGNF5vB9+tfmfluRvFuEKDNzu3iVlxBpuTyEhVEH0Bfynm1w8i/s4v9HPp29zhZ7NXj7
9RHrj7ZXG0kTcfqM967MH0KaNu9pCM+23yQQ1EjJOJfGY5PTJ8GLSAvEe4+BtJemyKjqH3svY3bP
HzzZcbagnEmfd14y2GwnkhfjKidO7lBxTsmLQ4C7aBWz+TgTcrXwCpmt0VBuQycsIx+6BzCXCQ1e
YdPzPWTEvMo0YV+843of6/SlfJtIE9I7Y6ZawouGqQZYEUpJ1RGmVhBVrnvYBgr62tRJI1mvNa+t
dwnBsFeecPxECgbM0mk2lWtg16Jkxky1H0NlTur2BJAq/ExSWmj6CFkaLBeg33R+pQ6K6slGnASk
GAF0B6cuc2An/uQ7w6l00n7wAiDPi7mDlQWPeeE/7Chm3ZH++SUwtQg59fkhAIIpE6nefVMjVxLV
ytuZBkHz+znaOZRh3umJbvQaOI4JYKBrMlzEbkcKXIX37SWq9fudFHNonWg2vTjZCOUvRiv8f1Kr
H8Um03S1SeJ6jslVO0mD7ChGcD8ECeR4XIt+ee1RY1+xnfvnsVzbGw5740yI9Ykkiccwk0LNo3CA
6vLlf9qwUZxlB08xyT+HUeftcPHnVzv/6gfeZolobAE1D+ZkZOmpZUC8RKioFNvXeyu4XqrYj7+4
RVEZ2SR/6xMSOQiul920JBfb2tvn8Bhun1MaJHbNtQIKBnHuzJDiOR64nWPIGUX3zn5lQfVrVQpN
Fe0n3ZRAydPK7CKDpdQiTfepPwY5ylHw8WbLszGujuhQIvnOPLZmzjBURSMAuevc+wtnafvJxeU1
eYnVas19URsOhYHg1YURa9U23wavPjGoYpIZovRS0bSTGp6q2O0iLH6WJ1vo4Z55wsgneHV9XFT2
iNBKwElncXOWMlZZbRDTscqXkUmhPjM/LRsopFWKEkoiRQ4LSm2BuGmZhn/BAoss5x0Pgh68olp3
AW313nxuCXQGMsA1lu1zslgMRVzpsM//pdh+JkLKwKlbFLFaeOs0CbiOpLioBGI76klDt7QOTcdj
PTBjuOA11zfbBhx0egckxrrntc4VEns2zJzGMo3wWENAuNIyPDg8/7Up50BS5o4LWuPQyQkmyfju
Eg2wLU8d5KW8+U2bDWEWk+LtekTvWmT2z0LA4QB4b1I49NfLiFTlAkJeR0WpojU0FN2Y3cJ1gAHy
TWt83w3VHikrTQutdgM0yGJH/gfdXHK8A3l3KY6Zr9zJnUlIYKZIPx3Jvm/lvRZz64cKH/lt9Hyh
72wLkd0DDBeJp64KpdMi7+vMSoNsZ946+aS4ERX4M/GBWctFcVW6XAjT4QQzaA8jLVytspZqO+CK
CiutFs3c/XF8JjHQC08VkJWsx2ycakspLuGDD3O5zSBP9zPOBjUipqgKNbPxb4A7Q+BPTeiPOxyw
mCn8pWcHBXGwHblQK2LPfK4wrex+ZVyZ1e23kLij5oO2clIihLTQZkoF6eUf8OqVxEQVrFXXvtaU
o8O4aABPB6PO5lBCvmTccvYmXEjp2tLuBmjKZZnteu/xb+y8s9+WmR87pM4ZkSQfYQPJGr4yLE1x
Mq5ochwG7yImgx6r1sLmwPixC4/pX7ZDifWVsiga4cx625davNUp4LYiSOQGCCV6yoJ8CLt5sp40
osZ4gaJyB+c7B3r3U3GYUoHnN5sHWFkQKv8BXn96VJlIs2hw6suW6PkDYduiP6IY8PvoalAGCppt
q9fbLuIDqb0gNKVdiv425hApFjaIbY7K8qQFLpj5Q3xITyDIDrh97Rrz/d85X58egPIBql1w0SxQ
ZTGBCfbjx92YuPdYrjU8cpjILa0ItiThvs7bzc65cdLTaqPX5HsOo5JQ1a0JoN4ltsnjGF+HAMLR
dWY0WxivGIDaZTpDED+oHunwlpU32zlCpB7ZyVGf8cIINhLgVI3elWZQNUk7Mg7WGdecT0ZOM9y9
/+84YyO5DCu9//u2fqTyyyjt7uPb21Q0w5+a+6KXkDELo+wZYQzvCXOgO+4kP3Vz4b7AWGGfcLPj
551r5rpZeDd3/ug3s5dZINwurfgyUZbAQnj+elvBWxqop4BSjvn5I0p3X3U7h+En115WFILixk6W
J945r1XtgRz1r3GgZkrfeQNZDbrHTQwmPUIjK7ZVNSPNOUDNr0Qt7473pZ8F8ZQ+xMQIh7R5AyOI
XDeNSv05qpDWohF+4GjXYKXxUITzVjWUcfq9pCq0xWLOMHCAqGCx5fQGsHKarxTFma6/pfrzj8mC
kYIDX5AicE5kqyt5WD299pXkPTveTMQDFenVxDqTrIICUnDAlKRBLd/jns0DQ3EVcTF7DLrrbpPK
K+n/MRVyjhv/tK4Cm5jVeks/yX22BxNNOZfVcbi+bN0AaRGlqpRwW9LoCDuk2ouvwTidUHVkX1ox
wgpr1pYkGti5IcsxFcEGeJPmPGFS+6G5TW9p4TTTDOebf9aXCZxSi+oUW48f6mi37ON7dPGNIoht
DUNqu9NM0KjIqlmO/2bU9Op0NdvB90dnReGqXrJY+SlKgK/n6r0Tx/yMaPqtSJkuRHnik6naEsdN
TeukhvO7ESoUHHP3MlbGR2+yR1aCMg6u7ROEHRLNxqtOJhFHAo5dcS+I9cKsnzwJDpCpAEDxKLti
Y4zXLeY3bsybm6FAaz9a4m8OAFiMuJzL7RuhPV/2CGY1SB6LIIGNx/K9vPn/h7mpB2Lv4CRF/xEi
/LTkiF5XHwmsG6f91VHACy71paPkEq/yW4sj/D3mFUrbNWauicpI5Y/7q9Gwzuropk4PX1+zWrqL
oemORKhxApdQZ9QF5hbFxt1YOusHifb8ZToZRuSuMUrwaZu14X/0po06BHCht7sL7J9u2wmiOxK3
zbP6EVpGAp4M9YwWkotzJjGBR54QKYn84j4Zd2MKOpfHlazgPrYtVUXJe9FZbe5XJpQ+xUCcyiLh
qifE+z7fj3Z/QThuycnSPgNm6qXyheUF1ROELHTw9s//uAyYLkvw14NK/12F5bMTnGV3bECJX/Lv
MqgJLciGi1Q/KvGmn0xl+CqYs9t9OWm2l31hgHfEujKB2Zpm8DU70MBqmFjloMH5XzMv0LrP+uKF
5gTekWtocp51msCe7mA1ItVWQF3C0fcTRnAJV2Q7UphV2+udjNqspRt94kc7V317kwlnzxYArLn4
CcaWN0q6K3zAaiVPyLU1eNAHKFmnURprmu9NiMrQewJ6vCCrVmEOLoxLpwslroppLpyEcKCGWcgL
1bqpUBoJHOuPzavCt7+hjLd4yhhcQgDxI2NOe4O3hhxtNvP57cWTxcaBHgorLo+oLyX8ZhGzCHUw
F9+wQTKnzmIOzcHjAp/RnynxpEqBQrk9s9PlXEuUW/MpzAl9DnfqFq1VOvW2Dtb3UiIfuVYVamk1
3+A6hx5c7qoionlf7IfIX4bpYcMzGkaJCITS9tNuw1f7kfl7ADalq9ib5vgaffvcFbzP6IRUrMNv
9t0XyJikWp9GzLTvgu237xkoXMyxCu6YCENJJ0i0d3UNfteTaNLEQix6tCm+uobAAH7gLYc0fQBm
mWKn4NLH/uKHlu/AEskhMqUdaNyt7Jiy+kZzYmMNz2secQk47pKgKcdzsTpVoTZ9pU8IG229oY1c
GTg2L6JZWcLujVjhNKUn6aimpdeYZAVhEUMqOOdYqzXBHWxSPPRtclgZGsMhpHwnDrjx9qdojaw9
sJF3FZWcWLCfCvH91ICEeNkGwC1vCj8UNFE1QCmsIyWBPxwVIInINdUAksjhJdk+X32SW4TQhkV3
kj9J6dSxbeDCJSvfaMXvZoMwj9eGHZtyYWyDd1rrZeRmKVZNIi+EOWEGm72lSAdoEwFITGp6lRFF
EIH2SOoUIejI3pM5tDVJhdM2s2RMk2GH3U97vk1YDlR4Mihr5g/f8RpFnHDPc+Mt4KplCmGGlxgm
9fkGitbH4rNM++2QF1WibLLlbitsHNM62f8/Qa6aYZn1kdAu/fcrWgdgmqrD22J3HS9eYKqPcSih
RPF7XZwKOTMK+r8c6r5+zNArAxqJYDgPXDlnP9MUoA4M3A9Uw0FGIaODVWklpa4EY+hpJzhaJs/2
YSFo+Px83rUImlJzQru/Z45sYAiL1yO1NN7OxRYCRQbOT91zKv3YOzs0fTkxTYOcp4HGQeagvrH+
uyYmzQmr+/mGJbMtLbQaOHF/Qk/+1FdU80VBj3mqMbk2rg2U0pZC6K6RR81YenQF+d/Q7zgg+9T0
VaMOV+9+U03J6/xkW28Ugh/x63JDN1oOqyyB1l9HxV1yTYlrUL47xafp6DQH0aVp9rg2UQPTRRtU
//o8QKKofp3Y/kbwb/NBz57OUrs/9wjbcvMmZGAFLuVqTu05oHXU7v0uKWBuFhBUaENiSBceCyf4
bMPEwco70Xdzsq1I1qobsBgCJWiN7MTe9o/wM+46ebYgl3HE7ABbfVdFm6OPVPsJ7kRb5kbGL2So
Wj+fjVf9jxKKuD1xyVxaFrDHNtOPHf4D3KntMTlO4AT7jQtzH4mgU7qaYZJj0fa5xmcqOKB7Y6SZ
nD05IcUbqxbIavP+IWHY2SeRxLMYNrbe+SGT9HEfSMKQHZevNROs/qBjyPogtkoy8Nbm/n8VCT+O
hwYvinU0SJy4dbO6WiwosCq0P3lbJyc5+VFQGspgKRhj/W6oRbnypOzuG1DHFCy94+Eizkpk3uhI
qA/HIK+z14SqS9Fks+2/5e52Z6MwkD5PL6ihoU5jAeXaUtV6LrRFjqcqT3FP2jjkdTp8VQ1f5Tqh
2rDC75xYvkiIp5SDdiEgbNEY9ozJiLBMdr0JhawarNufLNNTKmUkWacOSP5RtH7il94bPd1kyWiz
Ss/Tkb+KMeQEPkHvqUFTqZc8qsFv5bEIFmUv0pspoUGKlNAaBSgLGXpkI6KHocDTZC6/XFqeXduD
fG1LbMR1bRoCj1nOk5S55DMlKcFSrGej20wIkDBGoC7F5EXJCn/h4LsaXpfgMHFcsGaFosY282AZ
I5BeswKqAjs7TGF8cLkUrg8EMybykz34mRfGO9nXTbD1TCiAmkWDef44jfJjTxBs/OifP7w8e8p9
3NuF0DcJLYJE11xPxyedqrePZ/yRzVO8O4vAYUuFrEfJRMI6uVIVIjM/4rPoM/OO5vW1/xiKJ5k5
xonTKkdJiIUYIXFKNO0bKpc9ZC0X4MYa+ZtKJCV5K+96D5A5SaCES9l1ugTTmsaRPtxooBSa8+Bk
Nsn9j26fVRsrjbm7RRJLhiicI1qLREfkqIhk1oTWFLNjmPSL5vpUZ6QUP7IslHq4RNra6ukBGSOr
0cmhzfzsnGJh15QPFmo12qvKjQD9bYU5CEfBIGD2fZ4B80qg9PQ0zn8Txq1z+IFX17Fqs8d9BRVJ
FEy5/+Tiru5QaGdH6YdnkC8lEs9Jyd3nIlZJwTIhYH52+n0JoJSZmdJ0lCtp8w1Fb/n1lgHtopXi
0puznMf5JzGmHR9axhSfVvWbt3jhoAPTEpxm+p8ymCjj/2xvYLZnJ4wz2PgHCcuYOYvFlUM8AZjm
CrSCBUhkvldRdQrRlgCg3OmKvwPRj6e5LayoS+f2PTwEbGsvuy7bmxtLYj56t4FIatDlL3gPHgPJ
SIaYsoJIFygx++5+Kk0v5i51DwC7pXtJacpgYEJj/mB5QU1eIWiFHeGM4g0nRKFF+vSJ+QVbzinY
pmpXbdaGT39j2T9orEXkNi7uPWEg4JSygepX4G/f/9keTBreCh8IYkf3y7WpPUrpjFZ6Eg6xajZs
3jOyhGQNLV24zasNpdoiW56KkMdRkwc3BJMCRjZrqcoa6ab9dsulH4RnBNp2dvHauzRY/eJbXKhh
KdYrdEumrowWk5EKVaXruGNn9u1nF8FCyAuya86ZPPDpAdgmQIa8en/cj4IzQxofFLSCRSpa9B2w
ECHmUwnqHhr+Lyj8RRKXVzjmdU1MWhXG2EpEeKtOog1Hs+tBOZ3X+mH/OFilt64atfWL6EsZPfve
psBRVqArN0gqza/q6nrRil0krY2EjDMJqJUfahZ2ia+SsHdbgi74DwuACLtTmNOAHb1S3KaG569f
4eeG43vAwIazwLq2T8NikmirogLMVzfq/AuVMHC3ZJoVeDeraYwtOCGtACDR8muGdEP2+LRIX1tT
2eBZpHDcgMKxhMhmwuMN2XWO/lGkTnZ33HDoNMY3dR7jGqg6U5ULKEySKrs8dEVoUCEZuVm3ctc8
wQVr6gojVup3C6m1ILhumeh7eltIwre/5q93GACWE0lDFMtfLDUVd/G3zryMSfvGcY2qAnzSBaX+
i4pgJEnxEt6Es9AUldqXeEmiWz+Gmu8Kqk6BvxyThDrdOrnR+nLfLyaaIZIYcW+EvAyGXREhBc3b
0kTBwLUHL4bf0hG1VUlnf5o+xsZRf8/MRNkRW/pLE/yywCY7S9+bVXpJJgiSNkhTiGQxlxpslA5X
8FeXaREt8PuDuIJqywNcE31bKwS34uQhGbd/8v7ZBBVUnfbiYsL2V6JaQJB+g7Zj36GhtRqDiJ7C
7dV91z6lyMsJ+hF8bIEikCxDAtY/uGr7gRwrC3C9pCRivnR3TLy8pOkAHtrR2rPntUIcDbC1BR+3
b+JsVGNFoxqO9Nz34eLRUoPF40OXCKpN551YVqQtKJF2kvPfb+vYi41p5F8LB28kb7xbxfNKxOOm
9UP6KWkZ5kCE3VJCymdCe6idfmdqXFXZkAt1PMYfoRc63JrQxmh6wqZDkUND24xIafdBbzifURUQ
O+PkCIrBfDL28++RgrqbvMfOhZ2IRBJRzqFfhpZYS4BWZolt+BhIT9RtIt5J1PCrCtJKsrgMzuM4
3a0SOIH3AJ6XHpymV8FHdnHVY8vQqdJOthYu+Fi6+m+zEuDHLiRRVmPRxrKKoVt1ratNhg6FutbG
VecOA8/+1UNks4im1x81dylaR2i8XivBmYwwJoKWkx/rAzhx6EqKPYliIe0m0MRW+Pn/m0qKJBto
7sQym/q7idbv5PDbxgfOq2RC//CMFy40EC+xeDlDjlRFAf67obkAzX45Ue2KPvT9QuFbldYSuNKI
bj0CErpZNpL7M36AgGtvkVRZbs1fH4O7U1ncKxLd7vEj2Yom7a/li0USk2B9eYaCQuXc89IP1njH
G/oXRYcjthrjEnbyNPnPTFmlLcTKky2IxZZWaCNGr6HD6kPIo5XvEk1ypvS3i53zUI3k5roAnPha
marrwRV/4GIFfrYU0S5AQMPHLsL0TNZk7vufs7OuXdQzs9tvuvhDqhynd9izMHfbX3V5M3FL4YuZ
FugDcSA4yIXFW+6mOa0BKOK83+yAAi1ssruEMNFx3blO7uVkfmezgkk17cgZoiDbsFQ2u7FTgDOI
g0v35Z6L4wHXWLaaszmkWRGlsHFoIYtSift3arKL/nAJt4MRlG8mEh26Weoc4k2m6R+l06NXJEgA
PItUrLLA28mH09VBIiGgpkxo9xiLdCz8fnCnb0UfI0bXpQqWIb1FNkUjxwEMFkrTm11ptH+iwncy
/VdGTb+mkh8tPTqeaWXkTFauvW8gkh0oyQaIcs5TNttDeD5k7oT5i5JbDqh+wWC+dRPk5eBAhed1
X1SCXxh/25DFwCA8sobcNP/rNAWarjkCiT427Q5yxQRUY2U/5MCSN4SihcY3vHkoy6pu3uNAnOYb
E3K2ooEin+DPQ2zK3Q+KrFBBFUOUH2wfei8iTYTpZlQjFzXSLp+xKOBLWmuEcZdjr3fjASEVyEBj
H/jjzchlJc/+Tp4DQHLnLxVk9FE1egM41DGHgYYJ5Gn830utahpkCJDJphZ6VqIt8VCM7S+odAnV
DF8evHAhGoyFcgHbRQIZeIQ9iBefgQTk6o/Vf50QyUJ4gADhrRdB+86K1NrHcuoOZNWTPgt1Ypem
AeWGC7Xj/HMXWshamas9A8fx0eQKnbpG6YT4IPobkf4b1BjLFg7Vf80grQRtdLT6kmD8dwykS7eI
wzhoRbDyrCvq11H7Bcb7jIzxdINy25uwD1czsn/NM5zixVri6xBDYKibeMKhugPn7Q+5wWvL1OFx
06L0n5ZOVzWspcHY6tzXEv5YA0cV8ZWvroUNo9392ch4j24bKxXYxnF5UIYbiCvPFCOfXjjhrYnG
cDjpdXkxaL1deBCpwXek9sTtB/9rclGtqMPMwnOhTb9QVNOlrpr/bk5xqDc+E93ye9raXvLLlZhz
Yo4JqVAaXA8RLQOvShnRXa2FcXEks6UGAP/6YNHAyAD5GQrmK0ugG6A0QHvPudcr0BPlRJT0nZah
P3fvvbyG7BtGonf5cBhpy6KrTnqyLuS0wFZQUriQMvSZQEfBvVjiGKRCQGOShrp/g9qmc/tiaMfi
XU2K89JbXgrs+9F9B4nSBF3FBRtE3TKYF6khGiPcifxw0qI0UR0SzG821nsze3d0+zOYIQgsIbTr
q6JHsZD12Dfo2s6VSIwaWRCCZbzg/84+7ae1m4mP11AfsMWhzwmFv5eeGGNOljln1ppWVgSiEgcn
rJtNPv+LBm8q+pMVPlVVM5Kl4gsLh/lHarO2eTONwYkHmO4wKEq+F+RZbt5qC4zKLmbwF6Q/tkWj
o3dBktqcb0U3WVQJP3sjJOvfvLCb0wXT0+I3ArKfRTcN/7WT0bTpbmdQfVsKTo8snu48sVYzuhtm
wxN0YE6jLQwLj4oxtI5/TYlUC+8JaUEQSxE+j/AkBwHAfRvOPr4KdQcN+MDvhX/VxgnCH7bq77wd
RVkquzBJHf8gN0iFUweR8YuHDOuqWVnPtYmxnOgP6+3MPpNsdcKlq9sB26DlQYpYmqFgUR+c6KxH
pqETDT/fTzoI9qayRIMSkFzQ3+T62u0/hvJM1nhsKBceWDSQv+Eoc8d+VZj9vvEeswqJ6kSTXHJQ
b1yPzwgEdp0w2A3oDNgzpkzsB/TeebBocehszJLpr0QnFegCuTuCJ35qk5OVgVqHSWQA26vwSwRr
Kodj62f+kLP/3QlGq+4/AaDeWa1KB75pdfJ12AZykkABAsX0FFD+KEiF/2ReT3P7p7oqoXw/QL9Z
pnH68G/pv9NUwMuaBf7HJswaqiI1bb5dT2Tn3TqxU4CtWcunXNCg7esKOXAymfTNIpKDBa7P1Kmb
/IkiyPxRc08QJDK3YbejuSoRjc8RgrIzbBzSvWFyW/O1ht7VHAJjE63czxxX8fq28SDgETBqwUWW
qz+QbFZmN9KfpNsyWj06qmeRddvR3H+6KcU+vjJCokEtDR/1XIXVmE5wiI4KE/7NdEsPuO9bEF2p
zhx3iJEr7AMyJmMcJrKHS7w8IBB2dJJ88zOJF0CiIzVoKVeMt2p5HwTmhNEJUoSllyOhQ6KRS36q
IcV24vSmQaqp4jTXFhFx2R4zgE+BNzZ6NlApbrOAH9ulZLPhfFJG4lXEniXVwQ7WtWlFcI6Uebiu
KalEDfDKSg0/8psgZre3sqxXFWU+yXHLF0QLG+m3lT9wKD7+FirQqbnjvQrV05915Kdp/e56iPa0
9vPryGKlLE7cJn5CS8tQAaC4pmlXY1mZBXmmu6Q8o+aR18LMC19uMI/jZ6dRwq4QPMENYNqsxtQO
Gfr3a28iKsJcZhN/2WBTKFr/RacrIKdqY2YVufKtxsEburzqaKaUcFaKE3hiNppMWAVzhjXGf5Jr
tY8YVTbd+I78pSXZh7eUtZo/E82ksq3RtKkdskVJm/rkaMuHUrQdbSMSgJm0OUAF998uzLDxJpNJ
pHMuNp0/rRqZvdAZbpetPIn7BguJGxVw04/Lqmmgw7PcrgpSTnbAeWdVIFr8vv0zLvojHxpuTp3T
P9qBlxHqWJ+RDBVe1NB7JPEafQyVxrBpkZwm/Vbhu9Oo3pHnbvp8S/BeNpZ1G/HZsSKlcOl6aK9q
msepiKCxUaJWBKts3rWgvadg1E2ayzczCpmkmKF9w6eazkev1XlvRdDaioJeJVr7GI4b03lWp75J
NSLzP7RR3VeB7kht41WMqo7+x6LqJUAQigLnnBcgqsuNiuF9PATst/8HU4SuGaLE4FZvXBhYIS1W
vPsCRro4NUFRrc1CkEJaiQ+JfKx5VblOlQGCdpxWOzcZbgo2zOatzWluRYbz8ASoX44jr1LZSFuv
g1Q0RgCGESCNRZrKytTzBnjeWRMmEyrjn2hbw1/VxAgTH8Cr4mwP40mUeRXHOEgT5LHjqqqkRsBl
IB8GPcuqsvKINSOhBQr8TMQ94YGUUfvdu/wROJlye16w7Szh0/Iops6VOouJscboi9wUqNuV4Wl4
ACaQ37Ue3Lgp8rANq9K5C6Z6XFmcyXWduPMAJgKmqKUfdPb1tPRF6Tfg3hMEn4K9XmNNOwaS3q//
BQvn+KmWEBB8zv1Dy4KFO7C5VkJFlLuFpdUGUMiJ7PA8t0goLOPTCKi736krjdkSZvWKmD6Fz3aQ
e+tTUJCEDIwqrOC3kDd3KNVowntE9tI+LO7Q9kuUQx3J8sxYyrsX8Bk7yZE9JFR4SIHD26k3F/WV
hVu6hnQkBj0nqjI3gEhjbHHJLefoEOSytPuQSYh7N5AJJE40o0F9yFD57ufrv6dmRXOxfabfa5kh
7VK5DpRl73BlBioHuaKxv+qceUBM92OIf4zUl9wHpSWDgA1lpdmLROKgFbDat91YL8B4qE337Dw3
b7q/DoAQ1vW/ZDfskp9JY6JdFkKjSyPRP7amp+bD6ax5MsieIHQd8VrXNJQNnoQKPWUf68gM/+KX
CWGKKShgANcH2aZK9WowUblbNdH1c3cgZr6UdUAatZuPS4I91Y1EKj05q/OUIP6T+j/yCQL6v67j
FQ2xk5FuHYemk6B5j5Bqo0FP1ymb1K89Vyc8hzdg5EKS/IvqlCRj7GGMx0Cclzc9/YHyMJMbi6yG
oLdmong2qu9nD5Xt+P9+z4tJKhB3FUyJMIyCDduT/+UNbB0GdI5YF8azxmGas+CnWgdXfD4F/T6B
Fic4MZkFOlS9IxwLamg28MIKEvi5uUs56N/nWTlkFEWzHtk4yCdfnHCzEkxnM4dohHY23lz04pxi
lP9vOD+ddMjfKtBGkaw8Mmri5hgY8h8gFtLENbU7B3m3yhRvVvVcahT6IwZD0qc6YvzOX2g7wNiG
3HVAGGH/KypTySRcvLKj9BmKO4GFuvAUqnvlBrD6VJbeBakOa3qBUuxJRsuoEg4V7fV+5o2syUam
EGcM4y7o1Bx+DFN/lxc0n3YzBfHRjefCIIvaxfpUE/QMnyIzh1AzT+c6XCHoQCEY/zCCthtoh4HN
9jyW6ObMItSTxthS7QLu2FPXA6qaCezzN9fExO4SCMLv3iSIFNymF8i+uxwNFTV2OyEVEPFiyIVI
Ej/ygKqK1eS0pTTRJRxWe+IHSdJNbCYx2ArdTlncLk0p0DH7qRM3NdfJYFp+A4t1YZnbHaj4laCa
/jSzdoeBw6pRhF7hHwADrWN2z7LNpWgrBpMxwRTxTXqH+DTkkhpr5UsNN8YlDaegVd71BY352IP5
1TD8IPvFk7GD9xWGmksNtIeAmMaeWuNidUv9k5O6y836YvVUXTtWw8m7weCmL6fiodC/l7DljJO5
rjCZLOH9AajThPtAGlrNo4xxRfbJxNoVEZdD20uaxHOLHYwqSiO5ia3rdSutdBrmmC/dhzTnKW+p
Ixrf78ft/LqGP/3LEx3HNlAxLaMZq/WXFyfEseLL/BbvIC+ZmexGGA7dRQDejtDK7wVSl8MBS+on
S/tK7A9st3t7ZK8MtZSdYoTs9F/zuELWC1jZ30x/g6nRmTNW0b4962JQMfFU78ZGpAoIDHuOLV3I
FXaIpQwkEvxeIopc+pMG/4FIPM87WwzEU7eZkVNKqR656so6hXBxEsk7v6v/bYffdA9ynB2jqkZl
L9lnoRciSHirgYDIOnqwO8AWIBDHmvzV4F8hBzv/bfiA8ZmS5FoBLLvufotsb4y3LXexXamGZDDd
8rttFygt4bR6dhV/fmqulbIMBdjjMLjlgXG1lDwqZ8t8BwkAPLgL/7Bustu5BFUX2mtnZb9VvWuR
lchJTt3s/e2UapgGYWKWduYlmBMTc5AHHQwftqEvksUu9szI4UGIJmf0F6H2qJf9PYeRQHVM19Kf
biCpse6f/A++nFOCnWCHR2WMszNUNx7JfOwMlM8QucPArRvuGMvZIDS0s7R6JIWQUgNIGWsTLZgE
ZpPUxZn6nE+tPdYkhGmXAg8X8ZUuuO6KScdzeqwBMpuVZtYQoE0i3/MeM5rCDAGrFMnn7B44STUe
gE43D5n1fBiuj/31/mwTZ9cU0QReIAdOrpCeK/A343Q+d/oBgbg1Ei0g3fwQAKyzBNWqlbtjbJei
+ue0zJmvzq29Yni51tLlP9fran6JGjV1ni3Qx7lF/JTFlQClGWb8jj6AzRgQFLNNQ2Qext8q7XU4
Dj005PD1gUv0jz2lw92kB60yNGleoyd/5BhIWasILRsKSBDeN/1V8K4KP6TBb5SZxeqtbIDMOYBj
Aa+uOQQA2hP8gSreRZ4jqcsc/hU+isLgtnJUhS1xj8len+x7nDzorhA0tm162EEQfydSYFKg7lw3
I7l/avGmy4b681X0n/DcdaE7L5lmjD3t26Fs66plw9Itt3VTzxIzskRQAbaDO7+M6wgukhTBQxkj
yBj+XhFZzzKacsKXulElK+yp1vGBJmBp57lWUBwOabFewVdB8BQCLNXWBhE/6H/QmJ4irqeK1kAP
Y0AaLVhRoU3IRV9pEjFGkeMNprXAqZaBepc7JdOFun6e60NgnED3Xam6mZZlVfNMLxPUENg2OUu4
mjxeWAm2n9f6gvftN/2vNDNnevweXDL2QqEDOCNHn367ZgMGWeNnZXI/x0rsr4WB40KDPkzJt4kb
dCxx8RONiH8Ml5RMQokIkxk0D+yknzNIBvLgkbRC2VOBEIkZONmm9nDdJvQ9dWVMCcJVU5MLYp16
ypv83Za3amPx/Vta0PCVJl70W+y5ePr0MLOIOZ4SmlJS5kaC+D4tkS2U4iQzGASd8asqqxY9c3A5
gHCslaQubfaB07Orx6Hrl2CcpE3UqH15/WucGIeYV8FrZTVyCIr4uOpSioqn7apqiyow/kNTWv/7
9DkzS8Z/lWBEbfJD5+AOLYADiKsCJ9j6Q1yWMCgwM9Izh5PvLGllANBDPKPjj0dMj3jQjZcPyTO9
8ohUipRvzzrpPSTP1WK4BG5/W33NC0lycJwU7yn90ySXeAKlCFmAjTA1MQQ+8JA/267CqIpZxERA
MnbH3iE8tGOHMJ8b8NbII1OZq5j/ZA6e057Q5xXCH9yQY+EmW5ILJSeVoPyZZZX+IjptMX9rSrQT
xYG3t9NUkCUemM8/j8dpenUykvXUOWBgsVZVJIwypeqbq3BfhEkT0sZUdG0+Tu/ACpLr/7PpMPxO
TiHNbOSfZNPqOVaeXFt2i2ng0r+6xokgNEvPnJp2x696fZhajLdgpad5cMC45il+2zuhgF0VfO7O
hRA+ik7hHoV0Qp3mdcxnJVsrBufnJYCjr8+gpivRTgDXzt2pEpJEOPcn7/UlSuX67DCbRBjxOfRr
0+ZDCu1gZXaHqNQw9ZWj7mroi1RcYbUNb+MREDRw7lr76fm/0/NkxOypKbPe0TJuoDFzuCn0djHc
sEf7i7XWDqn2FLSpymNFxWqxFFSVbQb+Ah8fqYFGLsb5A2d1/Mqc1p8fbjJCKqmPrPikqYaVv2Ml
Z0SweXLCBUTPTCHBdDJGT23YZVwt7PWkMtXtHVyLFCDA/xpaJNpHwL7yty6a77wtTYO5NJUcH4U0
KeEeMFsc7ATnSXYZd6mE94wrOfdH6zRyDNN3u87ACf137Wdj7gBnS5N+RovPBn9e2BxzM0cqirFe
NlPc2NgzuPLpTn/2vug7LlUfp0wEov5hIgNFZ1D7RgEyjJPgBsqvXHgIup+fXShf7EJ3dO7AxBlr
zJmLTjVH9EcICJx8Rcp0L/ZI3pD4C3yoiM9BV04ooN4N2DTG3XwCKqCxiOyU1dvxMQyrvUbG5Mw9
M2HtNFjzxArEZt4MYBiNl516ZrAGadlHS2kwyCwPfi3t2x84+hBPw/f30zhOzCog7Q9x35alOh9c
m+E53rvjb1zWLclH2G3/jG9Yig0y3TeIxoPFQcd/9GRmcuvYgUkMUkvGjoC8bYUPUUtKuFZdTRcI
sno8DrXF3zTPL1WU//LzRjtV5xFgoq0/jlN2wnexRVvlwCEzxSLO5wZaqfUimIV2+wdJnBrT+HBv
B51ERIGNuloqtmA8uHw4RAdRr70TiAzqkgKuirwTMC70JYVLfLWjx2Xqmdd1WtdmQ+0E9aDguirO
p8gWZ2H8BebACfD8URwjeL4+Xd5OcNoMYy+M9/46Gt/KI/Rns+8518vZgDcfiXDKQgjvKNYAANGa
mMkK2i50HoHg91XjZ2A/CpQcDxATpaBZevFgU/3zN5fafUcFN8O+2gl4fwALjYOU8ad9Mn2DomcB
cg/dWmjBVYkQ+MNF69nbegLFdo8/otUHUdsJ6k/0olrgD4SFd5yvP81D9ngj38RC2rafZVBZcvv1
FPL6Hv391VEYM2KsQdJUb2xtXvmNqc8sWpnmis+Mky9kc1Q6gc6w8mIGeoDZcbk6gHr0HGewtEnz
LiDePuw4hCVwy4mFSqriWlNhIwvVzwDbvA4x2GSKaA/Edyuhb/PDDXV0f5YLtilvHMy8Du5pz5ac
hxcnO1EFYM4jtg109vltAYR5lPiz/jn675X3UW+06V5yfL7jfr3W4Fn1n9kenyIPeVDCkceBclCH
kDUEdwRr8ctMRocJh2Nr0fjPo/UFP+jA75zU3Si8dG0EFGb6D4izKD4iiThTEv0XhZtfd9cfG7Oz
ErUosR3xQ3vg6kQ7j6TQ0Ajl6gkyY8pZOglc8vpxUS2dELmAcxSMQF1eIJWs9w+1VJJWKBGxs8Qk
2+/J4vUUJ2Fimx12EYlnt44Oa9kQehTXTEFLw29t4NjDQHZFsKuaVFvbGgM7W1bwkMPYZUqW6CHc
yhGwdvXfWEKJBbdf7J9/nfqhi6WayR1Tt/VAd05reut/KRCcJQAJC0mdJaC4aKGu7U5k16+NRuOO
4TZgqKSrbw8nEGM8EEn3poXncUftaIeHH9uk8poszHxba3xRM7zxPirnEXTXB9vzM1f8STvH2MO1
o3wJQ0EjrnZaajbcTuNScyBPto8c+i80AH/064THcXqaX68sLnzh9Z+TZfiNlytak7ucLDmgWMdN
E4lAdelELWGh93faFk/kiXAqGh3eLnbpUcJ9Wno1gmeYyrUC8kjSj8oFDIz8B0++PlLBMeFI34mK
waBZ83K9KUpbI0zCZBuILb83Tat2HLQOjhrnZgnAhxn2GAaBXIozAIrMb/jrHgAo/hfG8dfys6pI
mzTAZUuUonI2SWwJFRnBDm0/ffbOVLk8hSMlzZzQ3mqPK/1Kw3QNyeCXoZStvrYudUu7CRjlxLrr
EOe3c/hH6DJUQ8EAmZxz2qYUl+gPQJNHE7nBE8yIlMjPPRasYcP76Lytg/xUzFyKkRX66u5jOVKF
37qAjE9kJd1yI6cZGJw3mEiyPtFO+xUFkMYXWMP7+xIYr/6dj3U3gS8KorAjcp8pkTxT+ZGxzDCx
GGUuChFs/eZu/8kffOZHtXfNuorjGB5lIKa75V/gvNPPYSBQfVBa1ABJgK5RXukEWAC3MEA7Hua5
Pj9IH2V6PMPlVKVVMaNeKdax4uBtTW5oEEjRnJpQtci73iqYgcQEqc49z9e3w7+p57Z1+X7Tgx56
Gc5e/8A5n+yWRP4W3t8oV1rZx2VtlUyT6JUYId+1QsX8TFo+m0LQtQxeElNX80Bk/S+x8b/lcRC3
QVbyTaSf5OlBjlSH1lzF0G4j3Wm+JyK5u8T1fYMYY/2GADv7tL6gy36GvhZnc7ClX716w1ySAuzw
00d/McdcVPPhgTWaAH+h/Nfu9iuj7tnAvoPZpt8WLMPDmiqfLBJVR4dQsIefO4aNye48//DEuh9e
UwWvXvxxJMa1aHi428QQ7iSQqHylEBC4xp0Pe1Qp1MhQBD2orCMiCuRD7Z+YONvp51a45pM5MXUV
zNEf+Ae6exppNgGSODtui773r3W13UZg1hXdyYkbxsIH/nWka9zJrr7699L7DtnLOaYwxAh916qj
RIyCtcJiYPM4tdHUFhYgM8uMnE5RSYyAW7iPv5+fR8E8pKisp8zXMOafI2m/yeOAGE47cfrVPYMQ
ZTEpbbQ5aHjzXb+5gkDIzii2ueJfIwvFGTCBQW0ybNx8YttjYO2NJcrwvGwqkWtJl0brMid/8t5a
0SrgHLP+C+Y7wShIAIeJtleA3KZJ1DykQwyS3WYeFbxV8uExgdnn+x3c8Sls9sb+W8qcEEvAzK2h
GWCPt12t1dtOgwxXm1iISP/5BSb+Qv76YfHBYh66KnrispAbFWE0Hg9o/SDh+3vEBus4IKBx3D9X
7YgDTuKqobEkDkJujRveHmedrsBwcimGTR7auI5iN4CG+GAZO8s4FunY536ukqisis3w1f6uA6vG
qu2NL1UmkDgbXGmKHK+zFMmKUH2ZNdYQaKthZ3E97iafuoK9HaNiYHyEShZQoiZ3BjgP7eKculiN
cVR7kVL+X0p6zRsd5rWjM+gmhpC7ClkHKikULeiu43aDBvEV9Ly++n1jCtZ1qO6HncdOQcoSpkNG
fIjZ9IXNP6FyZKR9w6E5JMFWHPISqHIObxhxJCGpRWSMmaeD/VExYGAHsWEof/1+Lr5QmN5Lh+Dh
oWM6tvwAxYIxoGDLsXrkNTNd2i/+yi4xNsiCMaJf+MW5g/p6HKfJ4j7/Kc1uVqWIdtJfIi6251lb
ErsXH1ZIHOv7j1otL0tSmqHNeDgxXuKmUpUD+YMbLC+3iWM45/n08TIwbmMskyztWOhwGgQ8qFAX
ca17ifUN3nr9S/tbRI2zjDfuY2f1kDSJ0/9irg/HoRhxtkkte51g0tZbfYWeKxvuROe7OqNsh7Cm
6TRwnWbcin3v3+QukunSxTkiKdPQEqKGPFUWfS91ej9PwAu4n09O2nMDqlwxjBcLoTLiinEyz1ER
/jepELzxrKS+ZPvFfGsQAoWYtE+MWkqsTOBaDKqbm2WZEntSkGNy+ZHQrvrF/UVzGMQApMo/axOO
6bJTa0hTodqD5xEdtyofWQiOOC4E35RA4FhlDipV82xDC5+6gFqh+Ndsx8siGKW1Mg3RBT420Ia8
Chb+mh5mOXbgkwo2j8NTs2CbubPPxDubKojojeksiTL5NGuJqAG8OLKT7N2H2oSxV14Ob1IbovCi
3zNEzKOEscQ4Gl5EO6nMZ/lUB3eAeSnp4RbZPqFEsvTWBKPRq6EjkMvuKtwyWbnSUquUi2x/HCIJ
a3vBRp8ylMBILeE6+knCMSsMR+xtXWOS/uJ0IVBFt+ajt7X5RMnmrVnAzamOH9kx2xTeHJ/bfVSN
VOzkn5MbaJ4MF1/ULzEEXq6xrOSf0D7zjZyvvTwso8oKmvNqwqI6DOvO5ANzhUxt8TwIgUqr9O84
zEnrIelw9YgAAV0M72zsnk2Cy/JXR25UC4kUUz9L0eck7K/IYMcRydhMyo6r8tt/jKyMlT0G7hqq
bozdr5wfItLHvMXodnf/5nKEMT2l7aw4BJfX6g/xTHECFz+KFNLFmy1wKLQ+cgW9YyYiXsc5HmNd
sgcetev0laS1F9m1rqTuYtldBDVZN0e2qz/9OObQmLhOrR19HvdvBcKQR/J9rcKdfqfIvlvBOTzR
v8KmH69+3hrWB3WDZSjjd+vS1j0+ERqhJ9f/npgKqYeZIIS8J/0oz1ahaww9GV44MLyFX6Yd3VFY
Na+Ttq4M/Zt1tS13BgHUxCQKot+KKZW7146SVsRLuwo1/tJrAnJV4WweQxsK4tXwZqmPc54kkFrn
cCIgkJzVtHY9WouBg77Ap40QEzC3gfDj9TWZHPcI5SDOTXM0kWyQNK5lQeQ70TEj0J6/jAyk9Glb
9hat888BV8yGfyMs+8tku6OTAWc2H74eiTk8ghKrXsP5WhaV2n3hgzxRyrtMCUz+KeAmtl+Le6nr
4hGpT0ZOhrsetwa6RhKHdjOP5ZMVwKoNdde4IPxs3cYA1qgZxmDMdlUbTzzIKN7ZlEWTR5lyZT/+
8r8r20QnIgu86P9zkuXzJTtJWTOfLSvmNYJlj71TZJQkwNT2OG7y6NkFb62vbwmsJ/bRgcSVUhxr
BZ8GiaiO9HPm3LU7rVM5x4lUCdWPWAD29d+UkdLHXScihsHWExsKfT5oLeZkfY1cgI06oVQb3vXN
rPS5CydAjhoXhmC1jUZRVhwYJKPCQURPu9vjMHVFoSQ6LbGLJgYdI3EdxAgIIM43us86IHkNklcP
fRubk1/9+haYHpfMAQjDcLDTeOAwDDHsnhBB9jBLxiIM2RXdjuQtDWZl+Mu1zSQKD6Tr6jyFYL9u
alkhQbUzmTT86umhYSiFFmlQLbrittuKPGmnZGzNkk1fLw2DHdrO0NehLjiLgNK9AsP2FW4RmhTR
o96YnzEAiD38KEymRiYXDcqoc1hT7M+9LYAaoo5loAZdTRRoWTWLEnLwSZxC6Ttv/b5HcwzEtT5d
vRdNRgLOMD0yovJ1aKAVrN3BSCU/nBST0FWkLgasEgd4K6Vwv7sheKhQrrESfaqorSZJXbt+htrL
umUUu2gpmHdO/7/GBuipdkAetRkGa+FY8povXaKlqaPjDl7vXPx4tBrSfccz/D+N+8X9o/20OBDQ
BBMxx1sFfSccmmKKJuw0Nmu2k/edu8t4rkISX040BaY8pmDDX6pC/uDqSq+1qE7IkAcj02LVlXax
tWEo7VRrfPhOwdeY16L92VAzWbHpBaiPm66Gc/WrUlos+PGeNcC7StR/7KaPNNkkcjxgSRhPo1eT
dH198BamiGGMI+ygFy2RXUQe6gQCeUshcCf89+bCBzSwDF5SZxlCeB1l+CC79+pwgw8MIfDrW9Nz
Krf8UflfQuK5lGVSJ+p6HeFeb3Mvu7lodYOHKDqpbJSGuuZZjilXl4Sx1JLT46wyEwLpif4pQOCi
RFIoXmD1ZjeA/AUUuZnAkj6dg8tJ+LiwXIf7kThCkogGip+m4GRO1JnTmvUddIgNQNzxFfsehdWG
2ZsBPAb7kGLct2slGMqy4AQhf9TulxgneapxXrN1EI66kCd/tmczoLBHgBXFmiF4jYb9j8Oz84dk
E+v3hVWUHbMvVH4bkv+6SpY7RN5+TKxP5FnpppnuOVMAmdCp4sW/4VZxoF65f4nF6yoVHU45jImo
V7vYNrH5rVStwtiZecTtPSBHGwwHNr4ZtkgkOD8yOwxviCUVzzySzOkDGYwpAev3FiKCvB1EYssk
iCXRuphJdlAV4g1Vt2z8gw/3d3jkptCVFtXTMD7AwCFElaFmayHwFHQkKE06cEoNk1WxkgpW68T7
hG4JQNrVgTGMcTpV2lVZ2hGtAleGtIsV3o0j7205uLyVoJqtChRztnohc5i/l1yDYgIMP6/6jfAW
2Qe6okUt3N3YVF/SJ5bicDYuUxyH73Ko2LKy0NfTczodpSVPbQdfAKymcQLxE2nUjsz9Mm5qep7U
oI9pyicPo+289qKosZrbp/QDsl5qYJh/R1a1FwZut8Ae1e+miTBgrQmUSFpq5KS7w0eMaYHTxT0y
ctXPNA+a6l1UwfPYajMZc6LzTNyqjfzK+o/+ENsu81DHSjBGMHVghP3eXVtyAD5B8zmNrDJumXXA
qgZNzJr3nmw03df6zqhahyPIvzV7V+u6Mz5SHVDKtxX4pZ+J7Q5f0DvWLKIOkMc8f7xn/f0NHSDL
FOevJCc9avPOMauStLaGyJ2j1kF/8PVCcl7qM9WOdsJLBTlkW/uWyhtL1h4RWRT6Cbbg0kr0GyOM
P/T6+4HAzk1dGniAd3lprUt2Tg+gXabQisoJBSSThWPuiKomqFdNifqYVN8orGxOsQ+fRi7Ex4tu
LeGCyvvLN3h7nVwxcY1Wjnf+ML2qj2eEuW/KDmGj3N1tuCCmUe+Y5rPjOti2oHW9PeOaPm2HoYn9
iy56lrYcOuJH8fktSMPCMmy94KORYYqYZYxujDI2XG89iij/W6J6Z+/v5WLxxdP3vxP2AkzevLOA
PtVKlXuyEzap+fGqjPoZot2Ylbg/wbQsmoJ3v7od2yyZ0FsB/ruCGoubccYp7SnMNKPdcBz9emWe
o9+5NnxW+fG+G5zgCe+H27c43DqyC9Y1uD5J9d1V0wyLe7ptero1oznLxlihHjI6bA1bevGac0TN
5RgHOVyUKSMEZ/Np2Z0MGF1dMro0YYTU9zlJvRbBjwEGSOFNCVCEFXyMmBhbuKkafUcFJdc4kB8O
+wGOEJn/qBxHxkuvjIRDz+3H+efBqB4Xp6G83FU4vSquoFOOtEajdRxkDB8t3igMjvG17JjgroQ0
MiqIZ8yrDW7//VFmnVc2qsNyTaWDZWmeBji1339gNYgPn+bebpeZyDUVFw5WnwzSNk7iGdQLxZaZ
XyJw9UK8IMsNIIvRf9p4LpL5ao79hJnIOkgaXRig1lxDbBYIQRzbhwmYQlfE6q0ZvxTqebvV99zR
9b1MZwpQ2npl6Ibp+AmTU16nnAV/GL/iMmOaMJ1OxBIwhKk0/3gY6oMkFsLwmI46urr/QxJ3oEcv
Q1F/NkumIA9o4RWy2TVFOmgAseQKtwoj0IUaMlNDuqw92ql6UKTala2V4pJ6ZCcC9GY/ekOqZ5lT
qun4XP0AkCZORQzaHrylzmHLMXTbyiExNJclQZ2Ua2fIUTHTAdsCoPKkaeIvPrLjzLq6nyZ6xJJy
2hEAHCWhQNgQiTBN1ygMaXK+2nxrUplSb8hO6tGmALuwAq2oap8iJhEKRusywA5/lBVKq0hDCgdi
OYezgsnpY2dV3WSrUKXKy2z3SoMOMRq1AHQ7BXT42ZNvSQ+k1hZTTeADl027lhIwudLiPfTWXcZY
qZs4Sv1Jr33TTB8cdoqvLKHJDUXsVCvpo6diYjHY0U7yoFPk81RQBu3eejrMDHU188535HIxSD5Q
/VpXgPmeCHmwiBt/gGyzCJ4nRqyU/e3+hxuKUMEhQKD6qEMud6VBANzUVKBtr6y5U/OyVWY3dMr9
1pLPSFaz9aRTR//yXcYsjFoHvDXdQPqstw6BSd7bMz8uJlVBfkGbDg6W0u6QOM1auig8NlADLGgF
Z2M+cdIaRPSWRp1G3gBcSwDs1TcqPnhAQnlmeGWqC4f841j/mh7mCqtGrLyYh3ILIHJZHWryRfXM
/YBw7RtvhWmTcZ4vNzjxMJ10op2+kSNwI7lCW9DthefQ7gilSwLxOAClvHxHw8uPLUgpwCcW1R2y
WCnJ/jF/el16fFpi8fxNhXwCj78+j9ysCV/+S7ghNp6lYTtB8NaCTE77+ybVGfScJokWhsgUBz77
Uln1os04gfuZZvm0w/O4wV6n7KNDJ6YcoyOqD3PvhUiIaUNU2J5YE2v8YYrNOAcrd+CwtHvHWLgZ
jKlkpRR8inqwBh6gpAZaitJld7+ywkLT9oha1pPKjAD+BijMKTnGs+BW8ZgaJ6tyA9DSnmtQ46pU
fL900OZAI8TcvL7tA0YzE7M+hRU2TvqXZHojTHX/BXYMUrqHugTE/RXEGFrjoi6fs9HXjZLaFut5
OI+AAZi1JCANv8LpVf4tj2PMK2Ci2f5Xb+ZfnTHpnhfAspo7U/p2FMB0thBh3wV/nCeWQsAfUeXG
5j5uYTbOcBpvwRY0fPz1xSBq+RFA0UcnPtxHbbstypU6cvFaYDxHAVz+fHGNOaEqhp+3C1uR3dao
pQjyvynuYPMSgwTbZBGMnLyC77Bffut0tu81XHRnNh7P/QIMuBsdgZm6EWl7ZmGcRJkA95ho1rnv
WA2Cr+dZqbU6ZKennm85lRi7Z8mR7f3qgspbklMNtzR8fJJR5lh34xu/4Rm8Bd8MaX6bUIPvmQ4T
BX9j/lveiZfRZVdxiHwteSxR6bR46fr/HPT80FNr6YlFveLfbKZIYDbImO6Z5GdMG4VOpgze5+Ez
ZbpLIH1IIda7UxHj2DAqq38PZHlEI7MrWUG9N2IWafd384yR1z8ULU1dGwpv6wDEi96pPSmR5L0r
1fC04NhxlCt+RrOgwawMRplu1WFthw9VlDWIByDXRl5+ucWsmyoxSLtVXLpXK6vpqHYxSFAPiL4t
nZhWkXTnxQkAb3Gkcp2heDdRQ/z/bq7CLkGEsUpxQl5NXdrfHJnQ6mpHxgv2v/bzYVW94BMQOnTR
EgioGYqWWh2ovTC5UQnrQobwV1RgRgeZWFDl6HiVTKGpNWhR7nHNWp0rYVIHd1p4nCx7kklu8RJj
bp7rQSHLLS6ZYNx5P+84P7LCMR698YoizUYUusFvp8WBRIDF2oE9VaFQmM73koi6lYwAbRXZ8zYc
qm93n3pwd3aX1coXn4IfA9nN1me/VBckU65FrJKdu5t1can1NjR7+rXYjNJNUI1wI3cYdKmU3ft4
cNDL3DLRRR7iHbCl660M+JChe/kjUcrJQKE1gErrcOqc10jaDZgy0Bt/yjYCNlL7ejuwuRPNfZs4
c3JDS8g2lXgvVc/bRInJrSvqhHidUAREUPz9AKeAuOwjQxjOarinb+aqXGPPepIRwbJQ4f6wMICb
4/AMG54XxtSphrDcBM0FgniVzCJkLZ2dEBu3NsilDVXTU7v6mc0Rvo1hrSwjf3ifld6m9NuUfZPc
zImoQS8cvJgXBXOgrdhqQAYgRf8phX34rfcB2MM22n+ophgFeJOngthxlnepDL3vqSxVWSWpvYb5
lawq46icOm4aOmREy1g9gQxupoQUIC4i70sAgIyDz7hDIrCpqmybDWjvEprpnHVpklJcrvgkyLA7
vT4F0hNfJY8ND8aV7wm/4MKZtduIl8pvR2qOOhnrzSrnXUNYcDNkxry+oCUgwEHsL7HaDM2b8uwK
TA2wWU6VrplLlXJsMCAbKlmR1XXJiuv2T/oUJC0hDx30mIkxsCwJKYX46TrqyPYykCQ4niOQVyH5
24V4bbb9ahBY6vPlKLqTLTTz3SB8xAni+nK0AdWMLwxmOfhAXIHU3cJ/RKGICxpMSaQme8ROfwZi
As5lNJOF6ti4M2ZuATthqGTI4A+c9VySJnlH2tkzE5uDnsWbBqtHvynMxqCqSRWbJ7n0g7+fmZfT
/o5YC16XOqeivnZToDQzGMEiNV500zeRL5vd0LHyy4haQvOZV8ld19H31acNJH6LpujicCd7BLYf
UgWZ2Pj0JmLkaoSf/Zsm2YG8ulaOzjbTa/vi1Ywy2v4xs7P8kQ2tmpjVAuyHRgU2JK1t2HFfD1oW
BwWsqNXbC3lHN5+wwvIuuyJlpFkCwjRuQpoByuvJxKPkpNcxeDHtQxUOiIpn+xAZRm4g/jm0u3YV
H1P8UOLYyU4EIYKLSinZUwkDjBqV15WpxyxZPW6JuAM9F60wWkllAZw3Z9oy6VskUb+zk597y6Gl
CQU/za9ew8ih9sGC/gOxEf7i96Q0F8/XIIjoXMdO+NcdAy6/Ty9E7z8NPez9cDFLsRaE8yp8YiCx
KOfXlmCTyyw6QRiN1VoopcQdXO/FexXN8fnStc1Q8ltboMCHKS/zujhdzcO04x5MhCuDWMaHENzM
WXzWy/9VeGsgALLbj5PDc9US/nGPQFCjNC5qFpU7CRcuXsjO0bciw4Xj4DpBQAavpY8YFPv7KxXu
o+vfyAsh8P2h1eIruajkfRz3didgxzfVm01megE27ZnXqg3PNri4pqlxykG8QTuaxyDJ7lCBwrLr
cIM8NimTN4ipaohzJIIZNe+KXSMYl4w5FtQl1ZniktsbhFt2hdXaN5LdAGHNJWgyLEmo7AH8t1Xw
JjeEM6W3IBe2pIdo6InhS0CjUEQR1ns919R5TJxekyPZhPY/k7FFydgBqnzUKL3NlSS5GcQlA/gU
v1En2XPfFxd9IQEqOsHBs7Pu7dPkkPKkBrrBGQvcZ+CUBA9l1Jw/oSbcgYRRe+MDE9Vc6Uraeta8
f3upm5F0cGaTOc52DoBmoaODTMH6yYujegRRP+axjZi8Socxp8sADsiKjkPUDJHeZjpc6ROzx61U
hhSYGbpaWHqPOoS6kUKOCqxQxW7dG5xzOB0gkb4J0CmSgIOulcFcAdD0bN4q8nX10RvHdcbVIm/p
Kjorbxe6GonrcD0KcIbtRIWiMbs5RGKJ/f/d6ejT6TTATQCw9Mr87BdHU/mrDvy7HefgyF0LEnHs
1Pi6SgfrtcCc/TDiGkmz7PSbENjtuD/UzPqPuPqUMo/kmH1b14sfAvnec7xS/z8IFrDjFoBo9e5G
syKt0twne9RKrV5NyWCPru/bQxiAcFp17q4p321eCzjN0O4rVnDLGOFNPYxAx7p5qkDX45H6JUQ6
K7ta2UPuIESSurUoCwMDWCTQgYXLjpsSHyU+ECqfeuttfQsN1wWpEBj8A3jIP6ia/PSBtZPKqdYy
4yaRbBmSDGPD6jE4avBNOCx7Z/zuWn+mUh/oLAcb8lId7VXqHY27X9/nbZSd3ZnmnZCreOoxM96G
PTnAHZV2mTz4XzTjI8SuMrYjQe/hjHgIiIPINd7KOcdbHSKCae0AlL7AXpv4PuemmfBZT+y8Gcew
cb3K6uV6QYNoEnAQ4nopGvT9d2nuTyTR1tNoeHVv4CkklGojjL+Akb0eVml3YaqWueMfX6CkPFNK
K1kz9tdJlJPf3IzJWB9NNtg/R/elRzAKocY7S1G10tSTduL6G6ETwBhHQhWj0Kq5d00ueuvD3aQr
QAu/rPGoVdHcU5ZF3CYM9/1Ak/rjGSXyLIdLpscKm6044GcY6HLsdi0zGHvhLE5FbgJ8qY6JCSTW
d235U2n/x73uxWEgP0Z0up8+2l4Z3DLOmMi7eApyziEXWBKAZ8CXwWa10/Iz123xuq55+9WNJm8V
4e7dQ6/3mOZleA5NPtJi6aSPUzSkG+SmpakMeaw1LHQoAc6HQZEwYrQrVVO1TubALHTHs2eWeF3F
AdPunhWndRZeDxsi7GK35D6K1PY34wKTYlHPCFvAr3TzF1RsenAzlmFQ/+n0KeoCrIPiLYwZGqpx
bBtLSTY4AvmtpDNRQ6RnKk1n2H/DyjBUfDvZnwVRNOxiE25SrvfFmKWf+urtl3AXvNKwv/ki+qUA
cVowLMU0zB1m1NRB+bflkYg9zXuzCg5QCoRF+WixYr62/AOkrdVXeVSk+wF/jquWZvpjAjRXGY+M
fz7QxzdCkWfvY6KhMNUuWlTUVJ5GKoJ972zzPoSI8IOAFoqApjCGR0JnK8NhDMPcc27ni0coSj0+
dxV0KtOuFBYsP4yS8/cxdyWrnafLr8D8fhy/KxECmN0E2GkAk4/hAlSBpxWbh+oVH0/KV9MRU0OU
TZkgiX6l/fxPGEP+9JmK3Rcjqyw5QY9UlJmWq21++bJhUrk/tJnSJp0VoczZXUd6ZXouSwOzfMgC
Zm+fDwwH4SMZqxkJ0M/5qUpjBPQXUjbpgb7Lcs9H1kZAXWjK5fThpCSziAbxypJomeG9CYo0TJc9
gj1D/NXCROUEx2OtY9UY1i8oqBDlHX1lyPRUkvx1Hfk/FdjW5zJfDU5DgM7v2QFo0LUtMR8O2dhB
FgsKAns5rMDac1uK2Bc8mzS1ULzusXAwcrrSjlQ9mKZbPxB+rggwjo5oQhiLYvGf5uxR7Cagv0ia
kOQQTOXqHsZukeEGNx7GpVHNoxhEvyyBfXkVWudk3FjIHdxuAEf/+kY1mlm/MBIy9Z1hqRW3c9Ju
/q58VRioKPcOODaZJaJYkpxGOzZOKv1pktJgcu9u+cTdaG99R44w6q1NKaUr4OhVpGyfcGxcTW/I
KnSpBM2WnGddn8Iv8bPPRks2M+u+oZj5PPeTL3t6E0Cpbat9kqx3iCQHFqAs5vCTOFszF+o5Ks4j
A4kNg0MMAd5cvCp8pvJAGOxwR20BWfc3laivXonbHEnJbQ1NgBG5J7/TO2nuUoQY7S/yLP6vkJ11
ESIufLozJnDRhjpbNLu0/l4Iy9R/kQJlUyCUwzrkTI3reprD9oeamD/Oo1I7TWzl7Lq8tT8f5nCD
gOA4UlyL8h4ulizLmdVKysrB6bi+XTUuawtpCdXUvk6AuV1q9niNx3KcHtBNn2LD8+LyG+CJayU2
aAyCHl9R1nZ6KzM05ILioVyaP5HtioDcWOKmcpvEMjAtPVAioABE2FMUl2EJ8t1JkhBv76+LGPNy
w2jiEmQ6Scy4CNjXmLy/4sRzR/DZEKomDm8JmY5D5GqqZNmi91MlvWd7kIVhWi8UA7invC3vkgv+
1+fbwa47wK59EE5tuzwYmAYzdqF1zo+5/X4bX5zCqx188G21e2JdlYA5WlnJfS7T1v0iDWDTlVGg
jUIJoJYcOK83DnvAg9ANpeitx8zL+NCsF+dlrqEdu1uuxYgHzewlfYTmYDO+53iHgVxo0X8+yjQe
OMaTAv4yax2G6FS5ycyo88EplWOgIB4wiJ8G0I5QeRvRfDUgyGGXe7Mlfpn8A8uFMUiiDwi84137
KjBPnQbk0eYy+a482yu0xN+WruQTJ8wy2YRXNFpYJhb6G4DJHlZblDKh/EKgWvdr7Gf6de9Ve6m2
baCqQxjYigyA+yMLcf5+NjGAZUKjlMUOgQ2diEgpaGXP/uV//GGEx9nWedcUUvuRagiriXliwYBs
5xb6w5695dKy8cKuzSyUkpASxqFynSD+Ywslk4tHpwwjSMe3rGnO6+6KHJgO16Cy4tx9Or1ODpUq
UInwwoMsPkl/EiIqvRwYp0pQY3VVesBQTomodrmXjC3VsIvvrmPhoOw9T7AGsV2XpaX2coC0TJxW
AFNP11Pxl6K8dKtkkHxvRZuuVcZAGkmVwCA+GW5z0jTknRLM5Coh6yWYIan6kBQNvr3dfvCMS2Vr
ammKxA7Pb3jmo+Qpjt8Ie/5RUgSkeMEc77jP2SOP2LCEjj9nc9lX6IopNsg6lIBPdgwwFZhvM3Xg
fcGaZZw1p9SMHp9Y+26ivYDdfK8ijUg7sHzqRVRTDNJzwG4qaPXMJgKtTZye7HCL75Xsl7Rznr4b
7WnVJZpaJqgHfpFNjr1GO6UbD1JzM4N+axWeI4yFC5Xv3GOXgJcD3pgixyeUz3l1B5Ms0cto4U6N
JrSAxh/TGlwajdhkssvhE15VUNQYrQTSemTfSqbnxmHyalQtUb9D/gESUoAPGuDSnsLbey4iyZaO
vXcgRt+L21ct9Xt+OgQl8LtXIFLnOa3VXF+3hPdVcQoBm+2mVOpFg9V3/Le0bvadVK4BDh2cjcAI
FQAHVH1fXRmtPZHFpgZtQhEqi3QU2msLqt7NOwjGKt05zpOAscHbma4qSF+AF7VUbz0MQ71QT7aK
NeEay+hW1GMjJxA4k8ZaxB7X0xp8OmrGD1HtDG7BuZSsoQ85YsjM7st74f+5tQhxS3awfnYk8mkh
nfQI9aAleQsYI40PhP8y91uZU9bGVq50+Z/bpJr5+aTh7km82gxO5jbJuaMUJhnLWsvbJWTEM0pL
9kWOCZAEjxGzk4FZ2qOMQfvFlt33DzVx37VsUBtJRDLpauajkqtzeCkwQr4T28cpx+v+WtO9nd1q
ZnYLX3lI/xGjNzy5Obc9AIDXfDdn57fimiyMKJSvtWy4gjC06CZacLI0WNFwzBWaOVtqPq6PPw8R
zAs5jfFH1e3POLkwzaDjFj99FUQT/h+YrwcQbF/FVjWp7ufi0noRwpsDzEc0uAtkcmbDk0WLiMAS
X+G/tYxxCdE+fZbGXwsFJ4VB75uI+W1yjE1zLGetqzL2Cd/Ndw4x8F1XcX5sIQuF5KUi0HMXjv2s
GRqV5SAyx3UsOKx9Vi3p5TvwPGZTjudpxtY6yUyV748i9Um/O8cBMJP0PWSoacJXNCCp65DFs5Cr
MtpXdaf2RBJdAOlRBHTmmzUHVZxk7ODRMhBxuS7xcT2dyMSVf1yee7UYZZDN8cRhXsNtQLVMBsM4
r3uYg1htJC/B+MXrUB6bbUK8kFCB96QypcyI39EyAPll/kaF2JS3NSBnNBWqKbrTlFrGniNa2WAC
rFdpjZ8u+R2rlAhNiq1Q0HoRaE3qZqSS8+S3T90fDtHtc4x8bPkcgTjzqR7YZ1jpI1TO+r6xLC9k
8e3qp+gNXFfo2Yd1k4ZQpmgxzzyCxNXTTNVAZcwfwL2ITXy9aY5T0EYkvunjpBp3WPN8FeWbaPUj
FnUTfMEesP8MZfj/q0Hvi+4bLvYa03LXVGMK4qhDtTikXHzA0DM6Z6TnsSFSjPPNn+FNriv8/b/g
OSkK7hNeYLzsTWupJWUuCpBNDk/Nnq3AosISGEwfg70UWkg6vnwPvy3B7vkqP3jCev9ubdCorbiV
l9wG+HKKpOTM5oX178TYNPDKcY0V+/Dh1VJp6XUgdRoYF+/FxyKG5E8tyMGTROtCkK8t4f/z+Qjj
7dqhGBT6R8NqVXgxEGpYIiAdBkOCnOE++3C7IRuKSkgFakZ9PJj9YkvA0K44QUf6tBMilZ7Bmav0
JFsf9c2XtmEERe+aogWxKGSLHh8VB6Mr747aN3L5jMpvnmwxUL4gl7I4369JUpnt1HmX4S45OWIO
X1BonNSMq4WTbG+c1MdCEt2k8/k4PuTaj7A5ey9VZJYEV1lsju6qu3g2R1YayouMIWKCEKIUp+L0
vfVZDTjgu4ZnaEhM3LDj6PHjFuCO7/Wu6i7kaRqJ0nKK182deRcsURkiZsur8tAU83jmpFE8pl/O
PZj1UM15UnQFuY90yHSt2DrRiLBF9eeQI+vm7Uu2lEqYuCGoxjTL1mpBtbWYXMRX9vMcQWMqmriK
c4QYPjczVmYeqlpDguvSZDracJclolg1Tj5B9rS+6oHWkpIS66Tej3gTKGIUSYIIc4HRqkwvaCsP
2ISsTtxFq/Fq7KpK5F7Hxs4CfMsNTp08cCV2Zl5Jn/+TmmbJUxn3nqY/UiIp8r/zNlRHLCHmVgKf
3EGaXiAtOKtCyQBhUdkiHlBZhhUW0WY6lsOoQEsJsVWbBcnwADkm6uveA+k2TcAzEJvHdGUDt0xw
PWfvCZL+B3bqynQXbVQihzBvZKv675dVJTxnuVAJaYYN338dFRZETok2eec78J80IUIkIvwtAxTN
37g0QOQRVaXoLTIz7qPOyAHOgv2SZYWxMJ8x8n4POIBvr/Qa5SH6CWyURP/VeqHQ1QL4aCOk3Uv1
GqCcmNDGggvN+7kNEpnfF1IrTfBBAKV7HyR6owE4yYHdwD6SqqzEfIgLzitilTWnOIzUAjTsn2OT
Ewr0cN0Rvk0vKGtzyRZOD2imgVyQVoRwcPUf70mABR+6NNFitaOyvDAeC+mynbluLEH+NMG4riK6
6eZUGoIrVen9y2Xl0hdvd5Ss5tX2uV2lhXZpWlzq5BypbrUh8X5qzv8CqV3gZhqAa0tR85DmfO+H
PqSzPGK1X6lI9hmIXlX81+7r8JnUNcpvMcuK7ZkcMzy+xFLm+HMNycSSgvYoNIo0CaN7nO1H4iwi
Hu43G2o1EVtvUaasztJ+LoaUiMgJclQWB1daVcu4rXm4Pz9VtHOqAmwe5c7s/DRompr067TN+/i8
qnfxrsFdf/4f6Li97PlBZ+SBNsM+U6l9xr3vKh+7MMVghfqO8uzhSMSHtXR8p1un7M6NIWdskjSi
4ne/TVive8uYlL8/fodfvKerfEHW4L27gMkmOjRNg+tCmpnARVrYamdjbaQaQmqB0tZxHgIy55QL
W+GBrW+TDgleZReTBzN8DImEQH51zB5vHV1t3Gxg+ww5xBkP4CXfsf8t2RkIn87LCj3W3u44dMII
ukbKCG031Y+zb4prlJC4f4LmWzHWrfoA1gcAF1ZsbFSSORXjFiZ5mWAjOF/mqrGiBuxmRvvT8azG
j+IgnXnla2b/boGz2Yb3+J3h4B1fcRd32FCzN+ycbEaGXRPG6gpv9ftRzOtrXXauEMXPAE96Z09C
5cIS/mMFsUt9I/G5ZnbIun5D4wfNYdxAxBs9TjR1HSMKizcd2vaAa8nRRpipT9yfIjCzQOB3JnAh
KpTdSR2KscGG7643+pTnJVlF3XpB4nP6hXmU6VLNgYhMLINKEd/HwiDeduRBq+qXvQ8NtnvevU8r
LLztU75CkPVpL+1CSNfpbomUTudTwf5affVExQIDJTpuc2ea5mGwW+4oPZdB4sl1GyUHug9AjBz2
UchQ1USPCvXFqSy3FScnoKIZjCt/o0hx6w29TCQ8wPjUX/TzCEx2kaaxOUgQAgJgyE0YNW2wWMxd
w/66lEQptmUFHi5i9QDBHgNoqd+1bavHhlM4M/oROOUJzpTGs4T3lJDAtUo9fVAUrUAFdrAsOCaW
+IFGch7Nt5in0VNzH6NaLzRaBowo1oucSe8KPZglKtznRJpQpn+qi7B4dk/voxudFmQeKmcrGq+n
Y7n5IC1rUtv0PL/OwF+JtGPB0sSbjd7JphayEu/XKFX8gTZydRMJc8MjzWoYInkDzHvbOykAXhoe
CiwuCwMZpTFi8SvzVQH0Uz4N5Y4DQVgjnnS5X0nBJ8Z8krqPa2o3aHY4Otpr0dPfXIHvCf+gm/3s
RdaYs8AsBQv4eFZPIOZA88/yFABc1xP+4SlBLErFjeUEN53Evq5EZg6TbSKD78XQ+ho8me+4BEc2
eKu5q87Vrh3JGxSKRJcDXAu9DXVXatP0edblz8CdQP0BOtgR9STz/0/on2Vk38k7ORKEDw6NbF+P
CV0M/Nmh0Od8G/aCnVwuB2BSxVNPcTbs6ZjTKsqoNaGPNbmFckm/ZpgR2A1orx2VGqSI/otWrPtk
/gX/tbHTIxGyT1jr1BEwusdR2yx1mFcbyD+vdIvGQg3j4hCkSOEjG/Zm4qa8MGVNmz6ohv+h24AC
Lk9rXAA6QqxBaoIMBdD+4BPWvrTtKF61H2j77ISnWnKDNyT77IdURrk/Hgntmr/rbhzlmtznoFhv
EWGXuGrDgmCv9/f4gbifJNGVouQQQqUmxivmqcq9GOoin3j2HuOM6OWyWjBBcuYivqbPHoctLhug
rQLBAZBuzYJ93bszrm8yFYqwhQJ06ZcKfrHrDXnq2rVVgI+Q0SuZmqyX7YS/btaOhf1WvWgAGVRc
oudimJxhIXWUJJf1RSJSh3mgf2z5qvP17OAziW4hFru1osxGPwWs2aDW15Q9w1GJhc/pdz61Y+HE
YwXXC8qG4n8fkEibyJ6KVdOkTsaTkOXMe1ql/1F9HtFDX7vtvgSrPVp5NlMuslG6/59ET/plTqtF
lhUy33UArrTxcaFj6aQQ6yIXVvdmlacJ9zTBk6u5HARD1F3km6ZqvgIOjOSjMk25V+PxxqLB4t5J
oJS9WympWQJ2UOhmM7m0rC9DXACbTGScB9ikrai2i8yZJk7MxAM+ZJdZ6v3IXvwTIS1NTMLXu2sj
4BKV6Seuq+iz7Qz6Np8moK/FWYZIDvPcItrwu8aTGQu9+uh/P8J66GkSp75dC4SLcuJ/Yptz0xjD
gLOu8lQ1n+n3OvuRqnL0OSpvZXouh2ZyQSeJ99Qo5BrupdVSkzlLGx+c5Jejl6r4TVocx4Did6XN
pS7Qb7xG4af4oa1fzsOI6vIZVtyQaqJi09saoAtHJFm2NlisPVZSv2Zdn3ljsWW2ZT6f1JwgdnCz
NSL8mifo5h1w7gWuUDmyCqFFZQ83CWYKUAvuskod+/nsAxYymhW3f8rzoPtcVlhKNM5cB6iNYVWS
X9y/4MPxJ3W1NNNsnaxwSU8Ea3SHxiC7GuvqzABMpzZUXwZiTWKb6/zlqtO/zkZ1WOUwviJzzLeU
wWGG4V/sGfnTqAzfAXUpNX2mVTw7nxIyi8apELkbsEJ9EzH6IVZbP/VAQArVD8oWU0WRhzy4agRd
/sa/8DybIgDJGCG9JM/HoAJIttg/JR9lMK6mVZe5iQ2WO3oGSt2SqZIw54CxOVwlwlmW2VXgIbxp
WG70sfKeh/lZGtCvuEz5iM27DiDq8VuVzDgJA4Vw5pFm1FHUp1wKAZ2ptSk9Qy49Jc5u9E5VxwXE
5gqFGu0hFF+RnBwYwGzeVgKFDeyf6NTAizc+C0qRmlVxiQ+29MnevLULnGbxxGEPzY1EG1BYpfIg
vSQzYoeD3U4FMjiWnw0XWLkH8ke+EpfB0g+eKw+sJ4j1tV0CsDUmPB4TAhoViR8EalMDCLr/PyDt
LS1f1gEnmSWRtX6ec1Obo49BUsnMs6CdPReC2DHSbH7R90tbkx9HJ3/aHq5/2p2qx8elv6sU4Q4N
4DQCkFDBjd5wkwKTVQrM9xZWPQyUfIOn6U3XhHQblUiqC89MI7jukCsq33f08H6luoHo14nKQa7E
Omgf+S97TzpsD2t0mligxzsuwkgo7MVtZ9++gMvwK9slLPfB4xjmTdADXlpAJg6X0zVk8Z4BoX0T
SwvRh+h40emm1KNrr9YR6u8wKOe+828S9iW2uqsv0z6lkQZIBnRJ05pDneBfEYg+pgPlVM6ojg9D
LONMtrzs0enVw8n7vVlyPnnEOT/97+zPIfSz2UG+fMDA21Jdko80gaO0qFqnwXFylQXdf07wvcWC
2aaZ4+eGqjZ+4TMwHgCmamyDT/oij7dzFhYXT4DExXc1HpFPNway9Wd0GbLEvnZFqJbaEVBKtxNe
MbsbaoUYH9AC6kpp6AKcNyc/V1j9oUSv/HW+Nz9gknRFgUyygm5fQChqA0xMdNEcpKZC0ewJDZiy
3u+mtAOdQmpeH2t3imyB4O7mXrQKq0bOmgnuhC3zbnS2sVYW2mJh4fPv1GDtBd8ydC4+zCQOV91J
6iJBCvcOG9zSEJM+wO5vd3pcCoYIoqncXZ9eYNAqFrxW42Y7XGlPEyNoDH6N3dNQGJ+Kf9ro4eGD
LFAn0DxTF1mOyOepceWR9VJSXFIxjxeHIXQFY0et9+jW9bamz3fYzsg5Fo16v/wgWC+q6xOwRCn6
s9ZP5eGnzOhK3zel0/GfAaC1V61O1e3K911CMQ8hPC3QBLAM9vFyWLHw8QoZzXsnOOsqbgD4xBO7
5NzTvpkuk1zcpsmRJXQcZPl+yECEegbZs9hTVQDTDRlVKGwdDSTpOzw6vRCNvB+tFIDaRWi0SCmI
NIlVQIp0TA4wbvTNL0vGA3h7svkXWjwoxSpArleByq8E1CuxN5oMUMrSV0PDqXY9s8Ugyn+xE7aD
GEP/ky4BoxLJl2HALAQ8PvwWG+/LKfeZQjpAUB8Ps3L7PO1oonYwSHvtI6yvtUboQxrJbrlDY917
OGO99fTzU/Dt/pybTcbFunKavSxotQhhR9bZvr7Jaof9USDgnXxLiBpR0yz7OQT2cAGzFvPyk3Es
cmKnqXyyT0Bp5A3Nvm3tXJuKdcFTm8gT32Ka+s7Y6xWdvI45wubB8IhrjmK555DZAC/o/IACPVVg
3JTTJOoVJvdnJ8LgDYVOlCvfEO92xRf66+bi9/z6ZHAqzIR6HKDsNOYG2Im6lgcZWUQeZJ84/k7x
RhVfD5ZoXDVbfUf1HDN4H8a4PMFe2RfMOk9ZkS5AgKPTXeekqqYesjEWQIgdhT73sU7t5pkBxe9D
veLnYI0IgD9CLOxMoPlC6jH9vV9VRunmviLzvwIdEPKO+sDu+sih6emVJ6ROioUH4Fp6iBz4zwhw
fhn9IGTfMAZMwEkKupLWzMV9L/Zq7eV2VWjrDN0crKcyfJL0u/8gqt+N/7mPc/jjC9AhhH2mRyZK
Vz07chL2Ik52vdG15IwCWxvXDwSoWQACmUIW8QWBLYUjY6Rz9nRCxxkXsA1PqcCxpgqiaimFRT+X
kzCqAynn7JSSfJmYFIjg/La9rkSo50jwscS8B4v4CjoeTSQKHrDxyhFUPrggNJMlI/I7lg984Asn
XeRXDjxtUWM0ikN0oflXWDqaWcK1MeA8GIpuKWa8qI0OfsJCmfrijjYqzIMPo9+O8fSAsZ/CsJoN
G+PurG6xFXC4SssjsOkyO9tJazRSQc9yppON8Pb52WvHpgGUbECQEHCj8YKGgAzbxQz7RMJpEQD/
S8lH057Rk4mPqDjRra0KuMms6kF/E7D60VY6a917VLH7bbI+5DzM4LetvrurF0lNLycxivzQMyq/
tJ8fnQxz2jEeB+M19o8x21LyozDkRkUvoPNpDjfnjs+Tnn+hNg5GtgPfGX2nJK0rSTXyQL7j0NZL
gYmo9ztcCQB0iiZz4ivohObaKURhTgcWs0rbFbbRL8VQDstgoKw5vVZQCF5xesifn5+h4q4Y002V
JwW/YyZciVROqIdpxYnGBpQbGAgV0uDLDDyu/X6ySVqc2wTE8CPbrp7QBBmT9TSlgMj9iJB2n31r
FoKzKjJwq9Fs6bffKc6eUVKr1iwIp/lbIFgn8REhUMOaANsKX+ElGyauP0LCiyIYTmb3bX2ZpeRc
mlZiB0+jmypFcihC7o1DIuGByW99mugakiTaPaFEjJg0Jqq0mPxHv1g5nExtr/FLzib3nV0z670V
Js+6jhitW9bi8pZLmg14AJ/VoxvmInMkQ9vSTu3qid8jbtNDu78lpk43VnPYEm608l7hgWiyDf1V
Zcm7nrVFCwJYeMpRByH2IN9BRnXEF9nSq3kS8eZx0ed7oZr0qXzOKmJ0mGvi/eEcq6MNbmS6/IZy
py0qwe/xqJQM6eH2066fZXzPe2pp3bEhTY2Nb7B/NzczKQczk300vFDvg+C5FeJQG5RnXxk3h+47
5ENR4SfkYZSKdj1IYpE/3MqUhEXavkLUnOm1y4lDbcWYL+0QMZQjrxaEY1JFVNmjVtkZkUEucnrU
KLUZHeDjfmRy170OGDEbT69DZoeEoc+vmcs4yVDe7hCvkxrg6iSw8WmegbcJaeLuW6UyEaa9zUjJ
Z97e8xyCUme50xoR64qdYpfHfQ/t1jhk0wOC8K9lO1SRAMbU3Gz7xd+ziEO0Rsl4AGVypKlt0u5f
zntYDQ6DSsyrUVE+9en4Q409VumB0jlgMtsgYWGsN7vVSpP2/BfGsm40ROyaTg1cToc4ZBdJNoY1
xanHEb25w0YLMi3BqJ4pCUvuDrEVQ+BWl26jHb0jfQf+Xj44y02Pe+KJAIeve7LVjxjDnKrYUcHu
ilBcNyKMmV/EJg75HuQFcAbbuWhZZy1UC7nK/fgBP5u1joCi+fTNUfEZPrW75rjRvCHgP43z804l
mBlDNAF8t03wuu7eL3iVcKFXjU2iYywzw1gt+dH9QETL3GvHbqOmEEtWHjZ1gzZy+DtccrJJkrzf
CIFtqm21WsWhUoS1hR8A86OwMzeg+1rYVyR7CcPZf61A/4K4CKX9Qx4Y6e3YeDn62SM0gdI6lUI/
ex6y6h/jUeBPPxYTpG4whqQC2ULX+Vw5YmX3rKBtALnEoMvo9cXNxGTeJMk3ZgNgQr8xazNOKquW
HfgKENpbU4gR6tRRli0CHZTqLCtN0S2xOPyTebd/oOAx/+7snjaSA85OfLk+pUk0XL+984erUoNs
KEfHmOA0bhCPVs2Mgs/GIUNErYN9bwoCIPyf1a1RWj0V0uk/qr7Sbm6o58jJEZmqT2f2G1of7U8p
4ximSJC7LD5RC+cF5g0mVphvSNEdh+Zrg7pEETA/cxKyDXfw1OrVhe/MThvkuIBlRH8+CRQcnrWw
m2qy5k1P/r07G54V28KSXNHXWGi2lrSndW325nxMVfXqKHec7jhNhZswdsHTZcd/y97skBBAJ4NF
2U3gX84IUUZePNoNNrOmK0qzNT6AbBBCLnl2QAGjmwLShfVI3zhskxWzmVVNl/7LI0vBln/iOU3e
7f3x9oszAHahXwCeeGfSvnkTUO/Z+rTDlmxypsdmxGT10PmBg/do6tYZboDqErwiPKKQrEUhf0G2
Vnxy1Sxm7BSI26FoZU4J8dSG6C1f1lBQanM1HUEk5n1a65yAbkdnqZBfSfiS1kQ1vfPfN+8RLx5g
PT/BMI/GHQBy+UfNQy8aRNsy8y3QqYYdZ8LLI8Q4L8wbt06No7vsfh3weXc5Zrq0HDivOSGqbxpc
vSPm1MSvQeoNlOIwt6qw/74cKzaDPhRtQftLl8J5iOKl8ZG7Wa2bzAVxyYU+wGEi+VN1m2j0iyZ3
c/CMySVpn6XIi+eOFi4iJl4z1amMFVY35kIyUERjnkppwR6xFDV4HecKE8Dc7ZUBXah0Ee9Dvlen
WW/0tBD4nJCyI3ZVPKe25xLgb/BOI0xTVrkW6NBgnWT6F+KMObii9wU9h35HOigg4eKxKbA3g17E
G6B0+sfiPukApmCjCAmNicGhLsFL5rUUDPQpp05pzAfo8GxTb45ZnQw7hT1IvprOUGGmzv1m16VQ
p5hL8rEfbmkKCajeY1Ku/QVT8nY91OxXazfefTIYNxFZSBgb26G1tw5PtReLpWSZ8d0UaeJv2ne3
Fb7wRmzyER0c3fKu4fm95yrMOb2knFtac/J2PFTg8eENA24/KUJox1udukAyJq9Ur3bsqeCWiUBM
lvMH4ME+YyBQYkSGmt/M1MngRpK2fFRsuOTdRBIpj5ESf/8Nm7eNaiAzXKxbAIhWMSsXY2n+Dkgr
uWeUSRsl8ynGsrTpk5kGGw0bF0RO4nP79ddLzEgetXx1c4dZJlX4/DHufYsquYHZk4keV/OudMP0
otYmx+Oh4ccBXhMorEZ/s+IvOQ2I7nX+M87P/J0g2dcLWRHWicWjr52GtaBZ/2hFl+sejF+0C6aT
ivkfMB3VePSNsO6kUBwjc+jmU/ZXRfcP9ta0yGyCEKnG6hm8l26XMvgC2kRnSwtbIK4bEnOGrokh
r+Ot55W3FxlBNXe7Pc7NgRrYBtsOGVmGmeWTNiNVT8dHBl3f5CBMQPmgBLwN2sDil2DDgLOk/I8c
NRv3Pcs/GW/Uds2GnyxbGeWx+Ygt8VPjesCpir/P7QPIPTD0wGizH4xJ8hQrdG54lo0Q4M0Zc8Tc
d6P+KGSDSWpKp4Kl5LQIbP97pn1XpQRrczM2+M9+x5EQoIQ7yrlatkmoS2XZ3uiJ9uoeYyRRPO2B
3uPwju3yfLSDoO/D6Vs7luOmhg3+dl7up1OMQLEtvZ4Se5u6DbDPHKmQVUdDU2WoLQ5vZw1m4UeQ
FJAlKJCRTbTdn2s/qzutm4ME3AKPpobVL3CQcFFNTx/ZJJnjXyL+7GWxjzvpu1aB6WdZbkR8LLap
aYrR53sMXOvi6UQixbe6fKOnB+Q+bmUby9X5UtRpKKg0YAWTjOyhKlzXpNqjj5RJN8G+sK6oskVt
ImZoy3odZdCTqsLWipHVt+FHlPQoHlz4hSE7BPMU6JA4jPZIWEdXx1MIBhe/d5pJIunkA8VecDgb
Jik59EcmelYtr5NWUvEhdSFmwCgk/1q8Pex76U8SnYR5PYOmIG/ChkQEbhAYbIxfL8Js76y5W+rf
ftejA1C2AaTEuJy59hERHD4YiZSSXt9e34n5Y8LpvHpIOo862V/Zg73wp3n0sqgEpD6/ZRg3KXBA
DLr4/JUryBPv2MDcxQjHGd+GRmwYmN+oXpjlADVkMW3IYQUnYbfptQyBAxnr/sWld+FVrChqA2KP
EbgpGBRGxA8mYafL7Yx244UKAoeNBPAvhTjnkyRJE+LbkuMjioAlV1I3KkgU8HtH45TEkT+M9RiB
MLcPPNRhQTVdV/DhsDHxYVfMgKb6RRY7VDp/rdCmwGevvA+hBPe1KTh4YJOUZjszkkj/0D+JsmqP
2b+rjVJ54W6WtsW8vqC3cgwZ6SvImAwtUm15KAh1DNrB8FpRguJq6x8n6WX0poaab95y9uKRhKO9
tt6uKwkpNi6Vd7pGxLCmWEj5fChAYLaGvd3rHf3G36Ar1DgOLGFk36nx3ZZx6elZfMqTq1aXXxMz
qGOpYfMVDKfXgyYhusZQAJEErHtJ2dxgOY+xgDc8Z66vZdkMNSxqPB4YQRrjRFnBt28pqsm04hkX
BESFQ3PxkRoqgTRE/xvBLSa8HxA9S6AZ1xUxsjLpmhiskadFwVytDOOWyhLus1Sul+y93VeGsMhr
6Ow2uvGVQDFlnhSnOUNYnaMTWn1uBjvW/FltwJ5bUDxqdK4MvkQqFPI2mpsa6o64IvkpobhpA+8q
zrTxRHvpNJxgXYKbcsd5VFFssUORxYW0BiKcEmP2AotYCXGtPYn2Muq0ifNqL9FmxtLijYpxjfVe
wsi7fnQn93LSaFm8bUKrCpE4NZ9tNQzn/aXy27h3GCAL3eMFMMuNzdrxWhDMWK5ddEUXliFMi50V
f933sxUp2woPMnLo2X8t1YcDraDI1EbVAG0+Bs/3QGAh8of3EZRH/7eR+dTPDYfDCuUnlFs/0A8s
QP4DGZFYmUunCHZY7PCkJWzVNTSJXC/i7AKqh33Odd3+kkpHxu7a0JyPOiJgcolw7rKMyJ9ZTPAH
9N1mzApiBzeYmbMEgEMqGXy8tVAnREDbmtUrQnFO6Xphb3OsQzevXIs9nUARfGZvkuWNL4pESGIW
mGBJ1XhLhBZBtmrqc8D0dSMqAe4A5yQ+3if85aHxy1riWteNkLlZxcfVW9YWXZMun8AfaQ6gc7Hq
FMn/luorIh9JiP/m7W1qCRENTBAxelTkjBrBpuDhb5zt0WQZOOVcCj+08JQC4Rq56nfkPJnQ31DY
pPeW1ngXwGB7lkVo6zJEmeWuSSBcYS3nQJUqYQB+DjHBl843sljeMVQS37KL6bILdl3el4H0n1Ok
7GWI2OZxBntuQCgX2KlgPnkhBeV2zO7qD0bTiP/2XtynSw51LHWBE6HL4hOpW6SV7AWuocPPWCC1
1NNT0Muohl6Q1SPF1Vvk4LnrZGCQHVDaGiut3JoqJq1TtgfUDqhA06Mn9eb3gdupteqVGkC9LKdL
Qz/9UD0Nl/cjPQP1xMWtqaZJyyNJJAyXjWuPvQQzL/HbnlWF1qDZKL2WPVQAT0OPxjXv/PG9NieV
Qk3EUJxoDAmnYxN00O2EhxJhZp+W796/dcpwZdWfCuXWEK7X29nqlulOfEizfLVbuK+bqzjOp+8z
WJtB0L48GUDFsKVM3hxdydQmVGn7OuWatTKnUZ05LKoAx75bfttsvdZaPPp4kPKA6DxwuHE0KuIP
/kSBAyFprmYZnofXP5UNz0g7CKaYVq4B6uufLwsekhG5bF0h1eojTfyjl7EMNPmMMj6+tTd/ZClY
VJmdp2YnTqlnjGTiCxKBYWLyuqkwDCqR/1n1vziIKGBJNm9RoYDGvQ9bV8PFnaMMxc7kF37zH+iA
EeMJlTsPDg8fdbsBh9vsp4eMNjyWSzp9z0rN5Jt9GksDBp1xL6kjuANErEGjh6uOA6pDMNBMLdyX
zRDKpY+GohY/mKG6hx0PZUFkB1qwgZG4UC3ufvY0VzbZQmmO0wpR/Nptk0IOKiBwgudPfPEBljhg
u4D5LkQDWiYJucBHgeb29heKU81phdStdaXChdlRZ1R+AlNBcMZuZbFuwgdOUcLHUyI6xK0V4nJp
7pDP/D9JSryFhvNPVxMMSoJBRX68l96R3+xvfoTS1rq2S88RylaZux1OqEHn5+KbTg8SCetdbBte
q4KWciPPxRSAle0ZRp0q/NN6jlQo+J5q7BFE6nf+kx4HoiwENqnW1KI7TdXfTPAYo2OIqqfNktMm
XNIsNW+5169rtX1jhk4l7kTN2hEeWRoU6Cegb8Ih4+6dk2Zn6RO7gnJIWLBb64zIGhRKjPXbeneN
hjPq0pfuqHHMnBsxsMMAUf8AITHxl0npMyaCI4MSXWNxdegUTPRPGHkO2zMKN97PdP59i0nDOSD5
Um1fCGg6pOyUzcn44STPuD7BJ5lTigj0t1l3OnjhKjTKmkTV6VhaeS/QM0E43sm8ttM3o273pUFG
P8iaTQS0SNp04zHvx+9OwvRjUWLPXhM/c1QDi3CyO0xGfOUtLzaC93Ja8l36n+2i8sM6QNxK2wPo
5iQqLiel+MwFkIvynVh1lXkwGzAmXLa+7JTXehofhF65rO5e4ApAGmRdlkONw/uIBphjpQozoq8S
RU/jtEPFfiVEImxAkV3d/f3q55kKJ4J0UjnK7UanrVOYpQv2iN7zKeO9H+rpj9BLQDRvy1oTJQgi
/aZ5YNeZzWXA5fcR3rFnd7ytKMD+8KZVi6JV7kOxIx8YA+ECGvY29lrKsGTkwIRNIoK+tjPvecut
dGoX7lUn3/3d0R6hauFpaXJHaWHAYKPv0MZoqDfkxblgorfTGLtJl8THxVB4WHSfANuj8p0/pkwl
NrbY3ATLbFAs4JOsm3s/xIS6msRwwh/asKqHN+EwH+rHX3T2VtwgetWbhHuXhIgoPnGh4wmW8aXh
9+UU7ybFiK8jFBY6BnNixQxdMxnot0cCoVbYGpYpE5vcJsNyieAVfa/eLWP7FzQHihGMekgSKwk1
n6EwyZDq40t/OVGuxIC+wXdaxa1WaEsQs2DqLeP2i8Glz75yT6njLs3qUq8YaKp7dJf2xpzCeBAa
SRTBn0YRuLZDGOLQ0Y27CA1kJFkX/KABlDH3ONh5+8REdOrwMCd3kfReIDcz9wofIPnFrVfJhqOm
ctPUo/HO69PpCSCJ+rEJmOFiWNgVnf0AU/0d6F4FyapBKa8Uo9+YmmTYH2mS6Lu+K3eG0YGRAq6m
Cyn+XJGAc6+7L8E6940+wW3vB8Hkc/9J6gQKvVc2uJexTQu4qp8aBjo4WB9br9SgyQGslmNE2vnh
QT1Kt+qCK0pJbOoemP94bcJWoTcnYX2KsNCPwro+se/H34SYfukF66Pp1qfxCQHK03nsmg3edZv3
WykbdfwBDZddSG0JShpk1OVKGgYIjhLCinwbsRRIiAR6g8he+/pOBx6c7tFI1PTnngwXaer5P6G3
RZfEk9eU65M9hU6a0BtJzL8njFDJFzcV8czIse/JdWjvSLIBTZU5kXL4q/bNsnVxzWGT3AIW9EZe
GtSrr5HvzMvKBSg9lVAqvOl/gvxSqUrk6BfaFy5WIbs/1Tw0TgAaL2GLoD0veaML849+9EVgkf7J
6xAABhowC8sY6kvJHKbsCGZsVU6no7Z5buwl5tfewgtRfkqj1+jjrTA+qHqR42SI4TYbvgFVZBWN
6e3s/pUvzZqKDrCTvDskwdVR7MgMgHHd3j8GeNIClvDS5Uf/QUdKkymXpGxhKAqLnC7E0BGTZ7P+
PkwyRW+2QrcCNjF+DiBf9okb0NlThHPz3x6LgXAoHXExxmJ9kQ3WD3DzjjBw3/CtUuvZmkB9TsCN
Sm2pAzjiLMgxzCcI0IeQw+8zGM2tD43ywjOXnOd9F9o2Hrf26C0ATCJnio7e2VdgLfm7bSbcqohO
9eoMhlektc8xmIvibpVNAUXcdh5lCiZQ7eDqJ8w0NhOgUIvlMLlYjd/qcbsFyViRrq9tG6eI35Zs
frNLUbpvkpd7lenY4+tslNSydahdIzReHHxLn1ap5TxbJFZ+XbBvsFTwpyE98lUYJyG9PY6dpRZn
GmBEwZltP1ynKAF1ymSEJj9JOUg4JLDBEJFqAbtE8O4/lPE4ZlpvfEg8WunfKTp0xw8ehggPCngZ
JK0E3SUWbeCWTDTfbRQtqTvuKAmtlhEdVJRy4fCMoRE9C3s3rnen+Tk7X6yaoc1SPfbOslMImfSI
hhSGK/j1j2VK7foF6+gPdGqUROkpMMvJP5TckAeTl2aQ9AQn2uw61TUC9SxYIrANLY4fIwfxJSgm
g9mLmSOfQBZoO9tCyR7T36YVqRYP9rUgnNR4G9lv/rie5ZQcq9VwcyO1Ae6ZGMHcH6Z4ktGQGRRm
UG98zTwT6GcqK7EAOOFAJ/a0MU2qjwa2U0gLxkRs0o32qwlZN0gCX/Ve/K0DlhRNn8aa8SF5VdKQ
k1oFeNC8OhdZ4jBvMspdWktWnDgYUgrn9LnooSTE95jtmEm7viTmCe8a1lTkAq8BUEGl5egXHlrS
OIjBc6Djv1ucRSFeNhpgX9Zw0nz3E0leRY+2uKxLXEqeGrAlzeduFn786odQFzZrg57KX+WF6Tx9
9LXifU95+1fgFEGQg4w8Y2ZbPhDMPL9cw1pBnlXNn7XyE8+famE8241dGdhmMrUblchOrhkgw3FG
KLvxb0MB/ZiZZfFI2t9G6C1/VZsN72Vp4G6a8sWB7pLtuk3o2aulgXYqT8uiCya9zMCRzQKyOLAm
zV55sNj6dncZtmqTotGPOh4WATooGd9C8zYFtGZKx9y0KgiE3cbi/BiE9N6S9J5bXT1t+5168WkV
I1n/j27ev+ovSzaFrc9BnmORvZuSSsETC+hV26t+EnkJiRiNBDPpeiXMXNX6bHyiQbyz3KVAq/ND
xuU06G7CESYex8ISV+XEEnrsj6Zfw57UyGk+Dx00KP+VPBMAGOT1dGho7bLsJbZP+gdI+MNoIYGd
ruo18uqea1vCBWXTXazOnKuFb3YTu7aumUsARjf7EdZ+PF5/g3uWSqKwKsrNmciFLzrfcMcwXO5V
upi+oxkAe/b1yzrF4m/TR/IM8l9+2mqm9ePfidnJSKTcj1/kj+ptUVaRMbk5K1q6xRGkCzkRW961
6GhCOHoF9ORoqEqf/gHOVNS5PlZScf9wn6voyX4V2JK19Pb1IIYRvP7+Rqw5PcasLTxE0iAzQuS6
e0Mpq/Xi7pNBUGdZgwMqSVhLc7EZzEfhf46w+ibOOyzEqtzlGm65fE4sVXQwYlT9ztIJRqmhsZqm
9msXcVfM6JPXBwYqir3CoPpPXHDpUK/Af466IuWdhXW+bIFVSKtMKj8SeIgsB7x1MsUxSu/CMWQC
V7qgwNwGGbHohIrUovbeRndRmlNKNAfyzpdSSYckwzTupl60vPSnahSjq4JTFFSDlTfd5FPchbxJ
6K0uUOkg34GvJHeIrZ3CrUcssK0xCcAXUepqtyKtNkievDY3ZMwPXsHMaSwY3SzmSFxegY/GRyGa
2GGu+2cXiPDiIykEqto0RfR84BLKxlesVgh6gsZb76JZLI48phOddkr/00jWR8ibqJUBFHRAP+fZ
6CYeTJ3piIA8lO0Tr9NQu5l4BvUepvX/+nEZD9dy6N3EruY2gmmQQMMapn7j0oLNjhYWFuEFqjWi
zrJ1ACUwI7iFDT6SuOR0Cp8mJfNoiRU19mDnz3+xEIKxKrW9YNH7YQE1pZPppUB5kE3ZfMpqjtY7
MrI8Sq7dGndGls4V+S9Vm0X1WGc3/qnn5NqKjriTbWWWDr9ugf/oUjQ2i7iLhOw1Tvn7YTopLLvs
zpM+SURHAcvH3iMaMwNh0O33ewrmal6t3I1tGfTLQ5IivZAmPdRk6lGV8O+MO5rUTwrn5MiQLo5N
n/d4Cy5D+RR7jF7WQI6t7p+3xhEIfCjeIi1cG/xVYMeOLoSXYCI5ibdegzL3OUoqRkElZwYRpY43
9qWcioJdBNn9afwWQAYi96xMP5OqRmPo3zwj7ZsjC7rQVN5DlcCF/oTOkMWc/GuWKK5DACp8vXbB
DOYfE0pFQ+fBnhhBc4Vt29za3Ag3lwOXnWo8qMZ1W4X+A9dW0/FTlzJ7vYOcgQRzeIkDg5Txcb0e
30IUa6Kov2tXLqoEJ0i6RqfpdUKfuYJiV/Eneo2C9gZpBYWcyC2k97qNX8y+fDD7/7Q5fcUsYuSU
7FFGNeJe9qiHTdhCAOwewSiZ3ae+PsoscKaFD3V3eOsaJdWMFwVnjdfTY0OQv+bwiXmp1UHCm+Q/
nmkAJ4/kWT7eEhb7r+PfIbXB7UIpdad/gT9iWXo5NilqE2YaHLCd3VwXngwysS10JsBXD1ZaXPLa
Hx1GvzzwSMfMx3rpTttsfTU3V6Hi0z2VlCOLTKXIo+vqghLYcQwQlWgC/EN9SUv+hK1on6ATMDRq
2t7gwAqMP15IeZ+qfLwUsuY632qeym5FbiWTx9OqWR8j9XnmWyPMgaUoOnWnDQrdvpOcaDr9eEaw
bmY+YXrbz8jPk8LqcHRkzdiMNcOQdSRKQ8k0YmklbYt/XaTKlOwoc3jLOOgYageRSPbifb/ciMVd
CKpqooz5HOL4r0bQrhlK9zVPB6fUFesOfLWiIau6IGebqcKKk9gUyJi0K62+jSKqmSZXgOpDLeMI
AKvsIQY0Pf7HbXXJ9Itg9cdYQcxC+s1+5LcjbgC9HHWizk1DMtrNhKXC3EDpK6cuzmD/NvRzXJOY
naASVTc5dRi2kSQpuMCNquW0pON2uOxqXErsNkx4widrJ69uDs/bXDd7NBGE2i9ja8ffvSHCY2wv
OQlcdtd9Fefk5LkEMAWhhYOHuvVlokjiDfBjKNjPVmCacxBwa6OrnkZdoHVhFEh94KNc8YWBaZhl
EHBpMMROlp67RnFcKbmEAAPQi372PBSqL7xkZtF6vgjd/Qtkvt53CvT1RArWirHp+CBwpFsz9Zh/
nzyKKPv6NY19GqTvexFg0Dr9/nhEbpVyR8b8YTtds9xPcYHvUBZLNLInUUazB/gkMxGjmFCdC2l5
5Xrays1r553jaZmSn61jSlMfRJmDm3yzZdIceAaPRQmRdsneR04eWYXQBrRc/CLG6e/vvFkprUtJ
ph6TFg3VERIod3dIrYWtadFh+FbHUpXg6+4c4D7QYxm5EFwdL+7QJpNs10dn3JvPKVTWUe1XmIeg
epp1VYNendZwZkbayp4Aq5nyPQ0l0kH+Za+PWgcPJHFN3pwBDJiEYIMj96yjeYNEdkT1YY/FaqHv
GzLHZSqOPQGFTj+0+iOW4+LXVpOnwFD3hl9v/7wvDLPkHvXKQ7dpSxFML+uBuxvyrGq2lBYuWwYC
h945ZxQO7q7BKJXFTMWyDSnujfwYisVckaSExZf0sYG3nnl7I6pQiFMQCWdgBa78cXcWpY3X/LTl
mw+ueschxZYMKUuhQTIpldCxIPNa3aWKU0eeVPuFrefX/JWr1q/6MRmcvpYX431QO1cbXkJgq+fH
It50MRJOkz+bXgFOjEbr4/fltmsQVcKUr0lq+tc6x5AHPyzQyxD1v0ubTf4yIUJ3o+j3Y5sFdZDR
q4bjWK6wBjcJ4GC1prCAu0DQ6OeWIN4Ze3zgTYwz2rnckdtMy5K7F0N7/khTHaXFqqeWqShg1He6
T/+2gNYD+Zm9tgOh9JNQPMZS/GycxemXFiyM9FHby7ehvURYbAQF8b5q03zNJaCx3mCR4b5UMQ5S
mvNArrfVi+mUgR/U+G3ESMjNLd0AwwDuWjAIF0I338+OPt7JKLjZoCfZNmURJJJeBtn6pXWU79Yw
MIGNr7j5Q1F46gVIKXfY0tbt7kTkzFDIaR38gnGXKNJatovHJWwnfQqb3DMe07nhQj0xYKBlRhN3
V/87Jcg+FkHg9aEzrBrZGRfBAk6WU9nac0ycHtua+i60dxPHLNOZT46Hf4OJdOUMXRdCcojHyTTK
U+kHi3+ul0HxT6NC8r3xm4k3tZcn565EzqEUWJYWMV0UQxELRxwtdX2zWFmqBL0q5B2GoNHIPIGT
5a/6dq3bsJlsZfYt06C7JAyTLCu6oVAPg60GLtqJH7pH6d3Ker1k35inu+CdcLseguNzt+VxBS9F
hbHT/lphBXoZJvvDeV7qJARuR3onOv5kny1M5lrdoJqwQC2FsW8eXUZv3e3OE0zYtggceRQwgjlV
48s42LgrdKnmU6dzvzoKV5EJoZWqZ92WggT0HGlMaj307vmDWUmbdv+gxsfSJQwGPOxKDR+5yRuv
cNw9rSlx4dk1JZfu4caKePKblPVrJN22MjV1c60NTn/UqGFif0c2Kuj87J9VIkDaUi6zc406xsEZ
cpHmSqdgQxLd9XmGn2+fc/ggdpqFPp5VmHDw0UXtbnmCOpw8Mdd8mkte+Ixp4hZtg7iDDZiXY2Ez
uX236qRK8icGWcU8wSCgdGKkpiZ8epFo7d4miNWuC1nN7BjJhzHVPEdKO6DI81b36qJ6Q1Xw/JWC
lb+uJ/l84nJVJmYKj0bF3XbkX3aPFlMMKDUH1zZMB9ODDu4hhXfykOFVr9vF07PhGaE+mspuZN5r
J1duo5W9fzdCIeFQECYqoOMpsNLApEYZKmHnuRd7TgEPP+1x/Iea/qdFJGBMl0/lmKB5iWdxXpyg
ysO3Pvj1rtrPdcyRTy86JZXLKBHRoGL8UGOgZhl62d8mZFa2Xy88riddN241bIhufhKz5QGkoTTV
GLyeZVCCJAT1DkVAwu2F/hcLlnBOsHAAoJOZYU1zrNhQlgGHP0nB6s7MKyC1F6djaJA4twFDkpK9
QTsSaxM/iih9ScTOhPQ4xq6gH1WtT5LfhPwg13wbuRR2lD+YX/GEbVC6lKRih8ppqILFENp8jYFy
Xa1ZUz7xThPi/xVGiwcC9ybmJiJIIO2sGYSjDwz58MbLgdLcmSWlJTTLW0ACz3p4oEwGkBWjVN70
DkUzXFaXq3Idzu/erI1BkjF5FDhfBgCnXkElu29qo/XivofRiYN7jFmCSpmhvOxCcCYxIIOqJSzb
lkbdO4n27Ohu5z/8mAi0JaMCjMxScZneSdnBMQtgIVVNUSmLlkFSzh0DtJDb640XJNo0qmyHFOIe
2Z9gXEIf1T6uyDdJgpU2Kf88wFHQAraUURZAsObO2hySykBTrc2MH+H+1sHyyFiqfqefbF/HTuTI
3PSeII9ANv4jt60kI1n448swL6h/RyepMTXx1RxlnhyHMvx5I/KjTlUVLzdxlWXvBn/C5Hzg9E0I
hvkyv/85tFskVdVo+n/Xq3h/sYOt+JSaEeZv46itAzA8FmUYV4Bi5vBty7Y4m7c+uVFHCdkxotC6
CT8nRAtffOiSew7ZXhLkAL8vit4bKBAxYaRWNx0bNxa8Mfi5tMdoUEVI6XCrZp7buye3y3+Y/HGN
hnqqb2IHa5+T3w6NKV2fiMGgFZZex02MY28w8P/QgPgcu1RxvfCoLxWziI/pQD8DO4QNhbj9kmy6
v9VntyJ+TFtLYNNSCzsmCzfQkjJCddNozyAmX3AdD6FzmulcrO8er3Spo7xBXMJkM/x5prC6XlOk
vS90P/im6QZ9hyCeNXWZa8cKaOhVy/EE/Y9d8VI7nT6pOCnv5wGa4eKXXOfg2fS3svdSrQ/YBLPb
AxkTRSbh7hd0l061h4b5YZkFXhin4ZhI3ymI5eppu4YQHCpxz0aT19+3KGbbUD/knm6hfD9IDwxG
oZNwktIsv0Ul/dxw2NaF7im3M3F6uzf0wkli42SGJpW3n2jIYiCyCm78ZlvL6JR4uxJxGjPrj/kY
yU9Ii6lkrpLAkE+lJqZlb9P9UeIeCu/jXUf1536yyeFP7dyvBit50dRx+GiPKPYlQaE46GWhNuW2
GrycwPBhEEyYWe8hY6hlRAKxXwCx+ws+bJnOygQWAYvlyaJqNpHs2yTjkyFGx1In1O+L4GPKAG8i
Frov2xh0MU2swBIpzFK8gwTAehnrY5Z+wxgpUIXsZPYivflZJ5868FmagzBlcZsUtzN9Bxyj/fq3
xA+RFmXS/oSmpC+UPVM0Qkm+DyNYj6wbux52xvKFyv3RPYx3ssJVHuQsuUVelB+FEHtwzWKYOC5W
Q6XNRSK4GYIHL8tUc2YSZeT14pDaj3eR5+CoPf7ADKYtZR1glfUCrKGaj4f8N3KVDARbheKAORFJ
iHmw+xp8qhW+zrHmp/AB78zCzvG6xzUoHHJGgTwCVBILMPGGZD9trMKvlftsVjzHExvOTabKRUDD
yX9BZ3tafFHB36PpWOQjj8aelF8dEpP7QzgINf9rvp6o8ZP0RWqku5L7zgKVivcNXHsf/RzVIHXn
CMlDZ8VloprUGJ3VYES1cfpvp5dh2mBWa4fhWBXVRPj3XlU5TXyt1SgRIT3DhdhLZPrVMUEeL106
bFMtm6jQ96H6BJx32+HTV8mIwA7gN9hE2czUIdcLy0bq+GDvR495yvh4R/cXT/cGDhz16cg+IHAy
F9/XjXeAIbgoBldhePC8gV0fgDOGBrN6mzvcNR7QnLHZJ2F07Vm0irvURYssDPefs9iye3U0J8Q9
7PU0/uHZExxwWB2fqAIXINn7ERq1q5THY71cSwMMpMKGfnZzFOvzklZeFmsKrZFmZ1FqToNntAGq
1P094+gVFlOt+x6Bl160tA2DkH1L9s/FV3NmbeGpYULjqERGYh0MvRcTUp2xwjeh3V9k0mlbwsPJ
9SH7/bfYDshPFM4S0TT4g3HqCx9iDXWtFxnVmxvGjNfhVsxf0ABLhFUjPqDm4weEejH6FZNwusaL
f4f47AFv8UM/h5eLGF1l7eVADQEUnbkxD1FucMn2v1o3cRpZY1v1aUZ/+KT0G4P/HyXlnpv4iwBg
/Cp/Qm4jZFe9L/5gQszpDjq/p+RVU1pxi5xBftJ1Lq7OnZ7W6BhhcMuRsjfGRYqcnltnsAodV8qi
tgT3zvoxtWqQw2lig4x4W/cDaA4WgZo3TchvhVNDRJQHxdu8Y2kQU9tbs8b73Jfmr+Kxy5+SiVga
8GXy/AiCag8ZFnyskpGFET/Gob6FQYiQEZzhB7GoYz7PY1uL+vgFlANEpatmdS3II16X/nOFSDsm
6ndmNapo++XMcehYySUZONYgYpXgnLkeri7mDkTr0ff5EoKiCEDBcRWX5oQxeJ5wZqbGDDclg480
xR3QRAb0CpthVoYOF+TA7FhzcK069jw4ybVEibb9mZ6DwufnueLRYxxRJaqxrglVPRRrvFS0YtsI
0OCoP27HpNIPXBWnWYR2kB6mI6bF6czPhZOn3vvdHEVMU+8w3DB/5qP5xxLYF8K3M7eR73G95M73
2niAZhouMajLf9/htg++sk4xukv5gNEhbHaFtsGmkCJ91CwuQ0xGb0fB21mpVb7LkedRt8qtCUNA
DItFNfo/Gw5ym9GuDKu6J7WdkHms46iqW51grs6DjCIHh3ZSoo7mUZ/Hq3HgDiHo9mOwT3tDR2nO
4aWlkSCTjw5cVgMUtu7gTgKWlcVzXbgSrcDwbgk5/cwk57yt0Uny0Z7SySXpQVdcKrMy24O1Bf8V
r2iYNxX49VY2eo74ed9xeW9ukGkAT2F6iN7Vz3M3ynYdymJwSHB64UThbMPg+P5j7mnG3di3iLKx
Tg8qSAzCoVSjWoF428lOPmW+art3TRyNdAkRRI3fBXEfoNR30KgWwy3vFbJDFrw9a1L+Y421Nljk
Vn6CAY3gdz5sQylJqmRqXK6rtkGHfgNP3SoFKNpXhLJL+nIXlAVbh0D5/B9pO5au17LvU1K61Ba9
FNdj07RATziQzWB3mRh9VcqzUtC3QNoyTfo5Fjki3L4/DK/SCI7l2IVigIUBZg/wuaWBRrdOqH+2
Ruc3qN4M9+bBpEYjmqM2cPpV4M4ahcOFQxQvIG+5QqMtHHsQ5j9PIrO5Xf9pOfbCjCe/n/dvEOci
33b+oenUvo6N2wSX3g65DJROxxsjaEQihbBfOwKvGqQFXbi1iaq4aZPUJjx1iMA7KPtws/3cc518
tiitQVaKOX61AmI6wjJiBqTup0tj+E9xNu9tKqRXJCeRJcpgsdNC/aXd8OTlfFfdchLDXfLjlqlt
jzPtI75M86OKfC3LWaeGL5uKZJ6kXwA8VEEPWoGb23t1fk0bLNwV7uHF6TUdPp6ARYbLuHBBuSU9
NjPbmZXWIa1rBlKQTtPs46uVgW3L8EqJx3bjIeWWTixtQQgl6kFo9bVnRJfFnnnVLRakYN6tK03w
hTXzraBbg69CbS2BJhv88FB4iRqXHCPE1VcDGCAPpnjIpD0295GFG7yxWcCs5oYYd1a4390EJZfb
JR/qPy5b8y93+27JrgjRSTulCt4JSAZ4TzizzDMJiHA2HgD/VBN38gdCeo2HOgaaE97QqosK7NzB
6EhL4NlgLtTXuTFleMFuY6h4zqvUG/EZ0mIONRUU4E3MrbqALJZjeA1b+hM2x7jbT9tZST2GNp9t
H8YlBx8NpD1Lc4Q8YkcLsC9Wx8bLB1KHrAILQaTpDRWPrNlnonVvy54rr67IHDPz1aYYbAYMUs/C
U2BKztiIMTR5HRvR49/w4Gpo4E20yglA/Dl30KhYkmn/khJ0RJRw0Qx82p/wn+8lJjg1hJuS+CiO
e5qgyGadAIMfvispbBuv8zR1ytNfOWnqsjmpZaM2KZTHHobUGHo+y6/BIA+Xk7nw5n46zTYUPmVD
RcdrvCMJHm9e1ns61ukfCUJKaBqxki2sdVv/UUBTZCXazeNs8qiXgTQd19Dzh/bw18MXtQhf2M9R
n6ZObuVv5T15lmH+mz9E4r0vUU6JGT9edK29UisepGZmEDUo13Cy0g+mmoycgrXI+Bgui8yc5OHg
zQQUVNXk1dCzJv9v8B3mndoOH8vLo9achfv73O0WtHkAewAaNsRtYN7HFeywD7evAyWc8U5Pju1m
zTgeUPS7fvkGiIXPo5AZbN5qHtXm416q2pBXl5PFqBRPVTumol+WxufWjAwJ1LY9odP3UhkWakvE
Q7j5cpk5MuOuirM3Q39fY79KTrt5xDlHKrE3vM4BS/lgKvOdIhgxrM7StRhk/HwldH6qJqn/QIKa
zZQ1D5VEyCKcdJ7fFtLsLYcmOXDB0xQrIec00ctzc+Hnz0WzfRf5YqnpTbR8GUZngysxHwXPKEnR
4/kpzK05P6sSlHrMcl9aw5MiI6/xNTgI2zHL8kxLZHfriRB8QgEzXXVDPShBY+BXfMSl5vSt1wbB
5ye1YikJAEkO6Y2PvkMUULjMOSqzNPdA6LSRjE1YUl/98I7xgpSkHh19VJDIdnqQp5NaRO+aJjnd
VGWC2zx8KdKq3T8NwbG6QNs+BimI+YVMbDVsDYfTp4ZKVwAK8GNZr8vUfgUzRRexHw0oPHa+34/1
qICSro+91jf5x/XdBcKqYEW/cOpr+CZkrrPS5NAP7wruvuikkrXHre/jKKNOACPfdt6nU4pYyLGU
X9IyafyVeEPyumAsDI1PyF8XCD2gWb1C2OtkmfdO08FthTPVDF7ElBj9Mwmqn5XtpsUByQaLtaB7
ujALy+8MYT1xT3RypW8wUR6GHsAejpFo/IfTecR+ltJou555sTdU4LjuR+yiC1Hk+yINNdaecFW5
MPPos7TZrcHXIpBD3oO6PskXjOW6BtpvnrZw/FtlhKYi0g0l9+BDyfeqEGAWbbHSW+wQ8jjs9p/D
wT+VO2jDmqnxiIXhwHGLVL3nytXd2g5hJ0YrbhY2gGCCMt+ngZyFbfVSqmg6mvwKUArfKRU435O6
+zMi1w/N8kAZe7OV+p37In50zcS87WAIZNswuJKzjeB0I7r3asMV9HEGY5a7Tw1d7h3zqy1SDyIJ
h+Ds7V4txL38/QSIFJlgmiPOzqR8APj8dtOe9owi58n/T4/5An3Y6PWIljNUKIiAdthOzfoEqYTE
PN6D1K6dXxx+qd3hS5UXvYux9ffF1XYQtcmL/30GKtl9W48QoFi1/mzGsI0xBOLkme/VvddfSijv
/YzvkbvVvFiArlho0rjhcDYQOgk0SVSWbH72G9DkBeolMS4aXXjW4JHG5/MDyUlyJYWkEUQshQiQ
6L7KgScT75MQt0pErR7eukd6Zz0QDpI9OJH2kriujepKIM9ycKWz19vCbYAW6ilnI2V7LwsjRcDG
hZV5/3GA/6Q5DwT1i7cyCFTQ0/IBlGrbe1RkjR3iY0I1rj8bSGEeRrG1yd4S76ps7uT26V89LO3+
isS8NUglE2iQiK7+pZrd4P2IC5MsnRv1UxWsMnMx4XZWBT3L1aj/As+lt+lMPGDJh0/LFbTA/p/i
c5Lna2kEm81mPlHmU5e23dWK/3n4fXcs1z8TWLH8vKbX6sbkiY7+DLR0bP+Uz+YBrnpKmxsyy5zj
uDnbkNg+y+hTfPekmlzlhkgaoAab4ta9x/4xJY1222JdltYkROdw0kJ/9ULESzVMk0vl3Z7ZtWs7
tQ2Fdk7+Hh9VAqmnM65Skfu/hweEY51fbMkVx4LPAnRPUwBu6f6OXXhvAzND3ASfQsNkwbaABC+U
3AWahg9Up5/Z78cNVMuV1upKVVHmb7ExvI80ae1za4LYK+LIfgdfOZB7GdZUYSaN3Jw2Ugborqdq
2oaCyneGABZXM9njW+yHcUlin9TQc2K+frYG4nb9tMqbbfaXQbchykY/Oj2Y8Gm6PdfjnGLp8N/y
TNeTQ2HlnimtVlQvtWEdPDNdkxMpMgkt5bFULKz96XK6eNDQu+xT+nvk476sYOSMuTlA61HUCJwr
whSoqCprfd7zjmVNtdoQtobAUHifwGW5ZZ0NmVkIHTRrOU7D2cvBLVrint5YBrRDgtyzxba3lP/t
oMaliGxut7+ckXg25+e3rWyrLs6f9+4odnt4MvHro9+IbEQ7UpmFJYx3fKvyiikJEUapm/uWjQNG
4zqN9rzDIWbqQT2C4BkfMgceX4v5O12vTI6Mj26FtkmsHqRjMXVbbhk7uFe/xoli4bTLXVlfNltU
oueiYKAxtAlsgBMYiFBirnSVaYOTkvdvmSmXytpWVhVVDdG30LAy1awg/j2BLQxL6qqMVWRshy+2
QqrtYkfyzd0DVdS/y3/tjaWD30FOWATGXnWPdFDJi5YF4JjWgihYnXOKnn94NA4wSyXst1upEr7D
k6MmweL0z9GxDWRPkEhkWC2cxMnHAjTQdI3ZNHl6oOJu6DlOhgzRFc0dqGuI5JbGaEnSTmQyGzyS
HeW1c7oBB0WuIGEllbg7i5sUavz+mKmELyCXUW3ocHmDFPfWByn02BNmbeeGBSaZ4RemeFuPM3N2
3irDCUWAo2w+pnJdRHep5bNCTz1bW10t1krvRtp287F4tEVl76qth97ONCkmfUlz5X8AwIQ4I2Dx
nEusUcW0Wn3DLwM/PnA7krW2zGqgkSvkyGbP0vvX1/JuJYjpaKygiaacJdj6KHjgECI3VQ5lx/Sh
8UQ8e8vrR3fy5SNTyaXtWiaJagnZy5lVFT2pi0876PzHcTxujfmmpdD1q+sRb+ReuXlcVT1mFyTR
MJQn6bgmsoIz0yD1qE1wwt9/IW+Vtyi1ec8JbDO+kMWc4tW+ObRJ0EAhBUDdzUtht76d6yxiX0u+
80hI1yk+XaZkple5yJsKHqVAcJEB+5XRILOJnn9z5h1jZIx2t9UHR3ikdSk3BJmPxmu9z2hPGd8V
Jdxu/G8ImUv24UspLzrE4MVHQsQfOpB84NlsHS5pWf6PJb4HtzA7slA/WoPwHcNf5whPVTxGLTqd
GG3djliF7TIW+uuufnsc87Vh7nZpSMYKsLuE3yy6cUXXxJUljrqYag4pVuP26zHYuoYpZUKspxQf
rUwx+skdKEQqB+4a2MjkY0MVZXGwKt+EpMnIWs4D+fL3WmB3ftr2DgDJ5siDwtc8x7mCnDzbhmNL
gdmbr0wDNWVbdSLFdtad0SoJnhZuBxXROmktAq7A/5jypJttogoN1pBpbq3r/h5Kv4jlh+EVvurL
hS6xhzdjkXa4PsKw+5x8/mbi8fauZ71nlRzn96EUUeP//TT/m2VFCqacIbqMPsAfwKx92o/tIXl3
qg6aBFLLTeq3j+uRWo6DDI0KsJy4mjNPI4xcJl7oElD2xMDkh1JJHnYHGQ4D1h6COuJdVGwolpOa
ayDb+OM8MMu6eUePdFzg+yByqUA/njuOUCXycGtstjOdsZdD/fIi4Vphm62rcuwupRTdrzfszZZq
sByWxgZPyqcKIr2AMMNl0eMWjFRlU6HY2ADDAMEOy0iuwk1ewb9DhNqbwxNg/bPHRckfmHTHDI+Z
Twoh0Fj8HTRphZun+z6xKDGCRZM4oqA4rMqQZt3GwHqP8F86tt9xoD5Sl5IQDVlHlAADEeajNm1p
gHSLZQLBiSYET+qjDllupWg/s4xlvVf4sIxrMOzrpyWp51vi/uk084T3WebRLJPs8sihLZRiw/Zk
SY/s2i8Bg/Ognum38xaQM3n7VVm0HvhrHmUerdXjNctMrkcJ5byNd8PWv+kMSZNZeLadqQygbnna
DfdggBnI5AVMAjNNEeiB8LjT42MZAQ6LcBnZKL3L/0dp9Z1F8Fpq9HbySHFyX4gnR38wQHXohiDr
CKvKLZAF07mq422tWM0zJ567bN6etfygVXUd+2CG0ohulitDcDboK5lkEeeCqHvwL+fFnSDcsloi
eaa10vYoTkEICq43adUxOHXiy/ks+7gcm/R/52hUKJg2EAMKFBgcvUDxEU5kht0YcuD3q4Asr9gD
cxKcLaUAN9GhHhLZWlFAYcS5WBW4+x/cAMsAvO/Z3n6+qGdzR3nZxaF0BnlTALSeMNWsynEHnQCs
4heXnUYHCtNDN8lJ4QGAncCtGFYlNU5IqDRP/gjm04kzBlCtRJ3tIJu43/dixsRKYgWS2XxSmYhE
EuVoqy7WcoaJNubB0Pg2gCJXBiH5V4DDftjXThuGB10S/ZQB6+g4F+ux2b681FQ9Fpl/xXGUyXTy
rI+PKxAA/Sq0+QY14UwgQvVNtTeCjw9oNq8D32tsid0Db3bWkHo5DeithtBNg6gUlQ6+mFW2YVou
IOgujZh7WLBy7tsNeYRKeBwU+J93frd9zeel6TnvcIkktgtca/Y/BhrL9LPZYDqMpG/n7HTKLYIo
L2zOH/81jM3AsT0hLfo0jERGZpIWNubM3xLY0OAWXrVtGgDO3twOI4iRok0lMWNUspFdpOBpu3vv
QAU8WfDVbONbDTfW5wKGK97qNh6K54kFfTEqlOvAkQPnOxCxC5mnsOLlYjDc+Av+fiQqfJbiywpU
q9dZd48OSGjqdZewEr4CmCfUhuxZcXbPFpsNz5yNosCEhqhrWjqVgz+2FfqYYbXqehkswHz+c0rg
u0q1gam9buANgYh78T8m78oZg/C2efeaVQiU1gUXsUz8V81xDWc9KCfh5JO0dFwihADCXwjhg4H4
UZG2xud6oOBkFKxxPkbx0QUg7KWsGfA74GYQNcL4nZ+hsO1qYcAtOR7S13UP8Edu2vQQZ/ojZuRF
Hgnvfmumf8pySX5Por1djPo6OdZU0LGzI7YojiNOeGSXeXp/iOspFrWmSPgYUu0NQoHLjrQV2N5o
lcjRfCIHp45tj+E2hfH0Mv+2joyv76LscFPmqYiLI4U6ZAHkx+l0yTauGPqgvPp/C2QDSJBb6paY
L1tzxMD1mmoZ0Ed4AwUMkrcp6PtouNigGjwcAl7SRvx8/2LLrYz3jRsB9YyEY2BaiNBfxoBEGAPy
nJu6t50QeH+YSXZ3is2+74A6EsUP59D0OpMk8aCCaMMIGGb1gwbEozPcqeOckCdsKN/PLWG8iAc6
30hv7H/64KvAx5YLucrh8lc9R4PL4ajHDfktrl7UIVpxhGaQDMsZ7UopiqNg/hxxDRrhPrlCUJpk
A+DL/E7O4Y5zg1QMUCjA4ekACdq/tgCNbNCfc7SmplA/XW+u3rVMaP5lNHk3KU3nn6xxPKjo8g3F
r1ZbEgdLCRaHaHoIwSMn7Twj4U6m7TuGu1f0Sj6g9ccdzkxUGGh6tDtO+B0ziyybuBCup6eqD6lV
t4smanUxp9z1xPMWPC7jmUjHppzgAXnDGDKFjVOn6kyxxm5gaPc3w71OFbAGJwODc1LuOAWWbfVm
0XxkKYtmSOTQB3woJgXbmmuYSmtx8vKsalQs0lCtlhAh3Y2+QIulXzoKjo8zxCG4K3WW7kzuuwO8
jMRrMqFtyyLc4WFGy9kTfyDZyGoa0XNE2LJFiAqAY2iYYJ4ZYIY64chaFdn1woqPrZvmq1JfY8t9
bcOBFC2XIvKiCXcGP4sCDNnLrx6/4JhbXXfckYTrILBDti7Ep6og0TcI0Fym+KY6gCT5pt0TI4Q/
VrVWuKyRp/CBkBZPC+NJIhxIR0xKy5sycLVtaE8mdyDWmRrS7EvMvyK1K03zW4z9h3ow8Nd7hNWZ
kMJn3uX816dpIccVDimruN/Ek1S4o32My53AFHbC+o6vQyzP9nLifwTkpmo8FHnkdbhZA6M80GTl
kw1QaG/92IBEKlkHfRzC6k8BZoA2cRetLPEMVtJ4pjIgFP4ijV50Iq0hZlcz9YbDCbo6riqljyQP
yVdfZwycoFVepy27G4egmbpI7TuaBFJD6S7bXwCWN0VTXlLxKr+RmxxJOaQaNJCB/W2+t1aUQx0i
SZqLbnSY6WnlDlFeziXOfS32Yna7+jj4Xd2MOrziSa89sDvSWrsi9Zal4SIXwFSF5eSHQPzYrmIX
AG3sl9DMGryd2/GHfA3g3zLaZTQGsHNv4OiqAqptkTFyO9I/TGPBV06H1+Svgccvj11YHZrxiAm+
3uGq0tHJJ61DG0yWtiqNLoOKRRTRf7odId4Z35wigDx9CttIvdKpKYVmpxdr2A7Yb6es2kNd0BO1
egP4Ev6fZAY+wmurU5qq8cZvlXfH4Bt8rlFPQFelYzeaVoXz68Yvulp8w20OaUucssZEvf4v9TBe
FndBn5xKh7A1fUUxaXYNiC8va6O7KO/zvyVapI874OpFtfTBLm/WnmpCcXan238lkGakW5hiItvp
KkyyDU9zJWMEV6YRaj5uXaspNDRkC9ndau6CSIDXPZ3+7ByUy3misGPzcYEEU4o2HFkonGy1gB5N
LMSWBxjqjSaXBE3D4B58QsEALNqUaOPMrEwwyGvgzCbpmmt7DVfveJttf2OnT8TKRcFZ5T5DIZu8
3lJPO7Q1EiLM4HkT7zFIlbDyH5xpyktPe8duloknSm7E3h8sAeIZK2CdX/jlMdX69paKEUx2omxo
jJwRZuteakJqkloHzy0MApQ18qHfWq64ijQkC4c+HPMtZbw64Qh5xINI5aVHOtK96k60GCRlW9JO
9TbpjBzhBclvWTKVN3kY4lGol0VN95cNXciNisuKxpOP65qwhU6F/vsLAr6OhzivB+XT2RS5PwFg
O0dNKOPvizHgUNzDm333HW7CUrDqidWBRNTed8B2Ncf533jKpOTPb/XhThDiMxYaTewaAKKwuEmZ
/vKI2FqM3ZbQEFdJURS14koJ4qfKanmAki1oOrudsdizklKldArChvTcNdCBM6iZmlN116evsc2V
K3Xm0Q+S3NY3lqRk24A2ZNRzwgadddXoeBZoKQp576jijCTr2wcIrSPJSADZgluqMTM6nPW+laS7
fuaL2cknxxSfNS4w8BLG++MRsgh6P1i/IYb1N/LORYLU0+iRqRKGHVgYwbZRKwU3Lqc5DF4d5+cG
0f7jpD+AtEYGzd2GGj5grGc1FN5ZHQvPPzJYHzTDecBCljET+etFQy3EXHFjGSLGNoJEIkXX9I2J
PptunWDx9fUCbvNsoZXrT6S8EkPbB6gb8qVUP5TuiIzorGepffLzjkDr3UbqfpPzXeHTcRXr75X2
znA1CmQsVU8E8IqMN9Q2oIC+ahOpAWJkM3HURCpPKAovAvXV/K5qRm8cFY7Pp81mYQ2uFHu0hCeU
ykfRpmf8mlJXZY1/HuwHGDxCFuSL55ZoGNkaqeCYBG/Jyb7TcmOzYZAb6KiWcOee+8zQLsjzRb/1
TzYHzWP6w8OaOOayz3Wx6UB82RmGasdpAwv0AclNdlwcg+ggtWH04aiG1IzXz4tl/iAyEtRH6rwN
LTgzHVvP6d9eynLiLMIp+kA7yYmIjWx30v09MlE+BQQSO99BXncr7ZtlF5T/An6KZ2PCF70PHDx0
rg5ZkEG80cQdd2c/0MfBnvtJhPYM2GNAtI6KLgpaopW32FnHeMuJI5aPpn24MTxXvQ8Ph3xEDXtL
fxVAvL86yVNMi+EVZQM7kTCZb/HdMAw7mDHfShrbgUabUU+3dDYZa/48XixdBZb171+T36ARUTpV
G5S7OvYJ1GHebsFFPbfnhBjxa3seHcP499PVXd/lnGfXUsuWJ1aqbxekvb86mcABshIYTg2RnmS7
qhlxzwBQoefFYFxqfw7JApLyS08YbgYNVXoHaipu2cBgsbZ1dNn6aOhOpoGvPJqRDHXh9y5QkOd4
T7wx24Rs0BtpPDe+ivkICthUhbuQkgX8A+J85DkV0fFcuhFt7VJ8dMhxwfUrlPjJsgaru1QWOlJj
ydgxo/kZlxw7NDaS76mNP8a3aWSNn/svSJUJCiyg5cDF8VucapdeLfjzbFC7J2Poc5lM8V8XVA9w
P0N+5ILIYUFFwO6Zr/hhz6RHQPxQsVrWRq8hPX9xzRG6giuuwIyXn/xKwZPuBbUaLFEB32rRYFBP
kNgKUZgmZkwIaAlE03jNM/+CFSIwI67Ib0tklfeczwXMB3ztEoWj687cvZZdfKJ6E7ETlfKkD7JL
qY8cpUcOJ1ifGrZIwdgKCZT927+KX9dbqDeiIdJWR5mrsYQQVGNNGqc130Iqvh6ZZw4NY1kzSgeV
cj6u6jcmaQxt7YyHaKKGjI5jm8wG9PqIBn5KU1Trz9+9c6FiH0eSdeKTv7k6zO27oAceP3tY+1N0
4IQwWSg0HGCovcuymkLh50zVJg9JfPSLc6LCsYBKlThS1i4d4sDxAM8VmjkkdUIHAAifNvFEovUj
ZmJ1GzjW/4gEGcxD8be6p8cL95142UPcelZd/o8bZnAFsJN1E/pxh1+wi57u+ro8m8+ki+BShLQz
0y0V4ybgaYbUYhvmaWzyj3oOWPLAbmNTr1ps9LMn0dc2FredsZ4RGL1l2of6YxVurl6abHeFnkHa
CquoWBuTqQwmHzDyjl7UVQ/UfQooDa5DyzSUmVymyhOQTdG1u3LLWOBVomC/dF6m8VS4aqlUH8GS
9uM5s6/Kll05yaco+Y/reUyqNc8Ym4rZITIBwAM8m8RXrVVrm4+0wkWRSx8+nV3NKhwhO/y2raHi
b0Oi+qWqiYdrI9jraGox1QNyPFPMAEhApUXhX6MwxJWl1AksJM+gIfcV/Q8rVnTqim9iTuK5KvSN
rUhAnPtTbdKvVmt2T0fug3xEe/o05uBjNafgNvrZe0icqAQaNUH/K39haC7cKz3Aezh675tiQ4jy
h9neIIhc9d2LpgIMjGDEyIihGa82PHQ4g1BAWKOhl/sF5dVcpIEnFbQHMohmyXSimh5rIq2sJWTv
XDmGq+P9Jrp+AW3OVEZ5p2MwALCU5oUUBQA3xKNH3C47eP6svVpvM2e/iJSp0o7NmQgj0k9hVjCw
tdc2YGTV+U2Gq+dgNivxk3diRVc+OZ6Mqiz8GwHOLbtr1ApvgU6Y90aJRvkhcFYaIBnXh5VQ9kqT
aDzVzsx5hAkky9R0XE0X3uk9ojiyB3u4eA4ewCKBAH6Jef4trVOFZKCws817mDO0+vYQ6vEfsS+I
9wbntMZv3IIi6sVEUJ4CIbWjM0yLA7XS7UPAF+AhPbWii2m0NjH6m26sXbzyduNxWBug2U9BVYCs
yovYRY9hjIWAMeFdjKqrYN4PK6PpGVyN1/P6bry0nUq2rWcyv07eMgHnOs8nTKa2qQEtLcJd/70Q
HfyDiDYpdE80pxC6VLGIccrp+iW4wZ14R6FAAkiRMksSErTzKexLQnj8vS5h1VPb30z+t8eu1gMS
unTbwGPXlTyHcRV0xtVBTHHIKXXfDiEVCij1fS/G3bnxhsDQM41BqAwnC5zFvUrivyQVFVdT8wIv
FPpszPqBJ7Gr+1sYNpveTmJJW7o0/KSuqo2NSXULJmWLf+HZX6qp1ERhUSePVsjJk9X3vyBxzfl8
H1sRhOSwHOTZOsrnwNnO9mmhKmZd5Ga8SN57UNbHtatCXahJ2X23JY34fW6dGkl8UFQltvfP4PfW
VioSHC3DbbUEbrQT8jDc04fWTt4goDhHk4hvoI0JldW1z5hdAsQVF59xW3Uenj1y2aOYXzd+e3CK
sl2DBMLkfP4AxITkceOt0kgKNBkvEyqE8O0VfpiInOFSulGPXDGInYuaHuPm7p5y3g6Hbd6jDBMg
5EkjZ61hw6dz7Md5V7pr/pPLYUsBs9JNE1E8xbyweJkB6CtRmVxwzJQuAEIGJdHTt6dI49GlksvJ
bk9S3TCJwG1zskw0uVZd12/DK74Kyj+0sRBNzFKyxYF1bnUkMY7LHxnkzMn4HV3OUW3h03DKv4s8
7XQLjfdMAqadr0G26mjTwmz7WZyWguhqCy4u8/slxkfmmUnOBpEkeXPbzFvZpw9gmlCfa9hc99m9
nUyqPYi/ZXZzkK8SPIA5qY1ukgQ/V4jxWNWe9RSSLNzS2RTmsaCWyWfZIDNqNGZcITjYaWLhxjs1
al+Wcv+d4lNdixra3dqLWHLAOv9q9hSivh6hv7O/pVTfYSgWnwr2Cvu4fO0PqwCMmfAYQH2xtlge
haDskckPL7Zrl15oyG9aD5FCxhfk5uA6bBwY5m7Y3ldkFuqwtmLSpSHhW4OC0TtAUxNEYPNWKUEv
owbZbhPbgeLi+unDEFvnS1tg41FhT6khEBe2o49AbESGt01QeH/skT87t69+opL7BWp3Jrk2Oey4
cegq5ZYyEAwhRr0cEpH0p9hla4kc3s1UmMnQ2JRngL34HulcIPAhkiYdZgQR7Q6myqC049qmfHgw
Yug+VnPKy+yDS+F61Zzj3iXyCSrgR949lmFpLSzYUQNoeOcRtmgZLQiM5g9sliJ9WBWFZRnRo2Ja
mtZM6G39QglsOjkMH9W7J+4MrZOrAFIBkhlBJSUHWzhVc0UoD0LSkwWU5785Ps8Aqf6QqZoSOL4F
rXq+O3xT17PYKGQNyE+b7wQhStZ5OyB8vrrxe/LvSyHO+YCfGbu1SRcYK60PBBnU7Zye27AG5jNW
zk8Lj56J56/xm/xpHlJEYEmN/4CAaNOO4hvVfaqPTkcGWoMIFvtTI84JJ3UUbEliLIhYl8L1X400
+5+DGzDrpZRPcCzwEQw1whHiyl0HdAP5tk8o2pbbnV1jLt33U7n6i2kt1InmC7mfeajYAZHUQr1Y
1SKPZl7afxb7Ju2SjumgGpntoeqi4uAnRO8pbF5Kdao/20ah8yp8ONfi8nCqXHiFZuqvXl1ydH3c
4NRYN23YB3+gjrBGenasxu7M7CCit0afXixRvn7ok/hr4NSdY8JvwIpYrF3HQIHxRAE5Ghrj8Fv3
R9Uv3iEYhq0e09DxiImg22CGiy/RRbSFHW4fmUnNG4T/cbwhyWUCheq4lw3C4qZCAKZ/wv/JXJ3W
zWKxFnXRiM/vD2Xadvhp1tbRe5jR8M0wZaDpNV7SJudLriYMqcLy9ZMKbpk61Us5xN+wtCFFeVQa
PbSh5c6ZXh81qt4rlWWU0KjTJie5ODV7f5RAXALrS5G2daRtU5mEz+3BBXIFrTKRHDDqTNyki4BF
sNVtxIZ0k5j0DY9wmDJiTZjxev2QuGFbyTGHNer0y7AG831u17hZOmW2ruq6+FlZwyflgTlv43Ep
e0vVv/676eQWnELIEII4mOxHeg4mTJv9h/sMbPndX7rttT5OUKVDLh7Kc4xyerBqZw+1ZP2zIE1W
swbVFOgedjnp5y4T3zZN0cZ7CdaZKuNaQ5tnAAfMgJEzxj6THDMXBPn6tdKvRzAXgO01L68Jzk3c
KfVYX3ammqRdmSuoKywTsyESqCphc48YINx8TH+BfS6yL96mhheVuT6zcj7hvXT6/y5PcRzooeUP
t3o7ZkltmlTqF1V/0jOGZzekj61ae1c831fcMX94J6GO3Yo2EwSp9uG+peO9Dd0TRphL9NMKk7DX
4Fpd/F/dq7J2Mim2EUwrfJhvlDQ/ACmOOB1qt4e+P+YM1YnJY7hjGNgbcf8V07CzxHtf91Tm57PO
pKgP7bF+iqi4gcUrClx+ItEYrMHavqqtemUbNqjkNG9qrEcYYNdUgbMOWztsXViG0JbNpLKTkZ8S
BvwjoIiONcdjQ+dZ+Q/AlfXn52zbgt499hEP22sjEB+KMu/mbN47zMH+nfhELYwKMB/KTQEfsgGd
lPhEXgueKnNe+vgwll/XxhGo9Q6Lh2cm4nemb1WUbWc9OfQdygHA17BxGMkIMVROFjgv8wJi7hZr
4zal+eFdspP5xIovWN5m9DiIVHvQU39mYjhuiYXwVbsS48YiGtfqkeVfpVimUdCPxWbD14ng96Ck
FPnfBfr5ueYmhJP86Jd0zqKZpytkz2U9LrNC7A7uxVTQJyxzwfSCpXF2dYXwG2Dim0dXkppNLa0W
pDAAcb+QmGYjK8Wr0pmCX79XBNWaK2LJKWIVpuTNs6zjjK9QTnhKRvQ1ZyZ/kNRDxUHNrIS1sWZe
3DRdRyJm2OToRHYXjaEM+4NP0+e2UnPyglT+DmNGC+jdtaYyFzfYq0r/7Hp8fwjcnkAYBseewqk2
yZEfqIEZMzez2chHFxFGU1BadSiFDcmGFK8RB4MMbtPqA+4I6GwyMnZAOw1SupOLMGvWrYidQ7/a
mPC3pLAbe1hAqskZSLdD/s4tSR59geZelxkFcEmcjStCuoyuBkAfFctnXnhy2k5DsaG95OpMOsUg
t0JTUYvBn0Hhm8biKBQ47LAKEkSbBakaPeTba5CJkBc+FMNf8vrxKDvp2RMnt+8xxumkwqgrQs6Q
JjQNIjiUGC2lFMUOfNDji35oFw1S+1xgKuc7Fd35SR9kdRNkBpcn6dXBzQ806UKmitJkVuBNF20k
RV2kv/GzXYwDNmSyotPNzvu765Cy3fabeHfgr1GKX6JU03kepJE8FdbM4oGmtzln2rvIYdLdwrhk
Hhk0Y8TdYvnyQfF5kDekCdI0q5qPjj3MJifoEJIWHQkw+Xo/2tZ7J4OKWHBPn14kKFi2O7TEsn9P
jGaL7iHxSZsMnuXt9LdakJwqKsCudI6dBwIsYmP12tc4p53D0MlGwEz2nIhDOI7Mhh+P1rmlxoQ6
WQZpZPKsXVSnOX2jzl0Ko4lvQCrlt2DQBoukZmm9Ti8ULDlXxh9D6fpCvzQClCn0ih7OvyapIazW
4WWvX49S4UnSQDoPp0MDo+NbAdPFKfj7nW6VJeScCePaTIV1i4wS1/cbwmwrKLsGtkIHusR0xeA7
F4hp7mOg7ij0q0DS1Xl6Fz6WKECkhMwmI5DX8keH2b6OoKxpDcPynE5FuewGIqO7yL1Cu4YvYQNM
PmQy317e99VaX3zYEXFGfcRIHvTZfUuEFPbdEBhxDCsCDPQdWBIio5IfK4eo83M5hA/zyY7ka0iC
60GhaiP+v3M8dfi2BTNFGlTcJ+uuNYaTZYIn1B88N2mJM15NqK8Wgv04DWz2hK5HR13nKubFGihN
njkZYV+Hk/Oe+QXU+dyu0oisWS+fYFGPqAnksfB+dA5YLEd27+scjV58n3Zc9bj6cqaEpfgxnVJ6
uZ6PI85ad7gSqHFQw5SrfRk8wbj9rceo5hwA4g8wFx7QBZANKB8xh6zVTkvpPUE+xhc58K6ADrdc
U3bzhVwyv9oWebkCtAunj921OtAM53Ank68HTY7HIuowUdg3aK5WkmCzhWdeVKNK74aUmRFVY5mL
/rlkTI+F16MC8RQIEVxjmG9VgH8PL8nAQRs13wClR+SARITRyrcyAlA1y7c0xraedArhuiWsE8xo
8qYK1mLZoGhWwJ1JMrUJawq7PGAPKePurdVqRaX7QZ07N+7rK4UCSflWEH5QuecqKjrS+AOp6Akf
jq0d3oA6fIJDT+rjZJViKcenffTQYNF0wQXRzA/bMIkYU0e0OHKDMItP3scevP0TvtT/g6AvHv9l
Lil0Xj9MAEj9Tj17zHSEo5YkEkRtt1P3aIBl+5z6HsHbXvs6XeHcC1gvN7ErLCPtcbpuf0E/68Fm
vRu6PnLAK10FHb2fciqFMjf5VAvrrwLqYy4PcT6fWYH+0qm1mjkeY1P/aX2em/IZ+F9w2zGtqtsT
/DxpSWtWvkFSht7B1JirpFCAVYNWoaa12rrrp7ShPnAeYJyCmJUDYbT0NbXMLFGNKIX7ivt+pKZG
C/BUOj+4QcsyA0OGVtW8wCUZUCyWVLZMDmV5ojJnMAXgAydEOAVaqqU7gu0gLFxggvdxUb4UnySW
5teaQ2S/IKmo241wAjugXRhrM+oMdUF4TOdNs8hRetCs0KCHWnTZXNQVu7WSkLSUcuZmFUPwH/X1
KC2h5zd9PfOMy2arJjdzTRaMc1PDlWabE0uaMYiZUn0LqLVp2Xs1rJ/Xoxu4KideLCP+SJjJoCPZ
nj6YNgXFgypu9Gp1O+i08fNb88m/gv/IIfZ7MqKY5KbXAURwj7zEERfuEcQgduJNMclHt6pBAI6Y
5Ca5gMD2K0kpkYEBl/gWOeg4/pL/rrgRSQazAsCJBeNg3Bk0hUA7Kf1yTLrnQIZ0s/5qbgRjrUfw
s/qf2GvLAHzkbEqS3Zi6Oos8bSeb+2LcnDP8i0ePFs3OscBURlNqdmkSl2BkG3phKN+4mK6RjNbm
cfXdy2ih3an9AJBzcC4nS0LoOPmw/GwcYSVCMqhcFrmW9KCqhEwtbn3OqHs8HxN/dFKkQUi3osUU
/GNg71PPxQ40lAy66tEO6AstPh0TamLz/U8L/kvuFLRgFjQd1rvgW7B3E8b5Sx7pyY8+I6LyU1/Q
xp0HPzjVT+aYl8mrT8dxhCb8FTQGFJcpIqluqiRaBpjzaTkHgpmgrgNp28ohEi5tj7zScXbrisgn
RDsmnvtOuvGJlOsn5lLQETK4DuREMxwJDMgSmJsoBZxsDyeb1TtTAnCsYZCKEWE8CyACH977EhKI
BnjnXg292UbnMqNtMTzRUXMevwIICVt4rpuk70BvpZ9Hc4RGR5B4GwOUrxAslJdmmX8SRg23sG9U
ETwKTh10SH059ZqOq8WgHBirdgHr+/2IcG0xScVgthdI8quSAYlw43TyHVwshxJh0sr5Wv0WSW2W
FaKGDhtOEAuloAyd1JN//i3vZ37G7lYwW2OzcNbcT4lvzgujv/6HtNBgS8/8kwOi7JbBmnpCbR55
JC2EcsQZgnVsn+kpLaZftd8VIZPu53mQsCjGoEOQk6/RiBnQCe5DPUaZiJ13pdyzqR29ufdllQZQ
fX38Tj06MKThvyD/Q5U4kh+Fs5xEo2LZcBPcNHnlyJgwpSkruHRVf9nZP992qY9oXJbIUK3Y9Z2d
fukZB0aUJMPS1KEZ3UKHjV8kRFCjQ/esvjPvFV5W0nySlBpxNGIOaoh4X3Q7uJdOdMoA/ontz8Wa
wW8B63FatYclu5jJNWrvRzfvbqeNyDP2UkoyWpDjpUzrWsuHDVotSe1PNCidKu8RkWpheaOuSLgL
4fQI91Ti8mItxzdWOtLQwNn3COZF9e48vGnns2RGCK6TppZWdFj9jX+fv1Qkmxwv2z1tZPyrFLKP
foPIhTzecgg1S+EzvYIkjAxCnJ90+gWvt3Eo4tb2pCYWrVyGWEJFkQ93Wy7a+1cEIFCd74F5/3aR
65ZMWptm0mzg60fw6Bz1NZGQZlz+vs1BukMoaoiYgcg5cR8OzxxzY4dfuNUxY3Sy6bo+nTpyL8ZF
bwjVL9VFefYr50J90RMsgA+PwINWDTPrbjvFWC7OoLN7a83iBbcLzOtiV3QBrQOstPmBLvsaaeJA
eTfkDT66R3GNBQz0L2cz+aYgJKVRhTjxPjru6zrQ3uSIbfLeybaCjhJSJ6uDa3cGvf+/vrBfKnKr
YWpAfOBfDTdF3FcgEx9IeId2p75LLk5wS5LEW++9BY4uMv6emKCThafxhFU+uYgHkCjdi83IgKH7
FCbuIoGSK5ldO3Wfpq2oWw3nAK17/0gm8p5nAfSR42UiYcIXR1VY5pFMLx40nYFOCYXAPUyMfpAx
XTdY0viEt59YbEnFXBFyjN+UDwP1iGO4vBXJPyQRZfSWV55ZyN0N01CkhFrQiBLradqDbH5IPhxr
T2Bu/F0Zu2B7xAzQtrtiGDLB1UPenqLpR5NcrkYerNgdEa/BWWJ1Fj/4UO82oKLet6Qhcm6un7BB
jawz+YHGDkmVy5ZeidF22yuMZhtvMpAWst9huS5DslmBaRJcS+NwutWcCja12JJf0Qa8GBzmOCUq
IlETKNwfzeQPEdBBuVE7wkZdaU0qZvY6/OydwosOgvC5INCspaw92YU9lnAS3Nzioqd3rqqvsYgA
M536I+GWptdj0P69wmlNsj9++CpoeygNvgXphfs07C0OZhocPqVK/3nNSJRWAcwVEum24RnuDENb
u7/yrGdvew38NSsv0xOp6USnUncrmRHwJlVwLZT9q3xspY5IxAYj9IZCUMahpKu7AOyCNz+ehYIK
QqtF1xHEOpo6mVorV/gi+knChscnfW7J3wPpZqwHzDlq42nCrc/Es6lKT+8VqJYdM4UBLBIPDp+4
sipMLhL0sVekp6KL0Nre1Iu5nL1C/YURv7vg7rm8cT505M9RDXCXqXUY5ASSjuZ1Rql7gZhk/xQb
NV5rIQk1iJEvlhvaVe4kfd6MY+n8hqRTiySbigy0Iue6dR8qcSms6OIRkNAb3Ouq3avPfEKWWe8H
ajo2nMEzEUyfUEk1wu91vRwKQjz0FEBc/GJCYSdBh5er/spE/1wCLTVmkvHaZEbPlXDfAdCiXJRu
h6tAlB4TjQ2w3QrihmjaQ/WTBr28P9E9fPQQAQAAjtWZaSjwTl9i/s8H2/gUnaG9NpqaKEv5x47Z
dc5KcEW3K+eJixODHuf1vyWWRNb0o6NojTDBgeYotIQbX3UQB0tnBIYHCqnV40kyRjfGttrDQ50c
eLMSofbHGfyUoNxq7iiTuUrvnlCVsqOT4NfreWbAiE8ZiWeMuXM4idDcofQixLROD+QeUekaKYqK
+8RdZDCjS+h+M0R3PG/dioRADALkzLWIctWQxKH+Bz8sO76Irh4KtEO5dDoooBd1XSdb1SOcYSrO
EFuEe7eKuOHmuBo7CHmq70Qz1rsLtiPelD4Q9LiEo2mgcQXNp6W+xdb26W6l++AAdJs4c3zJuHC1
yjU58nts/U107QAaR6i68su6+vaeoEuWgS39RSKDbs/IX0mxm7vsm2qtVbnXEPguiA1EkGtoa3+/
Cds0CBkUvt20lx7vXofKeVN4TiNVLRrC9u7tVNYnyB5hidqesQfggF/ucuZSv1YOGvhMxBrwAAXc
EGjJsMbOtwFibpzd3x0559PEaHR/GbRbFoZWBzADKfQs2cL5/pZSB5DKPW7LOaG4/SW9ks0am0Gr
ZFlcvPFDhw8AFzHakXHQBQKwm9Z95xpJYl8EdNsZx5X1yXb/OJN1a39BIgzDe2uMpaTZqVRbFDqF
5Mu0RYe5/98XhOs9VyKx/tqcsdVLfa+qpo1DDsieT1azJcAB+ULbbOXMmjWC4HIZB89ffroZ2WE0
Kog9hJn7ktBImf7ubAke7BDUefyJlURZMKSNeQ4wH6pe8+SQcBXhY4isaKS4qnTjsF/DzBrGsXh3
XfkN7+lEtfxgnkHb2L7Nb4pGG1ZhA5O3EocDfp0t15Jtu1SAigD62PYygw3CpFmT7LLAsK+7amYg
rgRVNKRpOMyASIpsL3HBY5oJPihTpuzFYRV9HKC9KqQb8INWDo94YvwzkkE8FuBSgpDTaAUkORZi
jO107MzDTZz4NZvh0+u8XG3HBERewPdvsOygi33jmH28m7d6dIW0gS4eM8Q19erO1Pax9ypPTsIX
sRH9bhaRt7+a5e4A31ghl7OEGhwLGRSvnKGmYTly2Z+HSIfrt8ou7vXZNbjdKPo1O2XWD+AzYhtv
y4OdU1xaC21dx0dN06J5Zgf8QPe3vZcoyqX+kNaGqDWyzmLZTEUTuASosb+2ugItMuLPLOx/Yn23
9RAugPtItkC296cQ2yyHfX6Kz0hqMrxTDZG2EIvpAb9wmEGmV6ZTMc8MU2ZKVIrsbqAEuff34sBA
zXDc9uOjHTro7SeLg5aTZU6keysW8SRQ+82V4vQWOdWaQqZx50QykHb6seAiF6h38qmdaPUOXYLP
z8bUO0ZxGtCrtd79x6NbXTNyosNtlovMHCGTifAWpab93sRHRpLSEXQkg0icR0xRlySBWGsgnTQm
AEse5sAxti6Me9xAN/SbZN+CWcz4D1Ko9JZ2LcB5IC7NNNsZQrfHaPd7qmH0Tvp6E+sQQh3VQ/MQ
/XeBy73a/cY5DdfITyHZCvzyUqm31BO4s/5po179bbtK4YT5vND1GaIa+wrykgrz80pej+K9J0b3
YJqVYuK9grBU9gn+jOHaMv6UpTQhEJJmv8aWgac26Vw4XPIGxRdwRJlIGIlTB7Dpkr/Vd4xmvaaf
jCr2ZzcKSb4cHm23pFTf76ut0QRLRi0lG+3Mzl09faOtAduicIyAuUJqCi7RYzSijLVX4XK4R+yP
swzX/wflTXXxAOxeCLtQLo4+Gbr+d6NxaW6ZdRK27oL7yyGJsMiAXC4T6NEAcZRyZUwSZpQY7AT+
hTbDdJoCKlHIgPs+JsaOQ7GL0Rk9W+3qs1iKZIBvvQYWRTJvGJ2YQLt8gKn279y8WS88whPh043i
3wKnDb2+pjDRYU5bAWq4IMx2kB1Glaj1UHx/uQ1uyydgQgMegrks3COH8wulyp0/XRNBMavu4bkn
HzmETuN7DgBEiXzcetZyB+RYni3vNvM+a2bFtHC5kjELZjzxdM45J9nm6X+gujlMJq5kQjSxRIju
DLPCthdwS99CZbqo0ukqVXy09l+C2su48WdglLsWSftWAhvpk765udYicS2Y0q9RZkILH3LVcH7p
5kxdjRvBEmF74BX5jI1E/Z5frqUAQTQREiAe1b4Yx9ZCBJLSdOMJ896N2TLzTst/I7TyG1ure174
Zqu+m5IdJXVga+M5zumNacXXD7LMZpXTGocB1oR0XbhJ0NIFhzQsC2U3Mn2a3pTQpPkGIzcA8myb
b2rW/oU9nJm8QZ/cH0w6ltCW5yCkmwGmEce8R8G8MHvyax3lZC9mEfeXPl1L6h4v+WVM4plYscww
G5Tv+bGfxlQ/BYZAjcLCIe/fcFRyJJElei4J2sMLGdieH/71GLAoEW76kSopGSTuD7JSKS1YzaR9
+OIYoonTS8R9xXW7oJFyyK881wXFJfKduCtNH52VKqxBS1X6kcrmlTy/UHA+VvhFLB7amNLmqgQg
2wciCAtsWexr765PnnVQ4zB0CSxGw9WyeeONJX7BKIDE9Mkiuz+WjNAIFh+OKrFngsMR0z6wP2ro
aG7Ar6BzafwAIJkaU0vnxRkNakoP9LMeVBmmlErKd9yY5x5ms47nTECTgSBFowPMZh9ZW8l/T7cR
+5Fu532SfKdtYn9LB0+b7t1cIu2vrFQTyVHqx0V7/iPsNe9Mxb3zb8e8f+D43aSa/UACavHCTPWc
ZS1s38o5ms6y6aT2a8i12dp25x5hSsXgi5Hvr2IjGQzjOFba1iPrNFvaZk9ARYatM5PoE9nK3gGm
3ivMwsupmfZe2YOsiiPnd06gwuYu9E18y5tED5D4XvdNqv/megdkhs7Jp8rdfbSjBxvCF+QDp+II
9604F1Ni3U8V/KjMEmX901T3NxnJNKXGYDYWxf7TIac+Osb5Zw0tUb4wP92MEL+1qKo9TxqShwbl
Mt3iUJBzLeCFdoXwoS+iNpID77NBMXyJHgfEHR12ANB3yrLA2fWlS8tJTXJfGsMV9fzBhEs6lwbZ
8otqWEFQgLVWxo81nlg5ulWsN9fAYwgGQiR7oM395dPdCcgVQwYERPYBAwmicT77mTl/KaxERb1j
Gi5XlgRPs4FWK0bV7BT6l1mDXDQGcrDIYgAqe+/4OqXQly8SRAQC/RCEQS6vfohKbvOreWEKOAqU
BFvQCB/UV16JJVjnAqSC8SqWuMB4kYLmOXpAQ25ehqE00EuiejtM8RwqVS7Ckmj3G3H6a/lJ9Pp/
cBk1Q1G53zCk8mUvSpmnXjyPjulOslDyxsS0N73pqaNiYlR8ggDcLcH/rTiOba7nJoRP8V1L3aCh
FNbEXe+dih2VS5Sm/Tle9Tps1Kn0gf8TkYOucPMmse7TYpjc0zqI6rLdgLZmOEao1zZzgXLCzU4t
QRmp9c4BmvrJ4SIK5AqGVAmbO4xBzSY1zXAj3UbO0gbz0bGb5egq8zqNdu7Sd+oIJUR+KBwv8z4x
Dd+1AX4YOlcq7rCjRu2O0OKJ8f87Ja/BsO296OPNDhVtrcBjp2H5K+fx506yHxVHzkjzRU8lyiyo
Lw8Y3+Gi6B05HNc1O2qVWmNGEAsEyryx83RFxhGa4RsNhBtoZLSHZWWrrb36YQZbz+SjYCIkG+QU
yuByNfyWK+sBFGhrk0fh4/a0/3D16lpKu7jrQd0dgJgbiICu17RFz/F7dNqNf7y1xc/U6ssCphQ1
kqNK+BTy4IRu31wWZnWA7jKqKkwlSTd90aW3I3zo5033FnkOwvHPrF91f0GyfDUsg1ISpkLtpDGy
vDMPsbGrCvQK1uFgFB8gdkxKiA9RT3adZZ1mAsd1zigQ/zz04vwilJWMyM4V5YILa8DVQdkuPBgt
ZA6HbhLPGhIrTkKXZJH7lcUabkcPADIFAv0yxHyO2WRk6WRwMnW1YjUDywFqB6BCv38g6KVY2u/S
dLg+zJyZBtKzkthWg6hubWPixsCZKmNkYh6b7poeI+ZL/IAMKCd1HHej/o5bFwwyNvmZPWifEe35
jf48x+HjvQum/KHlXdgLic5gcwS8ytBRO53d9Zzbt4aXWSFNVyFabrh+v0FVLbhKPhiV6I6W9NJi
K8cYZ8BbAJJBd7wyuRLOZ88+arrCHC1eCtbulZjZOOiv7SWyAhpKZYE3Da20S+JdsAcOjeNd+KxF
QzXkGTlN9JEDIPPS9nUvlfjkFPm8Ln5r0QC1I4RnemWp376P8OIwkuBySd1SbyxwkxOdMO3ZSX91
ZCFPb1gPToN/Sle4O/R3zIbMAX4WVjatqEwtVoEUQn4DOKvRHy0ekTNNf4DbBT5T7DUOL8cRVzc2
8QB2tk28zhokQKyUh1DBFzMa2QvmcSRykcxX7KXQsBA2wRHRhx+erobOhKXD7bY07nAbvcJDjkhe
rKjmPVuBDjDPLn0jY0HpTCkvKfe4XyKmlX2vHWdju+eOhiAGvHKdSbZ50S2kqIUb9wnHP1hH0+AC
70e/HPf1vIeDHb/jPfxU5buNb8ADwvzL2qZPRd9B79E09Kv+pphGqwkCCqte3Ik9I6zJT4O5AiXJ
8/2A+suBBQmuC8OwF72lr1GrOlTyusRHDYPBD/XZ3lDahYtTwUqV4wSzJO34jAjkHeKdhxrAOwpw
PkY7sIXrXksbdb1PP9Iu6BqnSnsQpanPu5/OmdgflrCeN8Oiq/LCERPTfhmAhugTNccu214W4QSb
pJ1WS16qQlVl5nmU5MQQRCVrXc4FE1eBymuxwSJybZzW2YV60yPy84iR6c6ByStsaXS+TUn0jDkf
twDfMdJxe592PyhcQYSZLW0BVVmFNAwItacJYCJ1wN1lhsiX7Nsi52JFOtbn6xLng7/eSNWNWuvC
9NfWI0zl+eMLQbljD7bAZo9Z3LlEuCBh0FKDv+w007cwEnbYviOIDfxidkBFLGQNWDa0lZ9s5KLd
HW1eoyVEL18fKG8Wvuxc6D7pWyekz8Wj9M1dtMpOhGEhPxvGtK4cJLVjsmUSk8J7GoIn3tHRC1iT
mhbSf5aK1AtTvYBdvwCfZ8wtOCgmsCiZtGaiSuKzStAlm77ZrZoqgsXWtY7BdtOFLgUN1YDx0kc8
XLYnWSEk6IYC6soFvO1Evoa5fsWJd1E44anv0N0ecaKHjJoMlYfNDXqYIkMMktGIh8n0GAZQTY4y
UpxLTI38UKjfaQs1zIdTIAPDdvSbpj/zMLOc7UEjyS9dC3R4qa6RTXw7mGzHSEIDgmtqMGp5CmFR
+tWoCzEbjrFCOiyxHdVrPWO2imjomHH0x4X9dbxYdD8goL9ptC6JG6IpWgKYfRut6RDdRalbKLbq
WPY8dUcWhIFXfZx3qntY7kSLDchHwsp+TsvqmLjuut8nAD9I1sqCe4J/ZXnv/WMld9Aw13Ult33s
Ao8x5gBOaQPnpCleuSJxp/BZJQVUqXKglhA0hyVRdtTllo1MbN1S3yHlxIJAJhWMz2KWLdzcqCJp
k71as/mf7p2xsJNGUs/pLT7qAEDRdl6Gigh6Ie/viaEZbrIGrpmfwfAVt68QEp3nae+MfABsid1X
snn9/SeUf5j8ezb7J5BflA1BuSHilbimAnl1KrJ++tTvIWUXnyPw/LMG2S9UqluasSJy9/Nf5b3D
cel9KgUmuWUFInxR2B4Oo6c4iY83okSjxTB2INkbvVowow3Xou6iXM7hJ3eUAG4/HxvRQ/YSv/Oi
kQ8WBMqjI7iGt/trOPfD/KvAQkS4hZ6/4L9y/xM+GlWHb/D5O6gqef2tdxRPJQ9ianW9d5fXt6YA
lVNUlvCBD2/+iSs4y/wvu5ZtVbNUQGwMWiwpmjqhEjgwmL/ei973m5CqOJ2Sp4CuVea76wKlw226
zglyI5BhAwcoSTV6aoi/31ymfzM/fuZXbob4IzmPtzmwT5XB13l7Q0bVnTtX3zAec9ILqsjzijHA
yttB8p7zHsPRkbb8E+2rTogHHT6HcsiiwB5H8cUXExdxTfN6ti8+6pmRqOSgRTlmm8fzuwP7oWEr
TnPdVim4CwWX9iCO/EP4U1e2v5GviXoQ+Tm8LrGZRpZVMxqYo3yPVDoBUxehRffwJ1ku/uGw0SFA
OSU9kaTqYZloEs5QImv9qJPg6gRige1MhLC2+LTEeagnQcxqonmcKLSm9zjge6cZlltpExk9LLeJ
Vdp9CN6cFtl1yjhWVsrH3/UbbMtrNxexlsXUYxW9QKwqupahETYqb7UCmLijsE03pqFr3jk5KdUI
IVbvV9oQlQHNej9Mvu5lCp/uQyZktmldMPil2sHk8MC9lNmrbAPkCw5Df9w6OaAKYorZ+2RBKJJ7
LXihyVw1rgsCUBk8pFJc7iauB5vz3l57RGmjC69eFvvgdcmEEKpQh40PDB/AjQGMbmvmkY0ZssES
JrbzKHuC9DGOdb5yKmQ8UDN34l1kaDBH1v8gPpU1j9s0XpzXvvSBkMBf146EPXuXWW3ElXMW5JIn
W9cI8T4Afx/UhfedXY2srt1KRyZmI3Ky2XlXWmDczcBbiEa7rDKhoJ0FR4IF2hyE+8l8EXlYTdxU
j6TcSTVNZP7TYjYUnbHa1pixWdwbMwHscW4oeR6eyG/J8hd1v/UKRyn+8eNSvDqi5jTAznY33ypj
J0wPeHm9AV9OfakvVlrDQ29WWbWoBYReaAL3qPskARpe7L4eYBGFspsjNXZPRVotg31cvYtHoN8X
x0dYiANXdDpb6pue4kFke51P9OnVAvBM4Cj5WIHjK/+CbPv8gkg2AyKxq7UvgrfEGF1CZu7ZwuH7
sAQK6KkB6jr+QfXnlymx3h/fyPFdMnxNBNTpzRQ0ab8NRiESD7SjFWVgbLoiEUK167jDjbL2h0fS
RsywnTjphOncCBlLEMaCFbgcK4iQAqptohfmq6m/kRJ8Xxwql3ZpOREfSdDKT1lLEw+W3gpwZHj6
l4/1jd20kIrySlrqdSgoMr5WTrduhsNeKk7W++ttWyfjuWlbrxHgR/Qv6cV0Pjcihf+yqyFGFLue
koRSOOBWxvkTQIOkzHocrfdfjA8hgtyjku5RRxwFKySWuqwmVV81UfQJEEMZNa2+3qYxW1Uuxyox
1dp99tS2URLkSx5XuwUdXB+0wzGn9HkcnrLieFDd3Pe8GmXbL2qkxtKcvbacUVlm3agcDrMnAeW5
T2RqSjYNeZZCPF7o7e9XVKnYMCdy1S1BIHNLG9NP6WuJT7B48ZtHJZ8A57r+Qa6m3qdfTFER3Ii3
2h1S/0spT5LmFJ4DKJa+2PUplB7odTBSHXx9LDBKqPTmOHlhUXzXzsAoxJDqODAvn48FeA3MhYgu
x883uHTABLSMEKNPRPkCqVdUQbM+x0aybgaVxj2xd/+V1yn8GFDI8IDdgb9JmPGDa1pEWBbN4A1X
2baTCAuV3HyOgFteSmMHma2D91l6ZBc/HduAKHenRbrr5kbzIK/OHSkdOP1Lsi4mijFh8kc/bbpG
snM8Uvz1QvaNb5Q1kiztADp16+hrceNPYvmFC2etpKiJ1sCN01uG2sZK2qiEg5h6ZWv3E54/LEr1
JmVJkTZRiwgPlSZo+dds4vr/8rDTKLY1QEXXse+AIbUbzzBQDDQDUikTEO5deFs57Obih2gWwueY
ptGnfzrrpFwWhd85nG6HyIaXVtNkcXD8dlxBn7MEYKSW4x9QB7X0pftuAHWuZBNGUBwHGXa1wwL8
Mh4zDY4iiBMt/vtNk+2t5fs7QwS6N5cCAY4uxUqeOdbYRaC6CETFwdNlOYUO6LvCAC0lZTbrkdn8
LYGqBllvyZ8V39tRpchrfIatXUtKLYBtT9i4PdxtKx30dZUHMrt7JFkRTAUqEnUteokPXDMTYTqs
8gQZaWP5szBNnTBdQaQxhrV8OmdmZNc2nekTFmVdnMxQoOn2AN0BDEmVSC/i/7tLhJ1Qmo52lIZH
PEQD4aIQYul7UJLCjv4uqNxrYTQ0ZfVMtxeu1733S9le/QOlU/2+f6jr4SBlkbOs7U+DTY4En0z3
w+aEY/KFyRfr6r0ZL2GNKDr1LIW6fb913exVCvA3GZRR790DklRl1coI5IACWum6veZi74EmI/Bi
hxvuyNy7n+O0JhXJO38wf10sbsrShQ4pntIbnkiGCJhV1BqpdUmmKl8dubQxYBvd5TvNAIm7lbWS
nL+sRIbJTlcQbClNQcW2liWA/g41jlBTDpzmf1YNmG7U3qjdv/JRA0y7YE64gwOZXwC+EPjA69j5
pSAUAqgACMVireKZZL6Pl7RT0skgjo+LeLUeHCNKKAa24ZXu60bfh4t0LR4pLdoHkR0XqeDjal0i
NwTQhh73vMA6pMwD1yAxM5fFer598YxCJJTYc/F2zQU9F5FFJeMW0dajJEGdNdYk1tF8SuF/9Se9
Rh4zWJ6YaOuzs7pi7ll3SYIfB0L5Gp+XbQlVADnn7RzloMZTEU0RcTZwYaDAqwqhSQXWr34QaLkx
IVF4zP8+tkE5yaUHP+tOQoXLdBwj90VeoYMROv8Pr6BKJKOIceVjwfCbTavC7HpXe3jM8SaSuIVi
e9Ep3zV/nAoEYAS39cnk/aA/jLDr/qbxvhTNoZU04EkgXwD9MJHyZtWFRqRmekEFyw17TfD4fFNg
nCVFkXYby64bKPJKyStv5hQHEviZEY2I0KyiZgCK1ba5L5ZjHkWHt0vkCCx+txu0Iw7wK2ZpbGtl
II4Uhq9hwsOs/E86zk7jt83JCumgYuA9ectpf/gN3IQSIt5SvociJsYL9TbLd77Is5Umr+AZK8iV
QuCogWOvL5ifyLy4a9KrStDP/0S3YgNHQFXEfjTSsbmXATF5xNkKtRpU3lqLm2RNur/e9RdVf9p1
JChE6mdqSqt3gOqAecRwVx3wQ0cHOFY3ofgmNDZ2b0gfcres1PsOVu6QMDlLVbZjr7mJBxzqAx5z
05qVFH2UeR9No8w5OE49jrycbrdsxvSPyfwT2P1GPlsA3V29LRt48bPCcWWni9z2ZCXLsdljZt1J
F8C9CorM8E6axbKLj0pqzZBBe8rMROkBywbLYRpbA+veNxEjRAgY3wUIyjA8ynAeoOQi/TD/jL4X
etA/JWqhck3Nrt1MMZhZatv0MUFY/FoWoG7PbpvgA1QiHMlR3MW4AnoOTmRy4JGOVxjUZyND0oco
ggB21yNF2XifK8QA03Yye4ovdLRxbYD/CF/JLk6BCZa81sysrb6sfY8ukXaXgYLXAoufDIaTu+Zl
DJARzGmKVB7fnPZvDgXV2n3vt2phVIKe3iIc2KNT80mG3Sdz9zP9oBgaQ40kz7Pr7afJPKlVKogF
dTgbHjPTFcW2E3CgPVdVLitxToDQZZdg77dDY19tY0eaOM1tNyusGeycgnVq4p7epvZlI11ArCYD
Ngrvt1lPOQWH+nMBBkmPdrewjfb+2QU7KBrHLQSvZd0sdiAaKkNXu54m5P3LHa5LhKHSV3FbO/iD
Zt2risis1TLLtVy2S/uukx8/RrcRCxEKAZ63jE9JGVkzUmrB3e5eOuDjp5QXJZqdq3CtZdl51l1C
xxNmroJxa7ZLCk5HBb1mS/yCdfr2xMGBbFYeJUk+9vU5kB2xmT4oJ2cwPOmhr7jxOsRhVyYoMyct
UkvtDetM4ZXZuNFh/pWjpv1Z4zqZbm50KPpf95R/LACrt8P+5gvq8uIKZBOMSL6ztmBIsMvcmTR5
l5AUtwRSjc8j9to0kqZG2I6tURx0L2fz8Ta/YIl08zpWxn+r0G+dJGx+xYWNcj6SbpCMi1CVkoHz
FpzzHJkV4KRXJArlTBRO9U+AfstqlAFdf450GUTy1I0LVtQ8W3VJZlKwiTESLCVZ5OLBoObT5e3b
G7IvtM5V/n+zaHhkigxJG/eagjzNxO6QJjrwxK3G5x6QjVgsEP3HgvIfWNrCbqOiGsnbD0MbPUmc
00o2WnjCcKs6io24eaVJj2YDTsz4oG3MjbtfUf0xTm8bhMqPwujTDEbVESx0hDplx03Y/2vbszFH
DWq8eH1Ik4yD2hN6vTYwupqD6bsMK5qJX4w+y0Ifu3ck5dyRsZFm3l20a5alxGC3FaiiaUC1B9Zd
9Aq+jV7vv23Pcg6pizoQw7og0n9vPE7Vz44BB6MSwW+qtqH9d4SHGwTNuv7cDia4P8LrBAgNTvXQ
OIFxNLhrOsahrHrZH2D0/MUXkezmkxDAS8Bc6WoD1TRioi+U0CuiezBpps0y2aVIryMzCWp237wx
Nxv8yUOl/RWjbg29m7Ccu8+3eRB0gs2jq9PPU3XVT/KZVsxtddc9TkOJ8XKUZbSERpnQ0+502RWh
0SAoKgiQXBGEov0yHuhVemvRwLC2IPKoNw69oQ8JSMu2TidqeNSVGLg8CYlbqJdMimaxHmEbPUup
gr/s2eC6njXfUUwBe1kEtBaVTW14z0eNQLtvzlEO+eFlr5DEGL845jk3CldiqNvA7BgiPH5QARuE
g83FWKBau7VQJ08ZmKmU6+W5CxVvY5ttr8Jfa1/ohvp7FqrYG9bPTtV+mqgjTZk/MIoRdEUrZhdm
heY41FbJIKy7kEtv1wsWV3Lziofp578e3hO/R1tvTEZ6B0wwypCFGYnbbA2sGkeheSjt/C0nbk5P
p+9YltwgeyJ253TBt7dHbN6UNCuNcgtJz87q73hAaD07XXTqURiuWrIUOtNb7SqG7eM14+7dcsK5
FZfBbg8cattN5Q9litrUXo8Z+3L2XXf07jfy/vttHVyMA2wAVvAhv5AMH6YUiXgEmf+de8xNwe3i
X6KGTplFkgjLvUkAt3PJyb1AqeHkbwYxiWZElUfDcooe1C0SYDrpUPoWgm4GgW8kMh/avzZ/luCO
BWFQyGEmCcS2urK47Z5zI75zhkbJEXgT6HewffAVAElAs2JaVggI6B7plY4tgUaWBWbvWrs3Q0nJ
FiaLrCH7DhYALl7Nkcd70I0UCe+nDLCjro/5sPj+g3EUjqJmskUBkRHYs3RThW4jgClUhpk2KXdb
O2xkEGNZ8l9yO+WIdgdKuTRuoY+JPA0eLLsYXl+3I8Xg7uhzLgFqH1J1KGS/Wk1fDELV0p5pe9I/
MMGY1iPS6UkvYZWuVBdNAlS0/4K04IN5AVrbsnj0NU1cdCJ4BVLeEZ3VIjTP3AwG11YevKCqzz3K
/zOWhmHBDEFR9TDpwuPHvSOFxrRAql+mlUQA6V/QQdF02LW8UX22pIwnepG6nqZ4uOPzV/qFuZFg
A2r+rEEQnW/Wb1z5nGPJWB+Y3xiOmD8g6sNNs0Td/mbaFn43oXit8ksyL4X8xAKe67tfJoxNHxEc
epCiXM3bt7uXcjJfHEfj2r2nCg0VBEu86F1/fXEndsDl7lURNmxjG5fwwDA/84zx6Wy9eFBbmrxR
M6GJ519QADTFEKBBcEIbNmHZeNwmTr5J/NVxFhO/e/mK6J2/Ld1e0LSlQzNQ7ObgyrJkndRGb5r3
V20i5GqJTeehOjFZ5bBn9kS/t9RU8BtbRAlW6sbR7I4GNhi+FSEffJ/pvkvFyUfSLZCVLQKiVQUr
pGNzdE4ONIAK19nxSl36dZlMzittRNWOo0dQUCAEZqZvAfm067YPBDTBWC9edh/tzusiLFBVL1ev
9XEdGP5tYwl8eJ60MuRxlf1V8qvGhCpiRQQ1E6FIKdF+R/W7p7axGdNLOH5o5fs3wVcvNvGpQxpS
OzRwQ6Ux+mhOPH7mOF3Y+a6Yc71YP8jWUsK+iePMPg8RVr5+st0OEPTdEWx0qEXJMELTYN2u2Kxu
s5p3BAKjx/oU1vkRsDYZ9vA22OfT26jPRjhuyoXTBjP3ID0Zlbjcv70crGVUvW4iAI5BvZFHCP40
RtRK+GcZ4oNqHzzrz1oL3NN8UTAHkk2fTB46Hix6iFtQARIqT8uUt2hO1dm4cNmEUIGfC7Ta/KaB
Fz4wTTfem2lHsv4soHUutTKEV277VEcKSJTktuRuHDqG/ttP6GaHyfQactARC9CrHCoLmZR7Gc7L
UrxmGE6TSNhMBAMyEqD07P2C4tJsLzfxnN/ejSuE4ZqgArEdHv91YCqJDn4hd2hFOKcXg3pitgRn
4MSDDzxZQU/ENgG90+rDw1n/92U7/7dqtqPLakZYhIlhZqAcZ2P+95F++RNRT3M7pvDnZeOaqITR
ou4cYD3pCi1sYRuBcvszu/CGzQlFrJpJVaMGPkmrZFmk0QUN7z5Ncvd6TR/BtgAwbBwOFfPapNoh
FhNHeV0YpKzOG6IapndptQC4i5gugsIuziQa2LpDH+ybJvZN+0QVnmBFPspd1oynuwyAiqfHTv0f
VfczGKqpY0n8k6rEICMQpmLC6GPvSNOQRyiE3SWQy9CvL17RCVKXjUWGZ50kZMRcFmZif1HV3h54
cCrCoLZc4hl7buOP/rOozrL0L8xpDGW0sEmv0tstCALIbhea9hYnEyQT2c+0VO6jMXBV4ZFc4j0A
HTryhohSh4LdZjoPcI35BW06oOeEkHfrdF9OBa2XOTG0Sr4E6P0PM85W5gAqS8kgv4Wn+BnlPIhD
ReSSNw7BAG6ant3DQjOUpuZYM2MX3kH3Mk0Pdr86mraAo+joA1OG9zp009xl3Z0xvcUlPsP5Ek+y
LUkHeCdBJWhR+gDHBXIYOZXd2kBmGdyM2n8pdPz98udVcOmbH6xw45Kce2t3X2fzA3vP/R8WfPwl
ur/E6BvQ3HsPUdSiYyz+hC2VN1+ysJUKrr4mXMfaTN77K/3TaYw9Z2iQTLJMj0sDkwzs2fEjj74f
BgzyiC7XYNLXPeBaPEY+d4XgdX2+PyNjKuqj8tWtbV/+cVB+h5PxnEJ8EBWLWX7RB2/im2j+H7UD
R1P8OzlqJcB65NVkab4XD36Z/orhVconWyyIfN22SlgzdzmSxrEEitBWIUBObxLln2mFk+LywVxL
kRkS9oZp5oHe+NKRtk72JJxGB28Ae2A84JaPZBEMBGSvaDuKeRBNhLnkjPJWoKHBWTsFtiGXa3M6
FJzzEKoV+yEhJGU3bs3AA/JEnqnnFsLyfYfzznkJcHizoB+DhH74wTSsbmjXdN3iguUhsz6mXOKj
TxoCOf9391S/7az7xhr2dOUqgAftQE5YIjT2JTZF9LXkqTBDuFR4N6FoRHWjIHqzzCN3IRPXQP92
A2bfwrGdkbLxtQijeRqKo+ikv66jkpYCnTPYtOF6OrL3QngTbSJkS/p9ol9Yf9UrRgA42C7DvqUe
uFRvWIejelNkQ4ZwUKn6NxJO9rffIHKgKc9Hp+clpUL+uKxmm74Db7f7VQKCf+cOb49ndakoCFD+
orfhEfnORawwtSmcLMgtr179PPVx20QIKTnwr+b4ZLrM5t1yeizJ2KDgSS9hwsW+GdWIIlYoIiLW
a/7PnuP6kHmI2SMgPoyrHPO6K/8jGnTlWnJueihKF2r0pL40UW1nWiWqzv3q6yocNdTbjGmgLStn
D0pMgXbCNcPpkQgi4/nTajcZh2IvSuSQUWw+KpE0N5NoUiEv+zbOkDu/cqE6UC2yjIPeerXJFwxk
951+HwDe2d1bByoMZVhhJfNntuj6U9Y1EDtMza6PiGNsem5Bhjjw6Y7pttkqiL0kxyAcGpLH7pOX
3H2AgYKiVXRSjkwSE8OmeAEfiO/FKk6wxUFa1gk2CR96v5ALPK9/Y/cu+s79mykKZy3pmrdJSYdj
UwDWLxFrvofqvo92IGtcljuZaOVqrmYV/I75pl/0sX/FsvrGCFijjjBznPY45q6VWVSfkC7BrN8u
vn0SYCqz+vi2l/tf/l8nVTW3/yxl8G8k729mUUL4GfxPmoaXV3xmZ7KzJY743EvefxJb9LB55zXO
plX74MZR6XtWpchevcc1wZK5WO/+ukTPPqWGQCogO+UgaOpo3xBG9Uk3YD2l4yd43akHjFFeCQ33
USgTBfRGvrR2UARP1DC/Bcn0+q7BsDDS3Ar9SQoU5yAC2ZIBBTss+AJWG+gW2ApxlEqq2+VQAd8h
V5TgxC6rx24U7rOA5IXgusaYMFUxZVI9moPynNad2lbXGUH53XC+BhJghbGoygOtNVrBm4VJWxn2
RdDDjT7qwT70G7NNqJYA+bDGTV/qYZkMAgWQxDrJVyhcj/3QngmlSD5/1FqKipqd2hyYo5VixQbp
jfrXo5YSDxO1s+Cmsth/a+4A0KlhI4fOQdFzsutdLDpBi9iqYX6RVihFXk/xN7jLPStbdLEGzXYc
NShXNuTPCwhtPfPr2u9Y0uaYv/OPCQYY/w+ytFse0Zq3ck2cJ0qRubozDDVqfX4SJ40FupW2dQE+
gddBenZyyNjJB9o3Epkos6X4kL3xhZ/xI/sOTlmWVofA63siq6vX1Ox6I0Kvngxa38bb6SNwqF5t
k/X7wi/Fy42ad7oEj4Sa/MDDDUNzeBRtz83yNOHKebvPbjMT0gjh4DQQB0SuBCxqdIY8o81fhnKE
m4koBxJzLF1PJqqZNiKpj87AMzIsai9/7dGFmNnJ1N41CSIGXRKZfYxbfenubA/E4FsCcrlJnbJX
9TzJwX7FEfbMgUxM8rmQgpoVDgcLUL6fWshGqGITGl0YnK7SEYNV5URT07jOSWkc4INemSS2Za1V
9PgtXYWWrXhM41zvS8PglR2uFUXYMzBM0JCxgr+vydfcRE2lcH2eXI4uHfBDB2oNgDIz0A8Gqeg+
KKQWMHbYKDNs+KkG+dxvoVyvJ8AfVXVZn3mPaG+azSQqZw89XIonuEnIyj4jbEdraLG3PzyU+HjC
MvNSYhpTRGJrmTXrfj62vm9YA9gupts6c22SDjS02es5jNT1QkqEr2Ysc4M4pwD950evsdrsugCN
R/FhJvHatqF4wXRxasGXZ+pfULij6GNr8jBKwy+egGwJCYlIRHEIFIWDzceno8dX3IqytmnbHoXe
gqlyIZQNoDeh1RT/nBWJXAi7LLCm6zoASrysO3mzmVMPzSQKXK+TVKePlcy5FuyvXUOIgyu+ITFO
vjRESMuVRoWWRfmekcAgY1/54bYTuPQxjQwKAXW5J9Kej/y9JeOySlFFbY+WUmkPqdKXAeXW/Yo3
w/VjQa1AuEhJtc6hhQ1s2eaIfyZiEgIWg7aalkQysy6wiqoA8MVJEkuIcssFL476gRQFJIN971wq
LcIQCAJLPRWLT7JdKr/9FkFYwiSmljCOvKVXzovqonJEVu1Ujvx86D2xPQWIfAMB14r0/JBxGTKd
A92hGQz2IL6O2G1dek+0/sc3If63jhRS2zXt/3fTIX9SakGbg7PPhly3cwZbh3IzuNJeCJQoe5Hw
jQC6XCPVFcLaE9cPK2KZHjKM++hAueTaH2dew15kj/JhMf44s98pKj6/TgU6HNOdFiyulHzyFUBX
+gYYG+2Nm4utmCN2MBAOOolIpaLgW8TYCHA/I/loIR+ULtnPRLmtEHY5xssFST4HzIWEbVMqTj6M
PDhEeEDugUpBlZ87OhXveZybRBhXqgyGw3nZrKCMhENxpez3dV5DE5E+JKqho2eQamN1IMlmz/aA
aReQoMfbDwSTYTp0aSXcjXy+7ceadegVg8CcFDqOmtVUWdl63SDNE2U1lk7sUcyQYWAGk4adhHfA
mTU9/1mKiI5C7tMMUTNFuIdnqS1G7lKP8o9Jxzf2T24GTsDSSPKDCmBWFOFt4SV1/JrcCAL2XRSG
6gseBeoDuEWj4qoR0zEzQcaqzCUISgi8W+5gObfAbO8vVDE2r2PM6dYd0cu3Yj7QPzSNZN9Y/St5
opuO5EaWDkCveG4kXGSWPPgAv8EsKb61UmWRp2G2MDKtlMnq2g3xT1kUhWCJxTOsVNINgm18ToK1
QMHDFsp16wfhc0j9Bstpl98lYI9495mu2V04ocvr2Su/nd8382OmaR+Umq6xX6OhHwB+oQWlM9E6
dXIzRXuN4HAKTYc/TyRhVZ9007VyvTTqRl3r8HWiZghyN17rn4NKSJEED3TdfdRnpjC7FGw9rzSI
w/72r77TNQDihTE5zG6t/Lh+DIV9j1+IEtZAqngpJxRnieNV5Kxe90s4hF7UikGV5GqeTANbJ3ls
LNg1lOm4TUWRPwQtAaShVW3b8FNmlIvDTUvhxNop09E2nMT4QX8hwFE+fpUNHWvjfWvJWTzPTV8H
o3U7vg2ga1OxssCMuM7sMYklhIT+vzPFzZZ4Vpfo8DRkMY9tyGM9PdJ5a2wygxC6kLCoJAY/Ezou
KzrVryxIqt7Iob0D9SlrH/d59Wu8ldMf45LWGOqPBr2VmnOYW/nJaqfnnrobEYvbUbb3LltsHXfS
Qt+sHxaxeTRFE9o4oxlOZ0pOIYyIRE9ALMJ6XVRLQjj3ckKb8RivM/Qwl/JK8AUd/dwiaVysEsvk
5691/G2x/rq0ig5EKjWedQ+ZuMppO6zZ4aNoL1a09VrEkmiSyaGuA+q7bCa/cnzLiWyYwu1I0yti
e/ERzTMY26ndup2Yz3oHbT6CfYqqYZehrUVLHeLsX8xvI2BZmj4+VEtkfzZze4TmsqxnivBBAGMA
Te0dEWSL08IR51ehdCzSxs3EuOAoY/hIsYrY7Rauk6cSDJepPiuXO3SJonTTg51Xty9ijWKEg7gz
tzeiYQBHYxR8Ib+/IUEwVY+vUUfA4jZzZyZb799r2XmjJUIuyj6LLzvamUwjXGkeLsfqJmrlQJyG
GBvbpaz4l75obV8WUImk/DeHp1K1onw+PtIO6DWc34Ta7FkcpBZRimkMJOXOPyazymw8E9Nl1LVe
wNhXoqNhD41NsxYhSDhuA9c19Sb2zX2ACw3AupA3LAszdnw2JmXLQDoGTgrmlnAFhpYLaUsrJydl
QGCsjniFPeC/BtfnItYSNNQ+BJIDJNY/M6UI5YcS/d47V4RCPPjh45Lkt8RcSxCpgNN4i6nPjOPw
4QkCdsEm+e8zwDFGOKl4thgOcaWMWZoajj4mNLlrtaPXUgBjaTWCdVUlUAKHl6OX3JpwzG08F2yn
rTQim6YFP6A3mFcgvijofatBKN3CZLILKtVf+vtdygDSVvpzFF9lKZYOOpDlLrmpt5jcus097UaQ
fFXviluubqMOPdy6nSuXfojfnBFz7s+tFWILw/V4JYKV1Ema9qsdM9Z877P2VNFVA0ScmaEpc23V
EylGfdLErFPY0aXi7MyozLzBoL7Nn6h1NxILX/CQXfPneU6Jf/LwJxlvi7JfMLr3LFAt0dBcye46
hZ53Sm/E1KBETY2FRvh76TLYssnlag70kL50poFTV70U4pcj3kSTB5TTPwi7iN3mF7p8HOX14Izo
MifAVKhs6D/85q6LKKIN2WZyvGoAu6dUPQL0ZNbDp+nsTBGoNbYUskK1DMPSgTVKbchgPFTM1DXh
sCnS+HspA9f3mE72nj18EXF4t2YfAKroEVy4+9Qsy06xVHpHJ8tAwVAFbHKDDor7+iCHIPDRIZ0g
uM0HIIuvwnV+oscNp4il8UVaQfzVBB764tn0iq/OfpYHgru/+FlvKbODcZtIDjorhopQ3D0goklR
KsIazp0KYb5TuHzhtpE1tgm22TwJ42u7M/m6baeOQTivUAMzt0Qt82jyyKyWUE3L1fALB0uj5YRR
2WplwXX2B2HSmsZZtYEI09h1vdUqCMCorLG1zKUjD1eZ8PF+TckHjT5vvBXpzC3fhXmjvU2t4uC4
ttfgdSkdH4fE3Rtw+OCpaLIiMce4eP8AKAL0YYX9AdIQUUpoHXxPX7JE/AjV+Vl8BCNi5Oc4zJda
1PcjIKkcRpxZrPU+/Gn/qk93dpO7Gx5lqyEqOD4C2lFICGrNdib4zOpmW9ZQXlIYVxWfy5TV39iT
P6wFninD34k6uLW5bzcQM8gKuk+BISDUNr17NwFdeC6N+A9G4Lxxp2yjzTvcsBm14q9ybEqpHlIQ
BSlEzEF9M0azMLwDclXNlsajoBumqWbxhNDWkwRLEBFp+aIBnoo1qMIiX+ltYo0CXjPX+LmQJesE
fYcGl3BZF6FakiZib3DkTYtMZ3rro9+ZXdyjdr4bClboht606DyC6axRMfnp3UwOZfoPIE6cfC9P
kak3GdEp27yCDY9SZ7+aFMioBgHhpsji+jY5msz1SNW0XXEcHoWUnLbp01DMbXIe80kdX0U/xoR6
Zlh5TfZhEutdODi3DqaFwcFlWKk6jLCAvRh/c9bsE08Lo0OHlPvKeyZ00fTv61M66YS8hDYpiDCt
+vd1PpMUwz9l69Xq5u8WkKB2iQcpU29ufYAOlgdCoUvzDhieSSK7HSPQLcjoPDMozF/CASfzcstB
4ooZka+sATDus3cu2tbLrsE6H87cBYE2AZu8cVOCZFYuWMzzX6KS5mU6znn/kToCbeJUkVAz9UNJ
BdGg4QUK88ViT7sfMIyI9uKhSmLv2PdMpLss4P+kIEzeEyQFdFfX0FlJtIV6D5sj6iA/69EUysjb
yohtg00euEYkuxm9Bc4QGgkdaK66WwD4XiyigwyLNkqJeHCyAbzEFoEcOzhXBDBcRuYzj48y0f59
ogvJ4pR8uPa6dlq+5OWJjf0Dd002UP7kRUoDTRAQ2gcnEIZQUo8jlp/VOAYOgZsi/aaYhN1mJggU
4Vz5rsdz4SzQfi3KBp5f9mvGqXXQSjEZuQd3+4EOap8goCL30X+oU3ABWakiJ7/fdW8B16ou/Ypo
Pf5XxZUpKoIiF++tmAxJGgtcf5PfwTbQb6BYlutW9gHxKmOUsPONMOafSNNdoHBRl3LEVs1w+nxD
qIpktDL3shLqlnu5KvNcO1GQxgNpUkz2QaUVk680Bdz9QO3jM7oQMs5bZRamV/ycfzHXJOqdEjHd
Ini1Pwzbn0nP8wUx/JjrWtYtdGiAe1XCOhOpIazEtK3JaJqvfP7N9L0V/o3d+8uizpdEF4qXZodu
AjylTVCCSr1CdGSEbYE3IuWt5p5U1xVwxY32dQNJpZiwDgPtpXuml2bq519ZPL1D3k0G7pE5Oc3f
teAtzFmqRfr6Bje9bZZqqK9m3rEJd2687MrjBr9aKUYT4MMd66h8la4CZHBoDhXA4KaEEiXSXDbD
9aVQjB4f5XSBlNXdBQuHWO2nR2avff+08FSpkU77g1DqWA/oXTZlk6teMriaREj+8fHs/Qi4nEEV
CTZcNZ/p1j6Bw8Ga9kXzDGjI6MUh7H3ZOVCmOGLydIjayvooz/X3jrdrDHGCV0fjxDrLDDzVEDfy
+uSUWwCQmz4JRDkhwyorTmGHK40BF/Lg7etA5gj9P1AfaL8X0JliPJ4inYZZqWcgOvroyssSh4CM
X7JPm9MxdJ8gUkpZIs532R2X4fdIl4ISbYwZgHZ8DJeNNhebXuHwMC/0Nm/nXS2S1egm8nK1jFqA
sicvnjpWFF2to2qowN6CYL+CLKqnI97RgsD6bQ2bgOjEOjFiaNLEwBvX9yDAcHf/S0ooSsSSCYId
oClL0ArmhcTzVYSU8Mag1j27rKazNLiG+m/wkrn/CcqMMqA0A9//Sitesm1n/WJZ4E1liIDxMHP6
QOIvyds9rgOQWdFedOs2ZXK6/MzhkeKmWeiZoQU4HbnJqIN+QQ/Cl9sKdEujL0bbYaqrjn+AdNzL
WdsTDDFzN5jlgr5OId2JANQB2MfZ9u68XBMXcx87DAGRmoPzgHhO5kI5ZTVyeYLKLB7zU+GFGuo2
aRhUlqcu6PNlerp3EycpKREYKftxwrf1Obop/vCpblTVdE88sTwi+Q0GSzbKbw6SwfXvqbn4bow9
IRbNU4X9ER5S5+aQXaRAPLLAZ+4pe8cKTg6qh6ubmTbyFMH3wqax7ca0saZTO3EQLQub3nnOwK3o
sJHhx2fDevVP2GLhUS9pZOIHHzRzWjdVuWlF7A0CK0trSkVQYhO12Fjt/SXVaZonMQfmk3WjXe4i
rb7uovr4wXD+C157KtuNtkuWkwui4JdBLwRuMUqjoLIvt64VHNjVu7ZPLxhnv06RVNvZrO7f7GQa
4DJ2BJ2FLTgquzfWsuOnUlo14kF8PsefGn49MCfkjtOcBsckiyZYqKD9s53NznercNm21D6xF5tN
WuffIYovJ4tHFbMd/DPnrOy/Qb2t8/btNrtWDraDfxo57cxCL89Hg2dOG6LRX/dQCQmQPTJ+fOUj
dbwvP6ijdf2P3pKoj3EQDy8zMug7YyespiucaEZ/RpWuVCVnrP3PBWdLHxWMgy02k3TBA1EmO81e
UvEECwoA1L/EPCoSYEBFGrT0B6ynT6t1g4IYWndCttPRBuzPxBoRG27TnFFcw9q7c0ht4s+kSSKG
PKnCfc3TMxVCNfbF/BidXXZ6BWyLqVyCDXKoQJNmND2qE6atV6BbpL+vhSEVxj3CVs9RZyeU5Aa9
udrQuxZEb4JEng1O8u/I7XjpOEz+dtXO2r5dcGj1ikLNkLk6kgpNmIf3qc5tgvhC+X+AxArJEXXa
6kDmuW5JWVbA4sERSwNJtAK+3S8CrKuiH12G1wXho3pcuszGKxMmU0+f8GirMiqUlJA2eRXPY4es
hLIp/j9kEnuabBvcHhTy4aTyiJ3UaM3YNetvCBP2J8JZKhNIb27H+xl9JcI1A4xpGkqHGIFSlyik
33EDIUwiGukAX0ym8FJ3KFC3QXKt69zQhoktcoBjOibDrGwKMOO9Y9vpUMuU2NtNPEETC83YKebW
zmoy8UDO/ZpcJQaF0+ltTAlgXEGwKXxeX08aelWz68wRHU2JPMVZ498CBmtGLVH/l9qjUVYz633N
JNsno/9ygN0E3ff4vWk13B8K4848tFJh3XgVOX1qoQ0UHpC/0J8xxf5mAn3SADJmmMY9U7ztZxZY
yciASCeLccAY59IOVYcmYSbHAdO2HWR8i2+dnveqEvGatf0iwL7yzRELvHT1DtRPduybn9qsmHDR
w1mAyfjP9O7y9k5GZYJ/WzkKTmqQRwrr+6TcBI/uhsB1bcfIRBR/ImtAseCNj/esYZXV/cbFpstC
Tk1wqGMta7m7wM7wH+ZiWnpFr7/GyNCzfEOLWxAZZzHPbkTGf2l3EKUaHNytpT1qxCfEOmjn3xTA
LK7ywn2WmYC2D2G+vPUmkzW+9KsvpxRJ1yhCWqizgfEr6xKrY52aXcnnStwRMUxbYf5gaJjYhIY6
YURyowi6FytlFf+RzZDrQ2K7iCctMI2rKL+TQpkR4UtwjAHG8O+qHKz1vO5D4LMgUJH/zHYenIfI
1X7tkR67QvxOB6Ry7cQMITPcMvUqSULIP56NNQQDIpRBX38Rnl8xcaxDvLVMK4yxAsMoUaycdGes
3UAc1VKgvUpI69eKBYvGafi7Tcqks3J18RlI5erQC6BduJzhEEWHae5LXZskoAJdeYobMs+r7Bb+
rw5xuFabENZxRXp/t3JIJF0xcBG6SURpaO0ECM/ToB24ywTYCu9bdZVxrcsEm2Jp66R+y1h6WVJV
lqN0Opc/cWUsJcrmRQqHjaBKOCQWcwDP8RMBIjTIEMMUHSILo5TkdSZnyx2WDfw2jAneI9fCt8lN
lOmdPAUzcj4VqMfBucG9KBUdEaK+SEzaSQ5JC1B2n67vlcCCECpkL1++ZB26Ds0+QiJMSaGTtV19
P7rsshaFA6iUOsc0P1DieR1xEGVgsoek5g9GpWzIM5rSdt7jtCkU6TmonHZRInm3jEdFsiW2CTrU
6O8rBcrnUbBrZ15buujHvN2A1H8r/N1gIX56JCGBgFPQV1iD4u73yZwoZF/z0gm2ICJk9RImM9aO
McStaHku1Erz8BWiH+lqFGs1u6opWWatelBdkUBMWpM66QlvRLE+n9z5V9JVQzbXIQUf7QlQAqFG
Cd9cpDoI9H3bi4/Jl4hxhr8NTlYoDvdByHILzjfA5FcX137H2VmCtMaL5mHQNv/x2GblRGfDMU09
U1VbknpT+v/iM/UYuZ+35JPxzYSXcg5KQ1ajccj++yjU2rlzBmCx9CYAECMo9fHNi4NEaPbHheYM
8akcaJ+KDPFdIdlSJ1Bh3gr1qpXNnnA6BbWpcI+iv+GPQpgOWD+lIVUD3V+dt6OFASqXrW+qHTSw
/vsQiREKbhJ5Yi2fylUaX2YLmvPqp19gCacNLbFsZsaKmJHS0fZIw3jerp8w0ClFi507hsMEY3Gh
L4MP+i1Gu1mJ5ETABjpcpVKnMyI7EG0Cz4fQivFqZEh5JLSK83zzM4l7FX3rONem7UnVFBXSq8Qq
uLrIlLuAf3IOLslrwXruLOx7zuMcXweQ4LJQxkTHypWhcrl7rcD2uBK3cq9ddWUdPCjHe4Io1smk
gTS/9aTG+u/o1Q3mTKR9IB4IwKoRLtk+SUWP386UYNCKvrcDtBI6GxBb63JCDzPX3OC9LmZ8kYt3
sPyFQNVyv0r76j+E0HDAivUpX0r1uy9oyrKPP57ReGLYMXKcunFxUckUr7I3USAk0A47URPsbqL2
RX0Q+UQYSk0XVWR5cA358r7yeKx3vqXr+iLtEEJVYktzrZKzKuDPto+Pmk7b3rWMTbD4317Gxy9H
ZKFVHm653yCOMFFOouYwzwiUr8wfXhxq29fMQJQ4pXSs1+QnC8IOatu+VYYTW+ug4HWEKeCCfar5
g4+P1FQLc58nVG5+U7z1wb83I683NOFj/0QiPOfufLEWdfhFw8XEB2DhATR9oqk8OfEV2gGumQ4a
2Oqo8TWkKHb6r5jEPE1ZiXi/mEAdltmeBTl5P57MDCi59IUAE6Z4mrEUulmduEz2J0oKtGrLayoO
eCecEJTCfJw/HllQF+QG/T5EkKtsbA7woi0zfLRatqeP1ARdKf9iooi2bGLOlS5FTSk4XMG2NXP5
OiY4IEHOHEQ1wYHwkPGi2jXGLIJjQON5pbI2NrFpB4A8cbTi/tEjweSIoCUb6Q1KxYbpDKZp5wWF
ZZDoOGplb0dJFXCYSrelvQIso9+tN1+LQh0HflidGNGS1T6rsrFBdYBj5moD7ehYcBre4aO6kss4
1Yh050Kf38SkcDtv4jyTonD6R51w6AeBfujGma1d/EyhNXiqW8LbCufumKjgpX+L1DGyM2V5Giz2
HU1Y1EvlonQqTNNBxDHL4fGPTwxQiJ+Q76L6LbNnZ7GZ+5256q2k23JED8OeNhHdEWEqc7pjywiX
mjkYao/3JsUjJZviJazCi+0aMZzlPPVUIFIkZH0HmuVqlD1eJHYUXgiwSAGeJ+gkwXh6uC1gtW58
RNNemdg+t2Tc9CAqGk2b8j/zbtysxGO4vhxi5Y+jrgqff3rAeYlaThkaYp4pPCpSonk9vMWHpSbV
/B9afpoczN8eUqHWoM8XVa8kUgdyEArsP3Q+HDekWw7+yrYz0epa+Bl5Z2fcgrgyoqJo/X8ZQlag
ZocuYmUGMbSXgqBISYRA5X83+ZoOmNc6MItuxQ/Q9J2FzsYFeM225wmRpzCwBhpEq1nst/WARZvg
8idvH4+OQMIiAwC0+tBmDcTS8iLBFXuSfJ+2Vcqb1AI94UXHxNuK7Q8NTmxs696VrnAi0oz9pJbW
KiFl3ndoaWB+oOlYdZQ9w22Z08YGt9lpd2chzPyzyK2i1ZdDSydWE8I0IVK0N1nE/pLm36M8yIGt
RuBzT9BLuspVAQK/vEfhShNgniW34bTwl2GUNru7CMVd1AG3Pbwx4QCIwkA7jfJG9Pm4t1u83d54
yNjiL+6ihduFM9n3MxJC4QTqU9/OhJF2NaufEaVapaMS+42NL4J5Xp6h2Zi9UA0+CV3BZqLwQZoH
Y+rsxwnTW60/SjzKh/L+T1yG/nYWkjAzFSZGxsRi/j8dEijfW/2Un3X6iExXf8ReUhE3Q0IV+IXA
PONii5LE8tpqA1xtjgcp7wYMczsxZYUBYLfEVfUyejUjBreOAfSxjWioghPF6dXOSuruKjQT5UQw
B8V/E29Szdxytga3LSFQJhSjgEkhfNGmXuITel+qRYk+LQlzDDP3XgR1upgyL8/R3p8rImyFJ5LF
2FSZOl549fSvO82Ad+vxNk+GR7SMK99uVOrMrD9UU2CQiejGkjiOYNa9z01Bv1xgQmBC4R3o72L6
MlpzS7LXp7FozFnIq6MGo29tLTWwrcXDsmSdZVcKkLlexQ2Fy3GmZzO8+NxxcFA+drniI9YqDQ+n
c91L/mQeVpv+NQ8vUYxTW0GpRdi1EqpNgTFtXejB1AcQNtEyPHUk3G0PCraPPSHahgY9xsdDFhrd
yJ84xNb6ZzG8duG6k/3iHqHZdhLkK6CeTAK45PJhGZkS6AGIv3JY1028OcrNNuzWS7epYu3Crahr
jFwYkwqry7JqyZh/AaREi/NTsQ7t+wNcoeLthOTBJu5orfMoa2ab/m4wsRa6Sdd+lQqf5ELS+nPF
9lyvzlJGt/GPOM+O6jN2VwBlH3HrFh8p/VPzHmn3HrYWr8dLPxJhC+sST34LiJCWv/0dp/PHUGVl
VI+FHfTOhenbU0kYEzSCtxO26NktoYraQl6B6Qbiww0q4mjeK1n1owL+9UnJqHp37uIk1UxdGOKQ
n0WUwyh8Nkbtfj55jji2SH6F6N2aPeRiqJ2IDEV/7i0G2QQMzbrG2oNQWHxZTwpk3BBijvjyhoEb
hXB1G2m5lcgxNvOJDuF0u79IClv9k/cxAEigD2armJPmGcs6ahdIWv5RAy3tAz4mVOH1TqTeZUx1
FI9ulrMFzlkZpQ34gFXcX3ASZnu6i8PMNIhDrH/DzcTUsOHrwqeO5XwsWCCTVSzOV6W9K3SxiTsA
rS9DGcTO7w1NvOLKJ3N6PDsjcF2sHBG1Chl87i+zUFPXbdLCx/kJ26HhMT/MWVMhhkuTT5YZKiCH
nO3GHW4tFt58p75SEBQW+c6dA0xxshogjZlf5fTfOVQ4aj/JMuXUoaO4os5R80phSBU28FUqDnu4
erxsx2+F47Zgkp4iHDTvh9jkYRHPP0BEsZPLwrDJkEVcLdDxyyV97tFszbj+dfOr04cghpVInWj7
HpCqx70ntqJishaEVJhYNnznre75SzutqBf9ydag+srUk9MvqLqnjlyQeNTNpS/MPgr8G/dgzZmR
RUmUfsyuYSxgs9tWSuDyA4lQKitOuSBW6JvljWJkVnXOvBujXGsPWvX5Ye8mcqY+/MKDNaET8HKt
Y70n/oYCqJQUR4saHzRGSCLZa3Poa7kMEPpXPrKgKpGq4iGliok6G7A1BpNJljxT1IUjD9Dltrh9
0fMm7ZHwgb5k+JOE/WhxS8YWdrwWVeBRXLz3L6vnlV5tkt59wmss03YVi6JNqrqlBWB6j6Xugp/g
rTETKSCYkFHtbgxG/bcr2EC1jCurS3P2kd+wyxQVz+6dzouSQXC7FUHK1tXf36M/t2zW880QGWUt
ZEklg25G1gY17xwesIxU+4kAcdXpGSTBstSscMqz0GzNebP/H49C/4Ybu+KTtPZcjw5nz9RfcKMJ
Ti6xgRIua9vC2EvkxTw0ehEYL4yIOVyvSo3mtg9Ds2vpUIuDbxBbE6GmK2iWdlU9I6NLL5xAXm+3
O1+uVnL5FjlRhMHmdS4C+Wewf/XBekl0n8lWMT9kP9zVqsFhOUI2EoYj24mcazdgOhEGe7CRJ+In
2Zw+oMzs0h3RFgB51ZlF2EoIWx6EVo8k0x7uFcv25t7SbEb5u1UFKLO0XF5cwaB99163bBMn+VBM
a+GpPG4svnVerXbs/KZ3TLShq/v210ddjD7/o1gYhtF8sf1bkgfnttxtemJ+dnDX1r5RYHPe28lp
WT0rOHF2W+CFs/b9CI0RZDDY8ZTAchAIZp4fEXxhw9Lb4M8KtMmttHc8kYnt0r9syiJUlpUVOXO7
xlbprHyBEUD5B7g6T9XLjDiGysN6tJPzp1a2fkv8hdq+I1RTnBSA2geTXnIhoUCrFuq/LU6SLAwP
oSEcjY45ecZU8nxcdcW2Sm7PCnKRHbYj3x7oX4VvmGZ8mQzrL6yamTHHQpaMX3p4jIjLx4OVnhPv
s+N9eWE3sav74SYdUGjGtrdFZcQPJ/7AULCDJtKK/SUHoH+JoZTey6OtI8I+OFrbs2j2LeVvPuWq
JJINbV2uZlvpeq/hW5/OI4UFdwPj8k9fo279+eVQ9d/WIskVsSH3abv22V+63N8d+ChSb5Nlnjv9
eQ9E1b18IC+M2WZ/7vgMEkob14vTKR7hXyrV7NQVeupH9QWShlcsCetVkQKva1MC6U87pL4jmHD/
OBQ6iMShfS34jsUVgdAhmqK6/JvrEhc5hU7teEMSZ+kiT75kgiHcTn2cSM47tF8HVOKOdm3G09bO
RJKr98Rd6O2ESOpbMx5xjmm1thD35iPzv6H2gUcS6JH7tJ+0aCUTYtY0LGuyF4Mt4jMQcxJ+hMJT
fZCRMGDeG0fyl+HAhzq+iYRbqsGOL8EO5bmbmxOmZj5EF3gX3dA84euzIKKkeq4QWini82bZo6wm
QbAf+n3jjPTLAkdQMZIyMjkgBzgjfjzi4Nylek70ri3FRtcQ/MnORV+nLQJnE27mbuS0GKIfgQIK
OKT6ErjPN22VKb1fcy8gm8P+H5MwW1H6PYDYPXlHNmmJflvF3ardmQ7NBnctmkTubJ3ODGkMVTdJ
SBBfYjufW+JRxH3S4D0pGeNNoGwVF3DkPkug3BSRExqkvq6udENME5RwX5oDkAFGaOyFETyi8Cvm
xXjB/XSmiIy8gBo346MmT1jzF0w3U3IG6ntzHRkUjHXFdEV6MYAGGvMtn5tn08zqUayTRbHhHK9W
LqV0LL88kwZ16yuoQ5ho1lDId5vm5lX071YDyFmU+Ak+lbSjwlL4nOvVFbUZ3gUAnoRrLggtWe8b
8j0TAOG7SmcB4wQ7XNqih21JqhPcNonv+Bxw+E0aC5eAXIr2QSNzav0XuIQUPl0V0xAqWe0CPJ3P
FePQszmkjSrR1mFgL5zuj31WVxee6Cjs0YxGY/6AaP6DiditG6crvG6VJYbGvonnBuFsrriSJCl8
jMZmubqpra3w5vLt+QeMzwymqkQvMJWzJomin6yJRN8SCMp0mfUFpa3aXaFKAgUoTy6gti84pUzL
eAcOaFQJ71ZjnVudukxNwF3UiENrpsG5d0kDDcurf1zlKWL6qyb8JtmXlZpG6j9WptA628vVOsVN
8ToeYzpfJcDRSEEZtQOGznW+ICFlr6rsp/H9RlLOGuJV1+m35VI6c42HyMwlsgrl1V1Ojyu/Chhv
033lPNyi4TjrnZdwPBEFa7qyoQ8AZtgWal6sb7tmJtD5+ee6pn/3znJwptQ5xHl7iNY/cIpOchNm
NBcQUehx7Yc9cGEOJ7RlVtJlDiISxPsllszRQOqelMwT2YpOQHSZFhHprZPZkA5ltofwNwMlFwHE
k+ChxFkzx7xYYnMNH2ZKO97ttgTlm+belEUTXMCwbv1MDLkRG2f3rksp6DQS+tTUkbj72T7HDO/F
vtf0Qdkvfr1tsbwKRYzig13uLz018nF1SDZPP0KKyebWB8M4dOTH08cr7nA4CwzQ3AgHKycSE9oA
JBghBUywkeEQIfFxx+lAj4rxXBR6tFtQzKXwb0YsGD0PfThONII6N2+jnVcpOY4J43Hb+RCZ8+zp
Aj0g/as5Dm8UiWyAZoo3TIOihOM//JX2SRi0K3hKa6LT+eHnb1eo6HN/vXlyzRtYjKzQetpVyQZJ
H0UKHMo+GYSqtGYvSiywOj9OhtkmxPANLDsZMZuy6oPfxPFietBIffp4K9Cu1/7VIc2eAlvz3EPb
VYTxag8v4sZYxMEejThG+ORPw0sG8mkcL67+FkkjjGHRkhKUioheBmdB28Jv9iA2IXDnpIM6X0X5
514Az2YCPUyf2pI1WfgNhgFyiLkludCGKejzz82/a2CnfaCKLx/YzMQAo+snzd7aH2qnel69Fybr
UI0DwtVJtppI6GnMRnQT9zzQzkLtble21keCajWLrUOR53HsryigSDUFvO4S382fpm+RQcN6l8pa
7oaEsTtSl1ts0pZjSa70zV2fYw+EWga2+JWM9so/0OPH2c08UR6Jz9CjWNlnBWwZ8gufkqUvDLqE
260L7Y6org9SuldCGVEv9Jw0Zp8WUc3o/MaoKnZX99dJRE2wpfGbtxOLpC7OFsrOVx7as/xjN2RH
fsZdXbXhP3fZsKyT34v1q1EIkSAJH/lOiOYn4Ojox21N2oj5u7h6Zk3FJzOK2GbWL/9fhMOHAVBr
Z/nlcFpxOKcBxshhG5B9XCiGL1mLaUE6HTG6t0TIkrCFeu5uP5rXlKJMSJuLFGr3HrwNWxYR5d3i
cfC7wuYvQUu6snY7QRlQx8epEz4k77jQ7QdahJMSKYkR7npwMrkxnTFyaKgjCDm/WzLLnUySFxGW
cGhtUdne9dgi+B04TZWD4WQZETzSYqpsy4LdnISAUWf5jPcfLtqLMbwau8/qreB3vQ3MPSLF/15+
kYHSivKenJZM+UTYHGn16QoWB2WBA5yGBqdmfC3/RcmAeZcShwpKo8XiG9tthQZyxcQ/yr466lWi
RimTSgHEe/nmgRdMSXSu37X9c6ZcbWWe/003xHLOOLP+kl45Vt0WxIniZ0dbiJqHXjcNXYmAHwMg
ScNKKvKSIovGyUzj4IF/Vvs5lGBrTZgKoyIlU4UHrmaXzwA7nolzQJAory2KZZ6kB7G6MfV+ffJe
73w0hjdsleqiv9nmbSfzugb3eHhe0+t1A0jAMeaMwiL7s6BfJ1wZzkWkiNcy5VNefG4fzF39M/si
SwbVgeP7YqJWxPxAmJlYanaMuJRjJcuOaRPJYeAKnYcz60mhgSXb6t9+HDpRxvWn4GUoiSko3GcA
d7ipEgYpaT4Ff3O/u0Oiq/2tlk4m+BWNskrfS3W7SbXlNmIT9wC98pv1XbAb1z7FyqgT5erd8yhn
jSc2sHhAybb2SqfyIUGaMz/01MPGaiHDQrPKF/zlk0kHhudR7es/VMePoBtI8RXszqYi9Eow3NK9
iCanRHM1yu15CZpO2XcEo0VHHAAdU7f4tSEWw8xwTB1xOaIwmGdgCq1exZKXp6ntHO93OTjC/+nK
v+ovHYKa/9z99KSco6XSfOECkNPE5wr44DBgy57nHJsWns6JDJ8Pqd5fyXLB0xb0p5G13k/l9tkd
FMuqT4+Yd51lrA5RVWQLc2axsaoM1JS1UyK9e3EKSfp9sp2bx6uCsTF2V16TpodCoqQbhk0c6JQI
ymvhIpFSSpSFvZXygjZXuyILJwftTxwwBpUkGAjW5+Py8JjhyrLrJZJGP0AhxZ6KE7YJQp3DG95F
f3kbAWlWsedy9hp9uwcazEF0DTw5NHMu0j3/DQs+2hBD8npvEtpxVCZg49X5YZ5geTDW/vDdcS1q
Q1ObtocTy/6ReQYsaBBD5IKfP/qLXv9vIUStCk2/bJvofsPKCIOqZoOg1ZEbhiL3EWrubVxWaPWm
05rpLftIfmIBOUoMj0tzOnIKm8O4HjeCCqo3kn/kCMAESnHFoivswsmXqRYQvaNXzhygLo7YA547
1tRQSrJqwHbxp9tJaavBc85GO5XG0yLrCZfUqb3vfet2Jm9Gm7JwtKYPEH2ZhFyvwS6tx0arTbxm
OKAxfVbqzPDCTLjfrnxSE8W++GJbRMcekKbCNgY3gqZoKWznBGnhS45A62sqzn0qBwh31PrIX6nF
ygFslqY6v+lqfOHYdtMoys1A7oDdsHXVMVicocHKPKd4cGe/4LG5fCOzOLvebBBrW2vLVWtS5CGD
bewPXZL9ypvRzg0YjRDRN2Gy8VTMSVvVq9w6JzuS394XqFex+NmKnSa9pNWdFgthTx4tmaSri1oi
YkvDtSOZGEwEDjv0op5oZ9KajyXb5UMorUU10o0ufOvwf36+mIfHLDGHfAVevjUA/RJ9UF2ss+xL
9XRo20rMBKijnnCUX53KrCa4VZ09Sb41agfeTsHB70leWqufxTSOtT5nuvhS9FhgRajIckrLDyhK
NrYZI6Bk91jCDOVsPLSV5A8Uzk8dbTBN8bGcOMVxfVItrFh/AV4137OIP+/lahlsvokiTsNv4UUv
47E9GCrTAue0+3HVNnRKnQC/ka2vy4zmTOpAryFV9+uO5CEJkveSjMAp/Lq/2fPktAqeyCHL0mmX
+2UOqAhdKlbrWvfcVrY0RA8s3IswEOinFTw/dUkZR1Vjf/M/9H1lP3N3y3a7q+muvPWC3hjND4nS
7f74NouJh2ZJVU5/HG/6Ib59dF8iVHKuBf3YPHM9CpbR3uvK1R1ZEBJ0u/oRkOpnv//qEUVtj5dB
BXMmoBRIBvEvDiL+/2RXniNl9w0Bq73pLFzrKxH5XjgYczaTu5+Yj7M6TL047NjKZvqUva45U/Ie
fv569eVHAYnubmoAW9ClMnP5TBJ6lNDWfMWR9zxoFhdfIVciQDKiBDhdTGUsyEFGV5WODogiJaMG
dWP8KBPSUX5nFdz+O3DUeFyOitNxIh/HWi9oBs5ebxaVYYi6WzqIz0ynUAbwVNAGFwRPiNDX6o46
vy/YnHcico0PupRtSExI2ns8P/SaYJEABnHzxtPibU2c8Hloq0viBJ+STn169QfGv7mIjDR8F/BB
+HHbLJTQ3oy+9QZOpwlULJHyhqMnUkhLJ1zfVvFLNhEgAnZeFQ0WmBrk+n1YT8YL1Xm2DzMTbamz
Qx7exe+sL1YfYsisRY5z7N7txYSNmDwqfWbqP/NubzxkiBhywuff9NexxVtOc350MB3ERGxxZVfS
/cK51GsfhFNvby0JoIACTprfvQ5StHqi2UcFBWauvhVH3cKeDzNnW7ACzOKh1p8obLjioJNS9FK1
0jqRnMtaN4we5h5l4sY9LkuRfSHEwdTJDAd/pIeoMcni50u/L/c0OEWwkuq9mKHym/SqG7mg7HQx
hPRAK6LlMAK0hllutqtw+r/NthIS5IztuLAhhYRwGRLLrzNS6WG15FQ2wjXFzDUBWAmk3m+12Olm
8bXD2RfhXMbRqf1adYdy7IdOIIm3cDvT5w0zNL5KxwPSKwXK/pRI9b9jb4pA9h4popENIlfiLmig
FlxroVCsnIo4n3iBqMGtkaCdX7rs4xp/6SnYOqF74P4f5GKKtrhPLGX5WBYE9Yg/ahUU7uA8tj6x
8xIJRIzUs0yXYsoFiL+8XTorEPKX4lAxucuXoLfzSDfYj7uG72AtU/UZ8gJOiUB0KDD2Lh8SpKdS
fOIYozfmTzN98djblUzyVjzWrsecBO87tJ/9tFxNy5JREo2woaevcNcdS2p5vqu9KfzrIILlqdJ5
AfZdUfVB+1wuY9O3TgJAx9I2wRNf9UKOYjz9W7d3Ym9GtK0CNst54rwVythMUlzAGdGe3UR7FECL
78V2COzEQTxhBwYGvrMKgY6GB8AcKl+QqL9exAxus3jxy3XTfFyzh0PRyf/u6LJEs3+9h/GreTX2
f76i+IWUvn0ajfG6ADQrtKTyKVuUpIL+j16NJ97GH0BVbG0pd/1bu3MP+GTiSUQDKkssHCjE8rCm
3ie7JOHUEmjv6DRbbf0a7ESJNFOMBXUWqfkzK7nVqGQDWhD6q7wtDCtmLtHFc4O+E64ZccOMUO3o
oDzMJIQP/YEW83QMdmUOrRBUgvFe4HnTkCOFJAEvtwPzaJYsgnicugn+RWT0x+YIKijzC0381rmB
cwa742Pnfn9B78+jBmjYoD+VFa4OaxXiQX5VFWOZ50nSvxR9qiVDSNHdegkUbzduEzwgp4F0CD6W
LnAu5pPs120tjmDeSjf0t7y0cyOAWFFJNvGtrHqJGXizPSfsrbjmzKg43+sZZC70pmebo/ZyT1sD
JcQDkkIShx62m3Fj52epar/mbxXQdlmc2bge7PIS9K3fgHPMCublm/QM4C5WfJw/kMGlsbAt7ch3
dKzUhnedsvsHH5QeBTc2nBybS2IpEkiawdlOg7E7Nt2kr8vu/lJuN496h6ikpm14TaCjMAyBG05I
XpTWmmMon4jTWvNiOvVNIwEIj+niHdwh/9wGatWcN9LwBKGySuP+4kklAn2oHWW1kzVbELUsb2Ux
huE6FeQ4R/HVI99DvaxhIpXyV7m2Q4sLbmgB9icdPK/2DbTWnXsLEqv4vjcoIdrDJG/Z5so2Byfk
BKUR2EYUk1EJTFWDGo4vsSBBwZnMSQ3SGsQC0NJUcu57rw6pn3nZz1JVEUvaePLc7XkksRet4sQW
vv1SMw7d52NU76mCDnHzxN6UYgM+1eRLpGcA1t87u/a24WweLE68ausETilojwv//Ty+FFfjxRLO
7XJOTqF6YMgnGIW4V1V3yCLK4ldqxYmwIvf98uEIXkEldV2TRnP5Jjj2Dxf2eUuCogCftG1B+cf8
gEqyOIfsUzEodGU/HjcCZVyqIn/F/nEDtqPAiNHBFfMJFC7Hf/mUwv7mzskWQkrhj0TNRLbVYyqN
9vf1TfD0mtPkmIuZ7hVbonu4hEfZ8yl4vkNtzR8HDv24KlwKaDOObopWC1MP3Ki2GM433UTHuZ2z
BE8cKvsPKVDis4dpcsm2eympwlLZHYfEIJwMM9eYNIdi+OLo6zsUi0V7E4oHU8mPy3/sny83+GK2
GBu8nd4JiHP2L2klVnxD1MmV+b3Ywdrk+EAoUn35gLGnEBWE8BuoX8FsjVpLwJ/70+TCLq7hjmwY
zmlvit6voF//KKKeauA57WNdC/fzpEV/VSghau1xjh+Cd4cNqixnaibMj7qj6lWcna9m0E2xY2Pr
E1JJ+JpT9Gv4CYDCUdqQC5uWeuTKD4UlNNOtnTWil3Fcz+6cVmjnimyr0Wi6PgRgfolSFLrn7TDg
hWPgrl5qcZUSC1xTFbAegrZv6/L1Zf4luCmlHXkpBttCsD5t70xM8fLlHT+ayvQpc4u+o+W1qLGP
1gl3fe3FDt9ZUSkGQt3+zfV+oPufUf+n2/uWRk843/c8dkYmQjfUXQkY6j9UiU5rAoa3um9V0uzT
AP43T/+67T3G+sap6UASrjL0Ok9qjqjBaYFN5lfWng7LexbkIDPJ4fVhljFCCx+iZi+QFx/4cOZt
+IoXPwJIEbV8urtfMQP53bUJmlRlsVW0jMZ85Wd1w80VrcNobxyWHOaZo91ehZ5MA95CdlTjYVNu
OLT+gS1kfEe4RpU1iPNXturQ0jxgZ1Mbfxp8R8QZJuGuOyc3yQeWlStWY71/6gDtekAiYi0K5HzB
1ySAFG1ej5XpmpN/22WLMYA9bHTzUs7Z+F+QLX2A6AWWfHgr4kBZjqvGuxzEe8TB1ZmlGF8JRgEr
hLIOMTy6PFsjYEFGIspG5JWURXEBiw/D5xatwEIvkqLKsfZJW7ItgJu5+qkzqs3EBIAaTftutqxA
lHzlpHZp3iw5c6qfrfVKsTaWUBTWqLR55wy50keWNBRXbjiZL5MBKubUGod8eMmVm6I/9bC5Xr4e
rNQgqut4S4OkIVlOSXuJ7kIgw6TaUaWf9h9qkRrydJ9HSJ8OKdeDbNZC/bMSR79eNFDVAS7RyAGR
+y1FB7eZpVrg2Q9eeyjQq2hKGoTNHJpibTPOz74PqKWRNqtmA03gKtIz5STCDxu2ie9OWyR62XHB
pCYxdcG7UxD5fFAel7u1kojnWsDdvdcApLR9CnpqKabaTAaTfekdpReJORdQdXnzyNALYc6vl5Cp
M23ZoCSCnVMU2Zb+hhtCzs69BQfoEzBA2sTxY1gYgsLbbwxBXPwdZ4+V6vz4/z9xeNR2Javd/pNU
W7k1IdNXOd9Zcwk2Bhak9MFxogmTp/57xP9ZYpSZ5GUnqiQ6p8pXjbuM5Yo6bB09dQbudTQ+ecMX
VhEitOrHkPtN1lAdYlUdIP4h3LOf+hiQX7yW+f85LHVXchL95AHPy6sehfBuBr8i84/4ezIAwgyl
4woYTAd5/M56WKgIGGqb4BjVBS0MCw3bBZ9m7Kumywv+EjyPNJWNZXjPcYdJn4xvn/8ohHDiMYsC
7gOheEiWh5d/hb8BYOD/Pn3HUCWdxpmfToY2vyM9z6e0nY8p7+1i9gY5BxQCxPGcOIo/qDYigzkw
LL0qCN3BNqw/RduY/6c89WhWhP9w98E1J2ChNB1sgUYyZMPMSPffgoQXiBBAECkHmrwO2xPOgG7r
fJ1CZFoRvRWK5EmjzhmHfvtv7w5xEefQI60Fmt1wJFMbklJcfvWvhoEpQpPflRsFqCl/6fXqBFiw
AE/a9p2FhefvRQe4wg7jVZKOFwBA24X0iECmC97wg2fxLlDw4QIN9qFPG6Lc5s9FumhS7H5TYFpN
p7aW0V6fc/viuNoT2k6aA/rQ6cP/oZm7nLmVrrUuNUmrxN38+Tg3iOCGFpP5s0+TmWSfMyLiMlyl
sORie7eqoLOwvPdhUtCtLApGc3IzIon1LJlJM6VYoFyVS2D8M0Ut8wo9jSjlzhNLUYcEiAZKgPBy
r9e95QN4ku3BKG5iPX3uVioYk6+Lf0TsurZJJwfLrpYLQ5he3gWnWy1cXpCmDSBuWEZkRGeiwbUY
CRaC2fHcOJ2VsLfSZZqr/JtyZsVPoVIYEK7jR7DsUX0K4zvI5C5AqpMZOFwpT2jrA0O8O3RnCdnS
RVPuITZQ7MbBx0csQo6eV2kRe7ukQvHsXQEnAnMDdCz2uirjLaUNucRv5NizDx/v2KER4Hyh07Vr
e27WmY70Y0jLbJ7X4y0frmPiWMqEnWEkJs2qHJ7cLZfRCDwpLhNWKSKnZfFJkQerSs12IeUs4+j8
lSRY6kEQzmbrG6ZXcpCFkYWC01phB7ZKVxVJrQBYN1NW1yvAZDh2tW7Z7MaCGoDTdTd7YQoXfds6
UNNJE/T8qcF+UgWa3Kji0Ss2nMc7zdKO9T5qnAxFAUjGg5ZJwYPuAZCf2SZIFpYq0o9RMJmtvTEZ
nqH7BR5y5iSoD1tfoC2lfqkEIKzmGJX+gmUZ9xOlUOmU1rK46zJGk3zQ6zuhS9Z6vtQQYvNnmDCC
9/R/yzN0ISqqcinZ/WH2HpAOkfAyKkQoevI0LFG7g3cIc0Bg0Yf8EjpT2CAw2k/GpzQrWKf948/D
FSAHbv7o/JrG3UVmfDD1jo8/W4vVFFt8fXd6TRs82tjOJIA0fMxTbSm1vDDF1r/W3COb68X8pLhx
SW4FuOAWOXeISdkEV4YespAiDk0byvGfMpFByuPlLnhhP1t5s0NP6fKnhD/ZbegDdtUuU/UhXBKu
Qu0DsVfSV4ad5umo5Vgc8/HDj6Ow4VFKgSQ4Zs7Vx23K6tI3Da81mKPgtkifod0wI2eZxMtEkjM8
FR3QKKowlw/hV2ByUi8o3FRTbYVGtFNzrvVTVF1cuffwgPt/sdduDIPQZMvfRB6X5nGJhfPEbOwJ
7alklTURHERNpc0oWllhgWjL63cX1H1Wq2RTEQBfCe3qqFp4a2IcX2qhSABtKLni6zVMOOHLeg2q
Ua6DiraAiJAPROgucehOmiFpksunYex8uz0P4DQFFLOxEI47NUkN+qBvQSc2pDaq62pGfZNy6xpy
gSrCChSHUTaQ2xEZny08vT4bL0B4dh4FeSwpcQ6RroEXlVxHExHB3z6jPisez/mOjxqJJoGik+ck
gzt3PkulPmyzucevFCYAeYqBV7BXyf2kNoKQz+1pxGjwzLk8ppJMbMDQJ37D6ANN8EIp1u0dJA63
fLeEGjrD/n+xM+pEqP9TCn069imKOSf7Jx4OnZEH65usHMXGs+g22WmTrC4Qd8k+6UU8eQB4PT0d
ny+6T+xHHzQ/28a+g1fO57RmXe8U5ndvhQsr5QRR8VAHv0lOYWLPCpfxQx2IfB51ry67WxdPmmYO
aJuqdubQ+oJ1nty4G84G5OMgG9sc4wxVVH5sIdsbVmRynY4r2T7A7u6v9HB2NFpwoo7LVTh30nFb
wJfYPTiZY/r1mrak3z9V1oj2rYtjhIQEepFU8TINPtRKAGP9yWEUSbALTBB/aeq6+pzvdOqjjNFf
jpr/M210myqZcAUnH6LWbmKpuKY1UVdx3ilQNXO09hdRWaLfz6wG2TzzBm980TZ8a0517+dE4hGk
ODrQr+yh/u9WtjE4t/FjWw2kCu9UpO8X0A23lmIz83WAIwTf5KLFMooqnJk28fEy80k1g0CcOmDc
sO5dyIWCN93XX1c+PDYIxxgMawuUBsd6ae41MVq+nU5Yvb/ApL47OcKovwTGdI2uUGLy72U7J8BI
G8PWckDyNpf1vCO545ig8l/yVbKwcLSo6R0OuZFQWGJPQNdTYbBe6Xwvhm+oqqlydgTxD5vLcOid
JPuQIOkqbVpOS19axiFuxhpH6yxBlwZpsKhguq4OaZmSEUzgOpvOzbPC9/yeRiXcKtcadI1MRqvg
7Ysbq8QhPEYzM+TaaSzHCnDJSyC8/4gjChXJtYUiE+qyMMEMD7qxb/P27Xwr5l+FG9FqIhoSQW1m
SruDTkOY5JwRjPfci3Gu2k1vO5zmblfkVmDuXQ3PDp1Kefxo1h2jroRkYPEom+PC04yD8K/V+wcS
0fjy5rLfN4XTdOSO+5e1BIP3MiEC8ohA3ezJJWTIoKQaV4fRmxiYplUnRL/6uuzRUO8v5Y5h5QYE
CjsbJUEWtse4wxJzymyhDDcVIIa3i0tr0VS6ej2ZgaQfl0qx3/q0fCEQaAafFaMke8ylHGbtIMEM
32gIqNF5AK7QIvNwFZR/ZsR/acXiLePL6lOLR05ROGdwQccBkDJH105WPZNHSKwMSLOCkcpwkuZt
pTfU7kG/n2eCmVSeYSYo5mSlxWCeAFy3fz2cP0iEvIREeeRJ2HL38uSzd1nWGEM6oIfk4sp3sRYD
1T3HWGyUH6ujNSjhVvhZnDVy0mCUrZgJuKv1NlC65HF0wVGZiuI997/4OwWqertQCPr6edV+BL0T
pO/8mISd4bAHl/w+O/LJFEWcLwNiXbT4+V9XE5IRP/8glKkarQn2janU7sX93KGNcMS/Xayg+n+x
4PwXNgBEV7mYdSsDORQM21kddEgAlCLewfAjuG66QYMIkG3rPpARHvR4O+La8Gd8YmxhHzPBeACp
3i8vL1VzjbDhtWCPZn9AyiDMyt3FqJNZh6GnsSlwPNEP9r/DuNB77csCFiakF//PBePq7JyIQkSO
a2vynwf6/KLxsbui2nk7NyIayODfGOmCh56kaxneE/6WUofCGkQoS6xfCXG0zlfTwCB2PllDEfvv
OM8yjYpflwtbQZkT1N1/oTIevgY5JM5R9awa6jEj2GfzjrzPvq+OQlhx4nCvSgufrDhE/ckDe9JZ
W3heGXy/nxEQkwg4hQG0JRjXKaPApmn9uUVidRbbmBAUr/MHlXT1Z+raP2vHoC0tkrpo0WPcGH0y
coQwXn+hiMnTPfOOho+x/yEQ6vmniISkasThE6XySIDgHKPpSjHWAtM0h+m0hRk23QX+kvMIdRl1
iQa14eK/ruLuFK1eMkPsLfWcMim4aHcVtYEsaKl7ccvxGdT4fwnujfXD2+5Qme18t6y/oXXXx+lp
4Cofka2tOsrlIYeD6SQ79YSGSFMTZP3OlThFM1EnOTnSNWdsCw3hnB0hdOmXFOQeR5k3PFxNJWAN
DEBuT7Dt4GyFkMtNduL+uJpR0qtbJGlVucD9vknA0pEiOWB29XD02KypIp+XxAuHlLxa9/YU9Qex
J5czo1t8s+D5lfSKep197in2d8M8wMejZG93tg6u/fBlLyjjIvMlyAYp1Gu2zH3xcXLzypmU+MTh
XHzO8vQcrd9bEG4RIe1Ojb6m9zU6/goXLBiZsfefO8o+Tx8boZa9MjJLqTmhOcTeUUJ+IgkQcE3C
BQ9qIPh039RWDLAoaHQouIN9Izd7NU5b0HXaTgzbAZL0xXYQH+wExMMOocMUlHs4vFWYPw9OoHIk
AF4h6esHBhuqD8dYZ0Y8Z6JB/VNV4DFPD6gV1U1TP6fgU5oBH4AnMjim6U4iAyE36O6ToYbhj0AJ
5XLxmEkW//QkqUBeoZGjtT863cxVoS4PYeIJFbS4hZ+3N0EPu59X1+K5HUfovPxaqaIW0Y00Ymjq
4e/5Mv+YTwqOjpcFcCdxaoriww14LOi8GBWaW3SbJaoBnT31TW1h3y2EGbD00PO1l2qi4H0Z0Mo4
FhlbS0cneIzDwbRrsZq+dwuJ0mtmeJQb5+VEnbjfUXCdMcUd6Bp4HFKgB7htFaKH5YXymu0Zl/21
/lA0eWsQ1btAtuLcdzjd8zSLt900xht0NnY2VU2MqAzfer2tqSdkop8XVWz2JvjIPM+7TJOBRdyC
wFpCHXYYOvmppcChkYFNAX4fBoFwNA2N+nnlP9nZ/M0gRTEEcYhRm+7KVW1vNRrLKPOakAqhxpdz
MjknyI53eTT/mc9VCWSVDrX3t0y5sDKogtSzoQZl2QRM5fwm5MtWogGqJzNdxsvbqk16VThFEioH
K7rR361umlptfnKJ74aMov2UWZqL7q2NXPacxn7vAO9uULIzLdrthR+W3sMjdRWKx7YcdfP1D5US
K7NVRKtZNM7VufiSaULTjPNWbmIiYXniGorTAriQv70QPV6xI3kIXAy5t4tkKyd5VszFnosNLUwB
mzkHELEJDnSOruQnJxxdKrj9XEEKI/u8Z3IR+QRxjP98G1eiYg+W7No1b+GjTUComw4cXHaelfYd
SShrWAOLZLoWYA4zpf8guSOIw0dxh4BLNfGkv4vtLX/DeoPFo5XmX1vKlV/Ysj5sh9ncLfLp6YP3
SBBNpA4ouq0ZYMoysVqoJvtCRHY7C1n2fok/5ATEeJKsRaSAgBZeYm/2zQDYE1YfvnTAnrQwuHXs
0NhbP0qryMU7vtbxxoppcknSdSQgSFekP7R6m0+mudo7Amw8c5VnyUYEbbIkdWcHy1ejY/AJzyvZ
bCnKJz+wzuFUq0owbM/cA1KoT2iqnP/4Qfb35jaY4YdEirEzrZ0nM/AdnIiBB75zlIgWt+nBfWbD
XnTbV00a/xI6Ja4rWoXsF8ZNZ4sBAHBwJlLLJWHaMNT1RUjKUYIe0s+yclQG+eZ6OUERsn+fAJtc
tIhHSfOasUGv21T3z8IWCfM1vo3/lr4254+0fUU0OrmuKu8KbW+N5vMBfM8+Xk6HZIQ2v5M88Qlb
toe2jqxw1fhk5QaN1qdRTh84bD01OfxgxZ3NeOjADT2nNfLx4fmASaHX44wq+ztlSgRMpZ61hHIn
CJVjeraMOq2u9NAQFW4BQQzXF9YhIIDOeClmODJ/2VoGIAGuob9jYEKw4bJqu+HqWQjsqcI8VpjB
v7DJ8iPjJ/Ymt5xOE89UHZArGBhSIZe/J3G3X33+oElIO3DrcAp5ta586AD8yNa/t4R77WTPCs+a
DSQcigW3Wqf5zu1gfdE+JOFJEN1Tql4cwPE3gaN1Zqi1yBkJXM5Ja+yyxSBb56FAsshbnCzH0d5K
PyZ27sGByXS3+deijbCfpqwo2sg0NVIE2NihjZM1wCI4053JHLGYsNpk+POM5DoK6MOBYI1QuLt8
No1r2vbya9ngHu12J1Ut9wlzxmr9szMVW4d1fF5CRhyXIHcsjhElFHE5AyNx/kX5dKGv1ym5PD3+
qizZXoEAiYjUWDhao3fpewOHJOMw0qVeXdcWraQsDZRYqIey28/N0AGPjMviTqlU8NHRD8kVeIRq
hOifdgYX4spWMd6A1sB/WlE4STjSmHrl4Vi1j9/LCAye0Cfgiiog9C5yCb97AOmwkGE5kY4atPqM
tZTzDtc2/SErFYH1JQMDkThWy/vXLjp8ZooEL7p3tLV5D7l3ShDAxV+nDCUdxKfHspaZk1KFdojH
LUOmEx7vlTKountJx98XknhtE7iGiNHACM0Z0LA8navxE7TbKdZ4YW5DUI85AFs6rXt/cMfX5OkF
3MeA7zXwbDc5EGygeK1nZg0FGROM7bGkg41sr861HeH58Eav60sqjRls1usxpIfgwxl08c6JbeyN
pCtlLPvG0/9Neqof2GH9bkmhD5glO/mxUCloyr3msWvJMsR9nPrX+idIgIQD/sOulULiY6Kg5hv8
LSKaBFXoEZvqq2qytfa1b42Xt668OVCFCVRmnhpH1D+M6hZrqroiLk0hpx7TeMEG7Pyw0RSNW9wx
ZcoSDQCWmQEWVW+2MT9T5bH1xtkMzSFTjVwaW+fKcwCOK2WGqYD7A5iQZOM9GkRkGWpZ0yonvHq+
6fp1onOzt8UMbhlUHGqp2o6wNBxmYXmkoVf2mrqVcvVAGwL08bM9cNfn2E9pw+GBCublxQ9DkBJM
HXYmT/Fgs8UybtuX+WwUDZ14Xhi4hbVn5RbG0TRSvEBRZ/2V6rRM4o38HqXhG7pKY3vrdVyMqCrb
RJX/c/sn/OgC5ZR7prblHA5xjF+vE6cn3SZat4uOnjSoLjEsyFa28dvKQFG3EfEh5GF37sm+PjyW
KZYKnb3wme15ZCxrtE38GNE6xzeq1qG5u0SmYKttOguaL0fnpy0cHFgYppGoqRq4nLd2JuaeF58Z
4WVZstzE5CO+4YUvGaecWOLc+ESw5sahLeFNkbHxtU40tG9EMbiIdMVPnov80WzTiZgZsXPggyT7
/xauWO9u8mmipQLA/dbAAyBmPrSkPgLF21kJdCtIgfaWimeosMxk62e3Np2Jx5A0AvQvW8nhK7qQ
J03dmSDm78ajPuGxHjFQNx2wTGsIO2BF+WiHnBGTDQI95ySkDZ1u+QXT9BvYSGWJCksBfVXHAJn8
Ef2hTxkwZIjgmXP9mJbDvnIovvrLBA2hOa2sJ5HDup1BQmGWJ4SftRn0WsyKOBN6NnBZjKAUcMLN
CcqRiOtuSqO9G8EKuQkBaqZKx231yViinC2Fon7HRdKKg1WAD0/klb2s/9gM+YgsjKZUETi4t+J3
hqovKCZrS+VspLb4sEtWlWgecnBem9AksdZvgARrhGnY7hyn2hCmcJxf+ug3J4ZNGK9a/E79G4jc
3EjWGHTfDw6Hs89u3BiPlY8+dzjZHSxMv6826Tzb0nEmeBhgrCLxYzz4d6BYuhd2TUod9dBWgKo8
mnKDP2/6hyDv1vnGZGVSz2RNrAqCPmUVoMzvvSemIbJuGmFrTGbds5XzD4Z5mnyuB5bukF490Kq0
80eXQXlXURVdyWNli2toN9fiGDHdZ0THTpC+2cpdyElWYOnRPs9b6cvslquFllQ19Dh2a4wa6Hqy
Z/gM7/C65GtF4qajWcbfGASAgblLksQobED3HA//SO4CFbjHMhGXndlWTaTZfwqRvr5Lh0HCAwHL
6LP+1EXW3A4wlicErk0NByAZbrovxnLQ9F6ssPsyfhbIekoA4BoJDTuwA8PxGvIiTwxMvQy4kx7Z
7me41lwwYvfCGV569/+XU8BnAnmL7AmP79b60NITcp5lf1AQXvuXp7fyQahlVfgQMqnbGOtpihue
ZD2y7LN+1Mf0epCdZdFmmNQ9aSyaRKUnVGmUc+Bj7BntWJzB5eeQULC2ovrMRJ/vmPubj6mrxMuK
UF/0RoHt1OVOOz2B6rOEF8vh8MLEXjtrpGXBxnppjp4M0xlF+UfZfkV3GsrX+dhoBbEZ2R8OoAbX
9L9WV3Eu6zOEZJkERjgG2jOdV6Dc570MXGxHfV9r56KXVdAWyiuM0A4WzzIQkcRyuojmRi74z+Bp
hHVXbFLQ3e+pRDj6HgLhiVzYjtj5W5FmMZTJKzGViz5/12VTjm8i0sdJKHKmR2Baq7X8tBFO/zuC
5HqPwEY2ypKmEVCMxssOOe4HWsC4PoGELBuYFYA5CdbkgWupS0/hCdjAFzY7WomWkRJ8IXEkwFBO
fczt3cNDzmW2kc7N0vHqmN5hiysCsFD/aM4MpD0RwPVzUY24tyRtcnq8z4iWSqLYjGuu33Sqnhle
kAZI4H/WgnX/6mTsCTsEq4DHTp+g7JmmzYZCe/SGAPN4sMxKME2GTaQKSqh8Us2SOceeCyxq0EtV
RVoTtIDWz7m0q5c2+R5HOfQjskvP5gzxFYR85/u00Z8lB+QlWa4LRIlOMgAc93QgOk22VKLUmbvk
aogE9OPzp/C9XxDC4MUIsVWAB81XTSRUPeebz8jm14/TD6jqgAHz2/sgwZT/LWppp8D+KNX1C+Gt
360cl41avZp5QpdsVLPUbTzA0WI2noqa4UZQW1IB7aLQuMKawnOIYTULi3BjE4iw1zdrBCpINROw
3OvRNpSYiMy2ZmBEVQkIC6uBnyRbcaRQwjANhO4yvpQrn9iFGVCl8rBgDTd9Cn4QysQEFks1gouM
HDdbxi5ZkF4EJ7KdNpScPQHSGMO3EX6djDMSWXb1yQy8uIac/OvmkRLuktvZnc5XRwpF0ILifQyj
mkM758TtizVNcL0E4LGwUbntbwUtpP1cnxyhe0swIHNEROBjk0xlbmnZlMZ+ejDRWpCOy4oZSNnp
eaPTaXFh60yCc9deaU5q5aGxmJZXPcESoaDzzc9bOQ1qaZA3mH7ctBe/Ql2IinGPwPX5LaWMpQ4I
IgmTaIFd1qs/eVczeTsmy746u/hZlkivhHthWilqAgfPQoZuEPie+NxuTBf+A4Lp/LGPcFZ1KmWa
0OvBJhS+EGlMVpIrSjoyMUiPgB6J5RqGLEH9gnr2HorpNGxOzq8NmMhBW26LAIVg5pzCACfS+J0C
gKSQ6rpmwGbF1Px/t7fKiVjh/+48kyRtQsnEfN2iVWAQIqmXAl/KBmlIHXkPr+TJzkbrnIEkD5hu
5N0yxb0slY2KKrYvK/DVivL3vzRfKtfgCgv7lFiPSi3liJB8A5KeJ4m6M0jKrMq5VW5q2/hJQ5gq
4rpYGH5dYwwCUtLDX6Jhbp2gXSprpPTqCM0FVk2mHUzNsgNQ8u4rc3NZSnu+pnFjCZHHww7/ZRU2
82prNmZ1mEvGbtS2CEgsB0UjCZ/g40w2piPLVDhNr5NB6K74xa42fyXi+wsrcn2AqpDC2gZ+tVbC
aTsaOqpQN3cdYJdljTUGa+SJmALO4eu2BHIzOXsj1lYbVCl+3740XiMCWCTCjDfzQQC5dyKmhHGL
tOJKcffhnw+qzc1SHXTbVMqWUGHy9JzfsWh7xMsj4bRaujoVbQbHakCexHmNaXRnbuRYbt3IiCD/
sIvw+JjaRhL1+BRjuCLU6IPY/o3+kya4S29Re04SHumjAKpPWLqZM6Mrocd6u4gmVrcUFdWgHh+m
FNeAkbXfkhioCabWZXX4duwTu+I7AUA4ql12VrjxJ78CrsL7KwuuYWBuTx+FBpvS0f34f8Et4CCT
9+msMx4LBMoKLfRqSyCl7T9NYSugO7ZhI2OVz/hnyIbChuNPQXV+9l4E6uw0FEOLsWe/2Ebb5/vU
FiWq8OUeaZW4e89JXM0r4y4I5vb4Ia+9WuHoiFx+eUAykz1Vcps7jOJ5j7uZ9phTkuCIiyjSlJU5
4nan8PpzEbtV5V1xTS5lwEjA5oesYhH+L50c4TJQ7iN59jclNuNTPzfADrSTLFiw/fs0Hpdm14yn
KEhBUA1dAweY1rnNT6b1oV3ls9EtqxOGNJCKesSqYWGl9llPWMpzrbTBLqPxZozObtB1+wdzCR4k
41D5GF8vFSX9A9VoFRGtiHwGriYCOdiOJHRK8e83Elwl6WnVWuboialLCSq7YCxDD0R4Nn8st1sO
bl7sso4w4APv2Jd8Jt9ZPRx9fxYBYRL/zgemeP2/kUJu+2ZhktJpxyH/i4t9S5XiKCej3dB2CV0H
C8muGhfKmoeIL1pWjGhoSMZzM1FL11t+rDi8Hyj37jAoCjLZHZE5X8eS2EGCj50jzsoYPr9Xje+B
bkCIJymRE/3TaeBXQfWgl42Dw+KlmJKY85cYgsnudS7bBM5aVbWPag6FWZDa1d5G819r/VadZZ6G
X9483XJSMJ74/euU4eaWrVDSTwEjZe7YNDRkVavHRWeIkILA0zyU8VZaLme+zscKieW9gTYF1Q3r
f0iymYUNUFKqSyRCKXkxIFakXd+7intQ2+YhnmzCpH1FFUSPwQkcIvghj79vPJiYD84V6LjYc1ys
eUHmOjbOmobep+ilAQWuR+2pBmgmk5RHb9S7wmB20edha/GyjPn3fLXASTCwmnMJvYcsYZAaB5WC
cyxc1aVWY+iecbdrR9THMigT1eD2UbdMY5Ia7m8SQoTtaIQRfvv9/dBuOMBnfiBZ0rJdwoKBF4Fj
JsaDbsO2Lr3sm/E8wJxQ1vhM6uzdxxiAZgOoj5RPBTeUK/lI2oD9zhY2rBXOOxKZ4oNoPrsPppoj
dzuX3iAn8647sJcJ15bjRD91qC+skfTKOoyGXMPNsMERZ2RUUjiPn42A2ieIpntyTwhqtAbAcdwu
3eZQi8xyUoYDQcZTl39MK01vQR591swVa7ZjO1nx4wX11S9URjB8nsjG8ecj/9QPKP2/yXnoTbUM
flV2M6vZSwAcbmkdZxyNUG8NiiDS2ZPZlFBgLdqeciWW0hzPx1bv8Uykuujzmt0Ks74+ZZVlxv41
+R5EkmRjHC8neIpZjxZijczlnMwo3a4zy9xLshCwByz7p5O0dch8VfTSnc+1S5AFPd9zZ1W6bSUk
Wi+F4PxLKYSePRh4i3URkFY6jEanWnGhzXIz8yGcpVeHxX251k3kGqoJ7xEIpRrcLZGzmxBTgis9
0R3k+stJscV4hM4a/Z0VOyLTSM4QCPYA/w/ZTT58LFRcgmDww6Fvobvpp0RPf3awfLAiCYH5XVv2
ExTQQWhCQJCQ4w4QQVCUwXRTxJ2Zm6tw/f2wXHCtL9Bcts0+29gIrZ6CHdO+0zEBjRFYDU2PJIPe
VxfkvRhn0Y28U7/YmWoX3FdHmOP3aDXoWPsJYtmcMsrwfi3Hz7JSzg23cQ0Yof5Ehob/2xYbreIl
UrAkkTwLzBTmOsJSj/y1ZerrKV38T2RlkbUV6qgaPIF11CJ4qX4QG69MGEhTCOmQJ9B3Uxv4M/eV
lt4HkfpZ/8lQBHijusdr5C8yJTVFnTWCvx1mRieaeSseZXLtSvbTDceU5+orW3++9jXrS+DWKPzR
jsxJykU/yHeR7x1oGxtcJtUpl+hI18VA5DHoMyNyOtZR3F7ekaod1lqNCDTaed7uA2Wtii+bVcLW
bsuS7v0mGIm7NQ39S4hwObxhNY+tKKhwlxYOA81MAWQSlEPC/cwsnrF1wdRVM/qJcpF9DjtZSPFo
qoA21wLk2KeeEF5EhY++8sr5Of+w0o90AxAhiJaRjyqCNymHvIhoziCIa7jRgZHOrK7BPEvDBHQU
Cj19CHXzmFHrWAMTN3F/RaA4Oyp4CfzdtUjxQ7y1SVcmjHAYaAbbzhxk5YOdvBgGXxeolxxoEoYN
jNpyBn+QhzXKJdBapMmlMzgZbwQREIndRK5EfLFKSHDaXOTQpjB/v6OXwUryqOGwoZteBzlvwHTS
kIueegiRQWJ26+Ha0Y5+sCSyJH/h1m348rNQ9KT562jHjLogIqsxwuAbiS7d4D0O6n2Jv6foNlTJ
Udpvo2MIkgwTc4csJDo6ZP20qpNh5KXXMPdD2ZjoS2WjiAsgQ5rQbeoIch/0hZmzgPJwu5jETRKM
Z4bJQjsYwDLevSYfADdpPxSf3WWOaDpVJksU/x0o7zHXFDoGU26DASXGdzkO8xvEw/0DIjcXIBc+
C/MZHOoImqIflUjRXUCwriLjuW/PsGJIlw19YVViw4FDZL6ACiZyXMjyNMDQ9/CxKw6CcR6yAJIZ
Uwmcj5BgfxMww7rgYdpqayK6ZOZXQP+X1zGCas+6glpI64Z5nkiFvUqktJwxsFuAUClBpfd6BCMb
EwQw01HMvODO7ArPTNmcbFWZhLCUn/ulc220QtrmkubDp4ScmjEytOR50WgovGLqHpxHa+DdRMzy
SdpqEzL0hBWns+y6Rx1qQI+M80IphGZnPdCt0q76qQyhzKQim4C+xw2HoYzmERFCCRa/8F44hXMf
TM6Tvb2F94JlRM84BY5ZWOuzH3/cl6GHaGpNzLlLi5APkBA1CIsunVh9wjRnIR263aoR2ZRcHnJn
26UMYxN77UxvwQxgVKJBm8Q4PhaGWq9EKYn/1eRCCN4p5QfFthXipdWUbYewQ07tz/LzZZeI0/eW
aG+aJM+PnaRxAUMKYw8MvDmMwZV2fE2RQxwcNKHxdGomILDp7dW3qW6ow+whTbWejrlZ1NX1ozJu
JaX77huNhfmdmT/2GHIw2URrqrQEViFPSdlcRqxNI5l7qifcPuv1HhekSev8WRyMoucFE9huGEsk
cmMWRWUuhQXbc0DNjChyGP63HjofWaycWwPQPe0viuA6pdyfQ41SRBv8akGZVvZO05s3Ul32A8L2
DXk92mbPAliapRe6IeM8SFBSjkF1qnHpfZ+chu0TJ78dZlsmmtivYh68Dy0S0C43IIrJFYM+mLBD
1aDGv1rYW1YohNE3jgrM/nW0AH0cl1F9wtTWNqdgyPCiCzyYdMHaEV0+S+MH2R/FlPrAc758F9nX
WIk4aAJUwK4vwsl6MSbJv7iqqyNT5r5lL8Uiyp8lr65jp7NrpqMjrvTJZOEpR9F6DN7Gr5cYK94o
Oy5e9BprCBKytwR/laU3d2Xv3khvIfZpvsNJIQYc9/Ll7UlXF/JCjDoY4lJCTLg5TbNsP3SSR46g
cEuy2j5fETGYqnUuXOlEkosBxeI3Jb1jH1Kjmwjid3CFITPUFLd/y0J4Ptm1RCE1Cka4/867tzBg
Ea7Pl497slv1UmLd5AFDiTfsxB4AccLM9GijkATKgo/wYCgn2IZ7CdtF4u3pffWfuByMrwWFYOb/
0jw+jKgJltBVQT7pzPvdWElhMstXPVhc5jSlG67HTpFyjeJq7NNTp6vsdEJ+hUlbjWGAGm8tXWWc
EbGn7LleU7lVY78DnQPhdAfJpgzDzfD1U2wZIrpjDRQ7pm+0GqcepPfHZm7CvWWVG2++QVdpak19
trb9bwtCkDzPHP+5wPMpkogishFN9EMH37DANYF1cMsU27henuNNcPnHlj+v4s2EV8K+/DupaAeD
ECA9sct22NzK4Hsae3/uKDh9fpffhFvuIe/ukfKv6K+dxM5wt0/HGWXnCyz11NCqKRy7ER4jq+1u
lJ6s+SizC5LdGI40tWBOUiPH3oCN3fRagWjmfsTvUlCiZ6/0UAbjtMgX3tJV5YhxcGbCtroIqXH9
miXIO2u4IRHYyENlHQNkLmUeChLRj5j2yJlkRXvRNmcgvTtBQvj+woBHhVLAIn81nVGLxFot0ewy
UAC8dueLu6+AqYgL03LRat5m7ygvz5R5MAQ+AfrdchovohE/nGmmecRgOAPyhraZ14bu4UbQBXE+
nMEtwA6XGNzb44NHoZz0xNRnfZqhTXmMIj4W0oaZ1qR8cdIyOX7C+SCupKrjixzgtXAnzc4+w/N0
c7nFb7bp1+pZHNRRGmw7rJgKwhfmsdnC401Gui8FnkHuezGeBi1cKaSq0ffurhvn3G3m5xv1r1Td
nYw7jSQDH684lQBegJBGl70oiKVkOMxqW/jQMz3j2lDzwC+GMUzTIoX85SJ4YTKTvR64wQnYLycd
cRWsHQneyPBLF6GMJOuvhQ3ckHKA0fOpqpx3yvq9kDNgS9fiP7X1jyV0ZQ3CYORk0bLPQhUayjIj
AsfIFhK/SctbvfjCmHhNB4cvuuiO3E64VZ8SBJX2eyE1pACx02qXGOi+nx4dQlFut1ph379xz63Z
Iu3jvusquDmEEmfKs9zUbjwbXm7rTUsP3fWG3tKykwTeoNmn1KYWkSp/Gy/s1d0Cfmvcce724Jmj
DfGiU79tw9iTVB2it+jaLXmn+gTRMkMnE0i9QmI9C20UxCMsuYjqg0zffh3tGXO7ZnGTYkPCO7fT
wYCwWIa6zU/DNKEq0krgDo8wqzZyGjcqMsq7VaMbl/TWxX6EPK/Cjd3srT4TlyBgPPpvTmHUaW5S
Yl3A1PeZU4GcgmnnCliWuE9KhfYWsLQc2qmHzfb1fB9tnNhmDcPR/N+BdUWcyZL5b7d71jyeb652
LBBjYKY7SHebhkD4Y/HgtbTdfpZkLsWKBiglismtZnTbLMxIgGvIZZ6i2H3c0zitgYIylFVW9Xvy
6xEZI204KzU17SuobBZ4ruD5zIpeHPXeVLWepMJmvRqNOqJmicz8da7ieqmTXj203aUrlW9jXDXT
UV1+8/KgMdbnKTIP7+8WNZ1iRK8pyyERAx+6R1gnW3MShciKybXzfLR9BQ4+UnO2v099hMej/Qwp
u64aftjWLS8ApjLowwweEf7OWVVyeWdukyEjE0uxI8Dx6KsG8G9l8USskVaA4I0u5Fwl2R/NVIYC
8dKmf0QvKlkI0rWUd99HPNrhpZcodvj0FdNCpZp00gRrWa4ca45ScI+cHdNUvUC5UO1KIHxg8ulh
ifPPrfJhOqLdjrqBsHyv8YaXV0kesl35OwNVP+V3g6Tm1hs/yXhTMqKv6ih7woj5Wb7UauAoFKVA
BdhenUwiDp6hIwWmEmQJW4x/jcCHBcL+WVVP4BYJvc3FkW6agbczi0euPNCsHeMNT3YxVc40wmga
bu/BaVpToIASKxrB7k36OT8NCUPrN4JHqoDdGF1CEep87Bx0f3nUfj5w8RYKeZ7SovnZidd76Chf
d6+n7nAj0Of6wrBaJ7QS24vOHQbuWypdN5NYMQKz4tQvyXQ8obPE97m6whpc6eiRtEaEutQqdunC
eCi0OGo4eIaY27b8lflYw1sGarHUO+OOlxVCX+IyFSF1feudCcmbARt/Vo6/0lJ12HIqwsK2Rr6H
tw3emcLmbaK55N59TJIxCJ/TgJs/RxL4iZp90mOcrXuXt/cNMzY5w47JChtQ+wU/JewE+/LQVHsd
PIiW7ktcZE35YQhbjGj9vBt106MwYR+cRKxn0Q1ec6g4m/hCmf0Y2yMjr+QHA8aAys4QCjsRV1Ks
qVzoJJNeecV2pNsd6g//SKM5YF5CdIgbywF7OlBzox4iMlcKC3DmnUZCBsbtfWke4gXxpadb1Zq8
On/pFKG4K607DPt+Ds88Z4hsFfkCShAroIWYsjOqJd9w2j2C/f0qOh2WQQIGsZiBY0pgOAzSo2Ma
oUqPPyQYVZsHe4zPH1oJTl9ULhg5Fk1hf3Tn/w3mNPteRz60FIssToW9FijfnsB033lSrp+bgZRz
JTQ0Tuv8EwtpZr2gom20FniviX2UwsOtyPYxmVnOrDwRJUkST72/N2gymAbxcAAyuRYyxwgWgWY/
hVcf/piuKi1zscavKpgfnE6gpXMtIGQS5WGD8IbPEPBqNR/oeNBPHEIJXhwMFon2gBqoLpX6LPcc
RXF/PWxTHZLTeHy/Hy4DZBGlROw6JARAL8WfmBbv5t1AZJpuym3PkOT2Wzfhx9Li+bEdb1FaXw0l
BNidu4LAxcDZjeXHIkk9Xo+awP7tWzrmgxf4e2q8wQwrOIAeif+NMMOfetkRz/yjioFcr2THAkZ1
p4ySizuu9b+CsfLsmoNDqkSD6xV2mw2vW/YlLpb06THYA3UPwj6304J3vU8XffR3DdExB3Y17ZQ1
TkBG/baCBacCViAKQhV4e8PmWVW9yzbaWVFV0Go4wopxTUCtkp3D8OiDYuEDE7iM4ScjSXXhGpr1
mj8K9utGtu9dJ6Z8+330zOctNL1R/FAVB1g85njuOKud/qrh4jWXM3MjWI0jXSWNkUll62SK+ZMG
Dgk8eZIR8LIIjtClw91rmDwWz4ydonL3bK45jUuTTB6gxhwHOo4mt3hkw+Y98QNA3upc+i6jphXE
m2eVOLDkxG4GmWTaB35kHboVamICjAl8XcedIagwHq8KU/vy/2mblQrhlM5Wm7wJ9gVrmpb6up1C
wNJgtnC5EaOK9Wmh2EQv5tQlzYm5iz9+rMuwwcR0sq5gWNp0lAjrVIKzSnswC3riveadTl2KIW4Y
XnhY1p/3oxsMNDULqhbY+fH7ql8am2WQZ91I/ffXPkOxnzpWMJWwzcGn7Q2WdrlB5Q5ZML1+J5h+
S7WRGRXZ7uQuYb9oiEuOT+JD4HYPRMV2ng9bSy0bywUNiRisJP5vI/GTIDv39FjrLcKTYpbRET2v
pR6g8XtmVhHj4AP6LepKGBC5EB+shTQ4EwA4oOxK1O38Wp4Zj9QXSOAnM2SdaV/URhB5NbM8o7Z2
q+2OFWoRomol/IiacuNCjxHwBy5zRLRlKHyB5/kK7SnFb5KilJ9cbwmZulgKPJJY8P0Ak2AdmgVv
nLbzrW0n6LRs/4ICn+QytiHr7YvrPBAklWOBsUJNnlnz6Q3pu8Gt1HozxwX21yu/Sgo6IBjspGCe
ZI2LL/Swrg288FNKpoY1R6VJFBMSQTvu4e2txvTzSuYLZxUYaLUILxxr+By8KF+3YsJ0qE63zTrJ
x+Dh3Y/RrkmNBDZyjaQZRai6l3QZzFhbeQVjzsYT7Nj+lA8P/EWaGrnzqKSg3waw6cwfeyzH1ogA
uKnCO9TFt9ab+GB1KdnyT16c4TaI/hfDZ66dpEZDlmNeop3Pf7+1sJMUKsbgKKfv+o2iAFO7FOT7
D5C4s2Ql6AmpJU77qpkVQSciC+Uw3V3v4CjAE/YYr3pboOMic643VC38w2OE3fXytBxHbvggTGAg
3I8usib3ATPUTJ744aM5A4b/g24n8FkEk3D4AQDS/whvY9dMMQq8WqGjYr8hwoSCNF/KeiSmi+54
b0CEfy6iPJkh0ZeQJFWukhQv/QbqQxRjoebwx9O584v5VpM/9tonUekt5zx8OjcK8mOzknY3krAh
tHwQ7AAqR7legin3ybGlFNTKVALicUIsytz1sUDaK8Olu95e/wPVvaoO5SM1Yf3oimpwYbpntdqV
vJQC2vsBLlzm4biGvjXgvEaoueTDIrzHj/y6TDYa7Vlf4hSGkGpNFcATQ9kc70YnO4yp0zjmtN5Y
EkPEJ6tnoAJ8JkiY5IYjwM5zNRPqOITN77B8xa+D7BP2vJYPYt+XX5zud2kOVvR1krCrkiS7kq/6
whYGMF2ar1FfP5viZHmASrXqpEbpExInciUgGkqZ+/ouDgY5qQjYmrAiwqc1lROb5gzTVpZZXoH4
bJRu8symDHE76FNCVhOWGid2LUkpJASfnm1MuiyO9WaGA8NO1Hew9hkKQ8lirWnNySLIpXMn6X+s
qMb44+t8YZoep331/hN1E1kKYui6TqjULR4J6oEg+vZbqCrewAgfuqm4Mu36AHLpnSAhrknTeJuM
qZWsXqzVi7VUa2c8Mfkxud2bGI91l+CSU+txVrLmTIfTx8duzpGgV0mlTV4zV4Z5ltOHBEilDbvP
a/oyQK1gSgKBwjRzVYK5KllQSIXRgqVKro5A7zvSN64jVOhp5mtFmc4UrWpq5xPhxm18m2/SlR7N
dVtdoKObE4K6iRU/TWNM6F4jhU2JVeizxMaSm9pq9Hcvv4VHhWN2i95wWp5dxcBdE2Of9v4TWzti
uUpiFYeU1w3RMBWO7l3Sv75oLoMw7J4zUVZxeHqWjgWxH/dRYpzvqM9dUOkNJ31kq88SpfCZD74F
FXQIhc44zrW+mf72KTeQc+8xsn8thbtsFS6sAtG3IefBeWF0086FsFk2O4H0D6UxTG6ZcuRH/DYc
9qZMfYCrbrYifnI/qMVc9Z+DCfLbnuIWLo93rSbwRsyzI46kBE1rERC0N6ooabPQOkhgZivJdbrf
VxHeDR8792pLkacq9cCa5i+MOs//Hkm9YwMz9HxNBZvSV3fwP0AA0OmIOzVaMOwtT7pfUP6c4srZ
hgd6PZNyXeiMwpGgkWnLFTq1udqptLb/TM1W1Aj004sHYBbrQfWYLbkufT3KqGxx9CkVXt2Y8nbO
0Sk0fbkfIXm7wogC7wLjBSdUUySJTmaixMjJCtlU/doyyKw34JR54GBLRpmBTwpOz/hIKYJxwC5p
g8iQak9+MTLO6nBUY3kbflpvJrR3j/F3njDyNFgy62eJstgqwq4yNXRY8sLMFAPMq+AxNCMbUkH3
LK5EUCda5whbrp6gE3AyA7FBglP4bKGSC6V4n/5ujKoVb+eGFSTCMDc/MYD6aiXhyjSCnTl1jGbU
CRyFeu0CtnM/AXNl5aWTGBVJn0tIg7r2XMybrNEi8AsPoFHrTYUFqzaveMP7qZDM3SyTduSdD+Uc
6ZN37aGd27Q+JwlY/6pxW1LrWL0B6wIUqZLsp3eh8/s0HD2oAQNQRSblLnjmyMaTLI27aopA/HuG
kohFcf/yyl8IdCHUXweVgRgeguscsqXuuQMKY0IJSoFruD5s06oEnowMZnyksx4velcINnDPEEiK
HbBRuqPW3EMzPLbjUL5eYrZEcqkU3MEEbu9+XHenJYq47JjUfOZYdPvNZVjGLNtJpGd9PYW4R2nB
wliCLDrIN1f8rWWQg9l7BpmeNEQwDXqo5V/8nMj0Gcqh4+PJd769jayQzUmM1UK692LPs3VjLn9R
SCqxjub0l9nNin8m2UOLZqfoZLnvifuXNkyZ0HE+W7g9u1qsDMj1fGirONLmx1iUfqqj+y848zau
Yx8/6begiQXwXlvGQzcOQwUjPrHpy1g6Hmm6+XcuPTzeT5f8WK17FOAHVeOpWg/YQh7QOqTo8Kwi
G5nFtkwKAlgR3vrGwsRNmb09GAX+9go4cLYY3dtCkY0ZRhzGVDgl0jWwbzK29Or7BcgI3nK6bEgt
RlciVAt53LWAmQpsxh+sHBykTpFuz+H2jzWdtPlNtur/WtPT+8Jm6R2dVzxcNUxoDoBCsFa1HM9i
MUlfAb0mXrMR6rfbdK6LgGWRGmk0rxYQ2pztAy705w/tVkciqPX6uNu0RWbCeiqiXhEMuvNLFZ7g
G+UcjNxsgmKZM3CTS+d4XXttC4pfisqO9KKOqRQJM2P7/mnJ6At/ybVnc3Ha7zivG/GNMuMDbm5x
yQVkVT/2navCWmBn/VU6xj7qpa2VtEz3LEaL7YsjkxiSvI3o6/HRDuhWI8qgiCnGrB/QVPm+rXma
qJxG8MCKeJc3SPrNcZ1wpKZIVMZezw2kLAhsVswjheeGBXadptKbW6ZR0POb8MWpBstfwqRnVDro
ZBLgmKd5bTSQR/FI/XUdYV3QAPfyG+Mu8+iqRpuq/COH4hDgZs9NdASMukYiz6gJPchRVCapv637
81ZjfyRvTvW8/ZM8uJ7oY0Hcx52/CXyX9a4WvrnRzLtuuKbBWq04Qz++SwxZBIKdemqtyqy9HIYv
0bMS2zPvaV+EmITpxT45bpfjbZhitJLytbYtsk3Tl9bLnR0rTWy8VWsgZ+CHeV8T0+kPazszgrYg
r83ALLjYbvkwgTfcL2u5pWnYsU6lJ9qLJfeyFwrRRzyrWHWC0LG3YvyL5grrh9QPYv4C+kYAP9PP
JXkn3i9HBq5vMxHtDW6D8juMcNeApgq8slj6f65pHomX/1A/o7jXbciiLKiATa+798MEVf3DfAFU
wY+blTj6vGUhUCVYJ2w7oi0Hrqr4Bb8zXe+2lvbu3BDqVSS2jAhRjqYrU/sH7zjx0SrAXGhXV5Qz
7/F4Oj6Ci/4bA8/gQ3XqK51K12IQ4bDOxQonvDMYnivsgVRlJm6e7Uq5Wyr8B5ybduWNsNY7RYvB
Nzaz2MUsjKdfanSNQ98vVpex2kdmX5OJyawz6bnhJw5Bsynn8/BqEtWxn4oSodXtPVKLz64sBToE
s/IlgSpYuSMpe604YlIFgdWgtIc5HqF5Q8/Nq3ed/WsC2Ba4puTAy/rBNun51m6lTL5psccn8Ct+
N17ykr5Ggrqn3ReQgivM05Wy2psm69YGFhElHdDotVI9YuyK0l1xWrbTzXBe77VLB/5UX0XpNb7R
NFW+Rho5uvyGKnrsLA7HxO/Y/2YiwhIxdt/yKGMYLYJb7Ob7kEc210BKKJUU8Ed6y8G+SPDlm4RF
Z7ZN01KxdEOgucoXn846h91yZG63+RyTMzLvte9uQr8AnQq0xOwxVeytEviGclMQVwV/nuWdxlst
4M8YnDjKDxvPF9PoCP0RZXbjfcJ5foScEmq0Hh7DxuNDGMBDtWjNjsj4bojIB0PvFNrOCJiXKgd4
UpsUZu4cvDBMH/CjCL6wShocs8YQoIr7X1VDZIAbIqbbbXL5VifyZCvAKqVcGfK2arFqVNAYY2ad
OGFXmCR3bqbUXaQvYoWs6Xcsam+qxdiMIxOBuIOJcOKIAtUubEho6erGMLi9D0wlahtFG0YHYglW
+TEt+Buu/s+wdziRL+hRsHhVWZR4xn/NeI+AJsaSwycRmjGwlpFMrM39Q481Ob+tN0D4DtyQmWCZ
xrjMLURCKmV+ENpbBOz/Qt0w+c01UalzhrndyUyuPE+vM4B+bHEFZh0njq0GnfxVtB6Z19um/LGO
JE93yCvDvj58+0Hh14k1R5JUlWhR0HfqlkLX2OadWP/5hEOUfri53Aq1CHNUSbA6itkq7D7E7WsY
VpoSM1cRFT9tdtgLcOu7Xc0zHJZYreesYO2Vhnr2mo8Fm/swtpKwszsiUx4PVzL5w37ytv3cY561
Rmd+4S0fbn4i1y4hHLl38n30yCrODP074zBEa8f9/uPEklLuKnxJWm6bfhwpyLMtBB03BHLrvzuE
8Ibshq4WreO2aJn0BVYuaO87Ue0vDl5AxKBsY7vPsvOTzpC7jrxIHus44IQB9RMUoc4pYPK7N46R
xFVCEECl0u200vofYochJemwLfZOiinssBTH68ZAwmEQuCKHOpkMo6DsVAZOxuvcvur3SIFE6xUF
FGHCv9/FnYDMhPLeqewVzOp3lJeFVwuS4e49zoG0D5qeNe379RkjY8Ka1HywNBkqbfO5RUK5PSq2
Lx5kJcfgT1alxPknnbwfLh4VIT2zRe2/iMAXmoE4UO12PDsZQCYUAkWhDcqCOgGjy/25DigiDCb7
1cLFqUwiUAbIwg7HEolpeUUAmhi7zhAHRZ5dKn9rQgtya27AlKkmbxSwRsdr3xZ+qZRQooDnsBVA
WXli7OlkGT+B+wesG0Jfc4CgyKKUEYRZuA11LnwZLTLbCNd+cXTi3RR2xlajQqrH3CXD8VDfYLPg
VP6iXNH0AcmDyZG8mx/oxyccf0vdo22fVley9feCqf9yi8etmugHV0uo8YspSpyV8qMdb3Y9UF7H
YW0e15hCLNpOQb3uQtxNIIQ87heZ59o3zbzyn/THxL/1lW5OAEx2BlI6UrqsXhQ2fjiIly+Evq4n
YoXiYJhUpoIFHOTTHCRnvXmKz+0JIoTka6IznMJjGD1mgTUmCLJhy52gpFolOcg8ormFg0Zk9mKf
so44L4QnM2qfQ7tMS2W0G11uKRF2h10ZNXzZrbcTbCZi3IqoUszfKjdFZzUiW5P85J7GbkEPIPO6
BlLd/1a0zCpYhft495bqjhw1B/asLWNDkR40sfNJLFjEAF9K8n3NFTjuhZcFfPSu7Yabqi/+nWPG
hHbFHVcz285EnO+/1AQnUpA9f1AudRUOFkEPD1jCmwJQRhq7/3ZTaEpuliRwr2zyI+YvEhLiphJ1
D3NIM6Ww3q8BR3Anlv7hN6BSZ6kxqczurDrPpMd66Oxd+YyGZNzlNom2zlNv55oAO+iyO3skOsMH
ETapEZAUemsjU4NkS4R+E3hDdm+P/CVwcKjptP2B7UA/2H+sxc8nNS5hbcuoqOUwsLInefOXZGOV
HPWRIkEtKgavcqe8CMneJugxHFTerZjFaQcyN7wMYdPFBk2z334TgL+i5bzcaYPV2+EMbbJUafcj
qOaKRKekN2WSFG31+Te+OffV35Zms/xKIscbuS6S612mfpdVJUbHuLFLpYN8I5Wxjk5WRlO96i0N
Wdfq1jbrf5NjEqpTdCSQkIccfZN9beXWqZTJxnkBiUxXFSsAYjRtlE1h+MKSmbTZ750yy9p7xG5Z
woynlTWDGGy6ryZYUpAYzKdV5DRWio1+sYZsQV1atpKq8uVXYryhvaclAFH+eprCBgst/2p+NrHi
iAa0N18kpKWdbze0EZkGsRsDBAK3jz4pHmjAHjjEVuRRSewfPqcrprmWX3bTz4rbPHBM8fdfUPln
AEEWIE1gVP0Hv1C590+v+CYhMM6ATa1m9h2hJoz1muMumJ/vaBclJgn595kpHmnsygsynjq5W9X2
2Dy95y2vEChe03/BzXX/PIFVHPMREk3L+Lvpr8ioWjSG7JQtf8y5hcJFED743dxCcFQBWcZ2J31n
qGqspvdlFmydPwMryuKMtQgtliKRxiwdE8Nk8mcHleYDcz3CMFFgk2WiaQpjQJ7dIyIIdZZbxJIZ
xkFXmKqWBIjRGH/HTfhg71jBGHwbdtscelTu/YO+ccmy1SqWRipkUhD1Fk7ZEbt2TQ9+mtYA7o3k
PgBVRHg4KbInNA0MXRSr8tT5cr6MZ6pA+NIDEfGfL3V6uVq5HWyqMX6NaDFqbrmsQg9X1oxFNVIe
GYmiLE4lauRgmj+6+dIEJFvATSokaLcFd1pqVDvpVK+h8Mdgrkup8rQsmtrYYbMq95ye3gTyx/+K
2AsRq+uSHN+NoyPXl4EmGqEE+8gVG4DPbjlYq2SPLpjNF0Nb72krN1DWHKdQnLf+zhSwjhwF9NKW
to0NkYM012432vGbeqyb3wPvtcQtlFxsGi3p4MFyiTKsXJByAVeAZ/mGuEiYFJCHLmm37WFyXE6W
vuxOGhrrdrQv/bkbJLR0HD4nb7eRXWQACxaOsuiqV9mMElIjK2y8fDGvYmGWbKBWTcb5FK3FdWci
pzybXAZQmZKGq0l2oNW4PBpGCvHgAfAy6LAW0JIzC3YjuXmRX5YrXWELVP+71vhCa8A4IPsgqQ4L
zhyTVBzv/R74EF/8X3wqa1fX9ydwKb44ABKcuhb9thh+jgFE2YeitiGOWh3VxA00ALMasSsPtahB
2H6wzpvWy5JqbSDDXl2wWffV9Ioe4AHV/T+4BZp2tnD3Qt8HL5IpX0EtWV1oBfbbkrlVNF61EeFN
oexXYeDYZ4LZ0F4ViGD49smpOT2gdRm7jboNVRdCHsP0qQLb1BwvMAwCrHdshRxyCdBjs2pN8f6K
u3gVFDPvp13MDvecqMSTY8Xk8E+C5w+4s3laMWFc+OnRKMK6G+hq0AcfWoo9DWHPrf5apGN5uvQ5
aKEPWqL4eBK5YVly8jZ5eof8LUsIR7JoKbV5jkvand/JkmAKKq0QUGKbc8F3037dqh2NJ+RzXh6K
i1l3ht3NPVZdCll06nNdFlnuM9C6uDKIGHlu4SmPDntWS5958GLezM7tvNE/jhCHItqSrYRHTM8h
y79MjUTmJXk3l+W3Y9bVp0AAylxTf/5bpca2waxeCW4Rd7iWWE2EmPLfhlUmAm5HCyArQlaeMWgB
U8YdxvGzHBJbYsxSzsGpBBhzvmgKehWmOx/DjpoAxQejFpizWM3ip8A0V3xyd70HzEeYICR31uSg
EpwAhlQtUOsmTYILSn6WLAOqnhEgNbZdDDRHF5Rk4ECfzyx1GJq03TFJKmQJQRJpdgS9UNCqPOts
7/ch/8sehz+389LqkwtUMnCX4DqCcSCqeyCD7O4QGBHGvtsT2UMma/wSkh9ZApqM1UQ83b0qfH2e
Fe75XKb0xLPQulZK1bbm1xpgv2EW6R7UOV014tgPeJiAB+5gkpj/cizFJ1jvmlBTdm3kM+pxXj3U
pFuDOWpCUbCA5ZkqfdXmjnIB5KrM0JQz7luuAiHfIlNnBC+Zp2S5kO6oPuNeCkBra/Pvd/njdGSZ
Md64Rtg6hniXAZE+uHHxYb3o761BH6WMY0o4QSAVfxcJxOFloaO7i8OvYMZIhvFDZFbKEe1cQs8y
O9EBVSrMdCuSXhkVrb5ErT55dTLdnfUhGAWeN2ck8cbx2iIHZqU+f0La59iOAgGcVKJmHoCKp3WO
HL8RsXRj+FiKTt6sb030CBdUKkmbchFDKoY4OQKZ0efGt2Q6QXQWr6Bi5jMR9OATFi9vabeY4kg1
v/nERoc8iW03DK2LyoE7DLKbOAmNLiyldQY/2A0S7vSaZ7+Qru8UV+ObX8Lv/sS77EJ5QSJ2icIl
1tF2OZvc+nXvPBKFLA0RBEJfpTLkoQ6e5rvxVZxNO9Xku+UOF0dst+TFnYKc9m7SQZ0oigXK39mu
GngkfagXqzI8kgoo8QMNz0AbIE5FePGbEdMcZpdJsG2+tfpVOYc2NX00izsrXRUwvGoLJl4210lP
ZlsRcNAbfoGmVGp1R/TkUQF8CWdMUWwWj8pMIix7+I1dK6mF6QHYAT7KHaaSKQxLHw6O3ADyRHL1
butI2/N+l3TSDt01U0yvcDlOv3nmdqi4d7DukrB/TJJzJ68ViSs/yBl1mgosRD4IXPosgeQMDMJo
gjsw0CGq0yC7WBnhQFLaRpaMfmAwAsj85vGPiIpadS21NqEP/Th4aUTWrbVQYNWv5+WeRn1BrtKi
2NPcskF9gzLjUkoj7N4+5vlT08fjEj2MTW0/TMdQN+7401F6bdwJHdPHG5//Ut5fgzxII51qk6Pi
YSeek6/KXVzKJUdO1/qDEUKP+RXAxdPjcgiwFCrdPyIIjRCY+D98woj0yw8yMylPUdPRYIsBeOSg
D1lVYcLK+Bp8wmmQ1fSfMaMHRiP45IideNxbqYLLrUorzCJcrebGXSmlVkJvMJaoZ0dM/OAyRKwd
jKdGlrXmVzyzr+TxZzjEyjQl4MX+6rGxdZ1z+xV/yhOt/xSiY9tEa+YwFmUjA8Ebj9IS/43Na45c
FimkWBiUI5C91UP/3ZI03aDyvM4/Df3Zq5/MyxPOQzBmbdt4XsCueQV3J3D9sggdDZ4BVQGeuYgf
BvDye0Va1qZfVq40MMW3xDZC6RtcEeh4eFYw/BVVw+UKtaVlI/2bzul3roxuEovg5iNOS/md4y0N
ILcYbF5VrnsAYiw7jorAoABbIPFg3Nka5Iac4RkDMC3Bt7kLSh7hl061s9VFsO5XiqBubB1gOhdd
A+sB8GYFubtVoYm95SbuAm9TykyrdQ6aJAanaEuhUJN18eoJ7wH33G2F6vktIVBJU4ES2Ui/Qkcq
ZnAyeentzTz+CyyFtK6jUT5h8GOkRHxsDQ0CL5yPedH4Ixhd3dY/W3AdCxlryahVyWJ1zSt7G7WI
ATBlbBVC5RPlG3ST0FR1pv8K7GEecCOX/Lw/KPJHbginOcjOmKTZpAp9JUqw5v+4zmdjhIQjJTJU
zqBqxIIKrXDAzSGUDtnbIf8X88KqXVflQPdXdSMkK6z5rzkz9fyxuGiz/9Sta9hCTvAHaz+tZErF
6XYzV/bRJP98rRjlubmQbVEsCuelCI+4eD4bSJF8Zh96fGMLUR5YnnnbsxTZ05liWbzku+do3pkE
magBZjGAA3jaJMDt0klC6FKHNvl0UynMQ7/48bTMgWjNWCV96HB+qRa+E8h1x91te+w6gj0rwEvU
R3x3hoCMxY3r+qnOnePnqLCrefR2qMvVQ3gRi3QdEzx7fh6zIJz5xBOTzrzjFAD1LuYuExltZAA0
dpITrzi9C4omIeHaqSIL7FEOny6hMdMdPDGzxAA+F0oVFByvSCp/+qwK+U0R+zm4gh5q40fofD+a
DiNUzMDXlVunhtFUEjA9R1PW/xDor4DX20v5lW/UijoAxO6Tqz4GRVd6Dh43id6kiYEnWbIjDyZX
fF2bgzgnz4/l8CeJx0t1kWB02X+WLfoCmNQU6oaOBV7Q6L3+z4/0TNibuViVHdQmDO7K8ufX2G6R
7bdMJSbwDy/LtI7ghPXuWCDJuvoPpfslfnRTXpE1Y5sgU0XaITJKf31R9JVXHQthWzYutmqdNVBV
OdZXPO7Bl3pArcfDIK2jXkwnvT1dhl3U3xMGjJIXlo6nKMSjpzkxWdGoJNA67zXt6GvaSH2+lc1g
6Wbk+tsbtDVjXp70iF3NewaTwvJ4qxj2paPsZsp2cd15J5t5WAi5d7hPdZuPhswyZ71UGgFfS9Ec
TpbGlIAUlIqg4cJJBPfUnKtsOu1jyPnAfNFo+/LY0eR0M8rqGRwAhipuJ/pLn6sOLg1QGCJqNbnI
DdejGkvft8Mj63hSEprSAVkhR6ZAlBDk3how5dJUiUnUwAZzDFHz7BYu2+3/nEfwvD855Xj3MopC
BdQl+4QAYHvJUgDqK9wzBEjRFISY5NJwayTrFyfjzSP5kHMK9E+zJywl741NBfbIqBsetq9vpV1e
lXHaoBzRdcjo3RUUXsqkHxaiDPGgbUvcBInuaDz0y7j+ai7k+2/JbAs0XcFPQ5XHW9R32TYcujQm
4ykDvImIAy+b7ciwQmZHoFAnGpePjqfzEREmkyZXQ9H4gD5Z8FyXY5ccy3K24UGXH4U1TVqdmsOG
0a7435H9dg1jGc9zFZZ5mMBZhPEX/Ta+G52Fs0NaRJ5YxSqe4YOj2t0lJZTGmKaspl8Sl2lVLhH2
rFf4oyHXcSe+cifZpiMUm8lFwY2rMADN4Z7LQZ+xHSSMzv2hadJTdVg7AIw6o+C2QLNESSQrf2fv
N9wbM5oyxQT5aRUqVpHP6WhNofZ5omCRvfPqC4k3/zVB30IJEsHq7EL/wNRt1NMSsJHwfGiDaNBI
pGgdxiikZEfoXXE27zcSzs+VBY2wJcs1kxE64q47xATnsE/Tq3K71JJvINb66BKRlBz5iT08l83I
VkrWjX/kZan+gcaUm65xppt6DLept4mea92afkRrJsWbR3eQkjbLVBWtGgBslW00R/hw9bM5DM0w
sZuGCPlur0JuAMOxYU+OWI2hCeT0y/WV+wy3NSKYNB1ZXg/Oek9sYBSbcVv46aZc1OsazrOPfLqN
fwOLf1bXKyY72M2U7r1RmTSBQ491UelOOmadnAgeUdY2HHkvTRDcBDlC/AAwQKjVrlbhm77sjZK2
fcvydBbrH1prB/AnphntMVXY+Hx6XrspV294+q8SZsh3f+3SzRaBboiBOS8zj9nM1KoKoI1Ft7eu
C4Fx7T3eNojWzURKd1Uq0Q/NHs+oKoLtPT2Oe14Q5P9NxOGVuSrm9LYaXDefXPeaSrxxOXVFPeXA
iWIS79DVj+LqGoVggyVxsU4ZVr3bdEKbxfWyBh7DC3KbxD0JwnDGFPglUObdFbp89A/XhvAAYHJU
pwU0Becbn1WeeeCRiGbxTgzi3ikAbFakp3ezIUD7kHEJp4JHYZnjRM8cbi1mL8ot/Kq9ovrWkC9p
7LjPm5cNvjiyaVaxyoHl76NBcgcIayt7t7iulZSyTYy60IFCY6cViYI6I7H6bUg/8tKlsRTICG6O
FcOIw3M7kyhYH9p6OcI52+hDXFe5nDsgy4237SsTtZnUFbY27pEUc0c46kMKSRtvbUEf71kuuBTY
fG+6+M67+wJcTCqjTQTg3Eo5IP9Fmca3hlrZJlkDpH1Vfz+OMr4cdCiniQaB3j3MMi+DTI8oDayw
oRbXMlBbbKu5/eXlEyrXrpgvHCw+etJ7SrlMNe+1bW9aDBjIyodjZJGbJhVsAELz3i2Od2P36IMX
7/91KGLPHuADfvwblfxryO9qdJKNZWa/kajgMWBQAZ4jREw6tEO9xDuGqWjJsfnhpeU/nUQdacy2
Kt5A9g+vXKLGDg6HRSEe7OLe9/m0fbTI0ATC8pvyKNMRMlByzf1PjyzO8bxwe2Cg/X/dp04fZjTB
MEHmLphEcicxf8/8J5DNxGXwnismjt0HKNsao9W1kMY/xloX2bi3UFdjdVRBfDHpR9XwTo8K2Mg+
jnZG9eLCFzlanh1+GospBdzcuH1CTd8Qu/cFmxJbdzIy+4BLzyy2nq1FtYhxAf7IywintJwNjoHQ
pDqbSd5rt12xFWTzkACpURUhpIvojobBcyZN+GJ+k/Puyck9VsNZBAqE3j3QxENBVuiHJrRmQ3rX
KfjMIKhe8KEnwL03goUMBtzJFJIJCaWlHpjMxY3U2CHB4/yflpwlxznSvVFWiiDWhZJzHDFCqaR0
qQ274+KVJEsRMbXF+r5VXRtGlysOSEWlkjzDe0HgHnb+yuF7ppanE4dwkf+d0c6rM+qNoKc+qCZR
9AktB7UmZQxxXwyyq9ndx6w+gGOWa35s1ri3HoIsMdLygVRYcLnu3R1v+wzDoelnCJN+JsRKx02o
X2Z9X1DF3LBNfTAH8qEPvHytAbglJw0+xFIYwlAZzcEA16ovwjgJUKWtQqq9yZpd2hmJdHCMHbAi
m+LrpxLxqCNt05c6P3yE+OZypK26L6Ttd287UmwkVlWN1wX1/60M+CDONv5BIhwsMQiCwdtykbPz
nLs06bY14IkpZAwWdGfTmlNSbtlIvp2wxSfNIVMuqR5Oes+jlmI7gm5uxXALQIiwubXVuk1OAzpB
zNm9tiaB3UIy70Do4ze5dLh0jtD4C9PCDoMHFC6pYQ6hw+wTuUjynRurv4Yj0edYAthFgJTcF/gn
2MwLhsNbIuOnBmXau6xI6IPNEtPxXh/varaVAucno8aqFlDBn2U3bLKWObc3eX7X+mZ5IZvVcetS
0nWS5KBqEvng7kF8IlJuN45CoVWU2ACpPCK3s50fILDm2r4m91tzkL83+hJozmL0hAWyjpvujUn8
7XgjxuQgoaqerZ9PPjJcyDlsiEm3PL4ksTq2MRH9bDctZgdGGmcLcN7ne940F8o2OnOFnaEyJx9X
Hs3yMb0jMKq8LxLzDC6wFBlVzNb8aRS/VkTp6I066CotAkCxfbnxrjhV8Mgr6Ca7d7xmnO5FfSRG
XP9YEu7BBCA/FlzjBKBGUcArAav0C24NzmUmcacg787PZmCxFJ+vf5t4cghbskF7vV/PnKeSOsM2
3LsTierPaam/VwxDZZr0DAd7gJPl/YK/ofRRis95wdkqN4TsJXu+gEaVKdrSQNy14arcfGPLYgEE
EEdSfBrfssclO6Le8yQHbOF38uyTG/8dpxV7tNn5LrfrO3XrfiIYoEijZlweZNCobhKW0/49BW4B
yhd0rsWdx3CgByqiAqHeNA1obR+EtCYWGVt+eKbVL0pxQe0WiwqnUT+FtEr5zdXnCHkf5yk4wACc
TLdY3p1m98dfCWTiQxM1ks4Rdi7kLW3CjsLx6dRjswXEL0bCOM9lWjtWpRbQvzZa0YQX4/002mXp
9L9n8N5FoP+IK/BnNarpQdlYkEmbS77Ehr/9qrvEDPSpxEIRlgoQUMMrsUiWisTfv1uYEm2uFyVN
Eqa5gilDmwUo/cxzAvDFlHCP4OXbhyhd2p4hH2j93gQDbNDfGrdmlwBzImMOHH5tvI34BaD4ZNzy
Mb9FkbLOhaWSvaGoVY1AqqVkxPYYqY/0WbGkCrsRj9Nfg47QTz1sfo5ixL8U9Iz3zIUfoOogFPL9
eHETAtVqN+Vb90MWmzc1tAEbeG3FwFZA9vxJuzfm9XHe6gACsmVt8l4RdN2bB+IfOK9zOWHirLPj
F/HY8ATFtpWNYaDyHL48LzFCH0aUDfbPpIfem//mmpsei7AGLSMoX7VaPmZhtq7eEzHwC5p1+bo4
meWTfZubPa1yfnyFt3TbuZDcASQOzIh0NsPseQgzmrWiMJPMxbI2WxRDkQBe40Qp3rGYrhAXkQzD
0uoJnY8d6mR5/7ZjpxBpO5PArH0kbxgmwcJx7LyxkSejiMctS1HXcydb9pnNCkHoNC24G5GRmNfL
Nxc8gG0GBKain0xaHRgRzL/k56mXDV1BXu8wLuJNGxHEMCw0dEIRdfWcIwJuRO/0FfKBmPDsedWu
ZfOvY6liKkrgpNdILQVj5sgFecHfRrbZjgmXzOKCSF9a+qp37TAs+tnHfaI4yLUfpfibzlqJNvos
b8adWldWfvmuRwMrhx6o9BZJB4XJZ64NLNXkQt36NoLf9uD9UsK7c3/gIi23IKkGy3rw7KVeBPoi
OL+4cw6P7maiS94BSYoBURCMXtF7apyLsx/tRQgHWIzDFh/MxMz4RM8Spp3trQEyPw/CKL/kTZEF
CLwi73vZ251MERRLXn7UZ3dLEgl2vJ7ma06H60T0E+e2wQauuU1pNGrmfsOlhfzju+74n1eWC9WX
0yhyFnWjHeSZBoj23hqtkAErVqmbEAwO6ZbHQUK6AYpG5+gpJcpVHBnYhESeE/PgLAIQB8tJ01h2
LWqB7pcpFBvCNHoeDTnw+tbcQDg07VnXjsdYb7iNtgn7jcV1xXyXs2BZXAXTl8BaTet6/i92Rw7S
5GGw4cDKmiLz1/FKkLskHN9NHzDazyZ0XEKTG4aPctv3W81arMm724NLzRZ2bR22d1gpiaTefJiK
xrhMGinakP40YLTyWNhXz44/ATPNR30HmaZWm3UXui/MpMyRlIikxDRytRnlk4mGtjK9rGJ+QaSW
fcCTu8kH9oaHSzLCnoj5/rfr+Sg9FbLj3I0GGzAMHWZUgewYjNdW1e7/LqqgzXHfJCxV4bwbYzbq
O9xR5JchNORKeO8b64055pbZQvZd2TiBWn3jipafE3dEml3Vc8TmXvd2Xuei2Dsqd3UeVNOzQIS5
CNArDs66F2R+RWbZPRWgXx7SdwiPdupSTwts0ou4eNxRUk0xI93D9YzVSxABj7g8G0j57W/Z4mPw
95/uJJ5xoH506c2YDnxegEE/62s4tdqwIBc8tQ3LjM9DkeqqPNZEpBHmJv60UYixVNqGoIdoe1tq
zLm0XTkzOmzFXjQjsOzTXhAyMbr8qqrr3kaIYCf7S156zNaWB6WWqtLv4FxG8Hb8a3Zad2nE2lIT
/K5H3S+JSCsLwwfzHLExUOIxCc0fXFvfqyZroU7r805S+adKLiKJAQE1zAqxMybIOlfBUWpcaXIJ
n5EUL+hbgRdRqbhRGQK6gMjaIUCN5/Cj9Kx6hHKQiomtW7vPz3VtcdmRQM+JRhjVtGYOm0t+t9NC
YH4mJv48po7uvfCa9T4doVzB9fxOXBNuYKbuoOZYpNS7CDXpM25ZG8BmpBL/C87R7RWBWeazyQ5N
WtkjgX/RJFJ39ckUtGKaePNo0HJl1jtcjMNak15YhkFQlLffLRc+k066OtYFNhrnTfouQu7ItkqN
u7GQzHDRIJN6uaHZdXdsEgPSIuYSMcu1qrIJ0Jvaw3SzR05Ugy+nbnotbCKqipPbDUiEwC6N0XGQ
1N0Zlex7XicHNVD+P18ynAIYLJbTrKJn1+bWn/NPj8lFOk7xXAJyVgHoGGMi9vlId9JL3cKatR5o
F4mYyCR6mieJh578fsvc858y8fq2FNjUFLkKe8eKeW3YBTpjSVz1F/zp3x03ham75g4GomYCxfHX
dvX9NSd/P4Mx6mk8CmP1EviukO0Zzre011IebqmnC2+Tb1vLQZjostyLuqJwNw0L1x/U/DljqA7U
nRqhOyqpRVKPu9aGwimg9KK7jT7Z+yc842hAm2MlXWCQFqsFcVeuYC6upAZ0mQX+oRNxqtdJGu95
2VfZHCh9QSWINXA86dnLtd7BPAk91OBqpyO7HAbRhIcM62hl2YdXjWy46gZQUQBumsgOUoXglt9I
p8uKQs78avcnACNVHyDfGZZeEi3LwBNbi7MZmeJWrdweOmeG8Q3YPNX07ES6P8xcoIFdP7yz8at+
GgECw8i7QKyhcjEdqm0emQdMi3Dq13w6w9yQMUyNYP4JIOX6XIjvFBzlfEtraG+WLayiSrYO5/eH
eXeOGadfO51L79uivZ27dLqPAksp2iPj0xHygCEfzlBwSioMHwtufQkZ7sBqYHvFXao6Ud5SpxLq
OwRAo1uPkrAaXHeTRwniabjSV7QjkBlx6Tl/k2bFODEDeLjzSF4oBnV/klXApkLHwzrjNBGsVIgm
hDdnN6oL/o6m7BvQOcPIt5il4l3ZvWIFY3OSrw7AGm3PZ0LEQlxV5Q2poaMmacNHabemcmo9wYHT
bhbqa7FDDgmg8nw1lpaQnzXaTrd6TJkdmCqncbwMyEBBNTTXyPd6EOGZ0hbREmIdNnCm1hlUMGHM
nzYT4SCb+Yf0SU5Z7aC/Z9eaHmE8DnGHZlUFXOPZUlS7UTxvFAYcRt5n9oSdNYpTOQc7mUcCL52F
HU8miBFt/4vpE75v2TBuXpl0w01r24cuf2OiLGKrL08MQqW6BtXHgxT9NbP1Dx1BLomXgfyahc8c
mwNFLwT2z+zfRNITsSnSO5ES/OFxxSPJlMRDyYfg/2unb8voQ8vqK/kzaRR1XwFOH8YKd/UKcu+P
2U11hr2HTkrrAGWu0WOO1cNT0r1Ik+4CinhdHPCx0DnzC9IHY8CLEPKswTBBEX6w2cqGo8X58kiD
P+Wlx3x1ISvbGvuD7wfEr4R4cW+BoqErZubFzaqY+4BlY/GnrXz1fBUnK27q3tMeNcoCAiaw1yZa
D6CHRG6iK4Zs21VGFn675kQakU8F9crEU40z7n5WaQAwMknOPOR6osENrUunXiMEfzMTmT2Cc3pm
T+4VX7yNhRsfCE0DZGpuMqTtidBelVSBbSFa0HSNRqcbjqAhN6KGbcKFdDAkU/1eA2qxgu/ZPqjH
6Xzu/80IRTkHSIrLHali6h0lsxw7yRF44GAcPwnkJOfESWFOUaEG8Cx7r9VNlZrBMIFqRNFJ+ktg
wrX65I33ilMaZrN1asRAFrCqekDfC2/UpURz/PFv+Vv0OHuG9xEJBXAVgwKQnbqxzINbBahfeSPp
sei1j8MQzzCa44z0gxmRiYgzXmFKkJGKxff/9S+mxO0tHSj8dNB4OInk2IkqE8mLD1TZ5IiZmlmM
KCBb9yE57nnj88ZM5Q5CBUEQwkjERV52ezPEMRklbZw87ykCJvfDrAXmeCSk6DG2elpf4cgJYTW0
moEl6wSkbKPGy5dVWbrOH3T5cT9jloPOlQobLGBlpAIhJ+rjr+SJnUWSiSN1MpCTqoyvCljLtiWg
PYyOHKWZUAoqeVnK2/AhTDCd1nkeozTt0Jvsu8o04sbp5MH1eDsy6iSH3P+dKDEjlt4v+1PGtVXu
SVYgLoEd74l3lsrb4OsAe/OmErKcpuTjwkhhf+eOXXhHQ5LMphl4CoW5dMI2IIYnSZ+3p/42vM2s
AB1nzLC9L2Tl08Npu0XSuRWpUqcRHOq0oULP+O8q61MvDkRjCRPDg+g7BLtV1uGkT8IG3NkR042t
F31WCGM61KtSQRUp5+uS3K8Jm5Qhw/CqNb2mi7gk+RwHrJAsLWIQZiLkYrjX++VhVkMuDzLrxrot
9Ljwkc+oEL+sPadQKyVu3KXsPILZWdIdcUDsRm3tTX5EL48mQAucZDD4CFLxh1sGyIfkfSUNbzPA
6O4cDiPT9STBMxWid7MiOnOKMU52L7qeyBcAgiW4qvGDus9Vkgvkf+8UWdcKpJMdOpKDNi50rHCY
iTf2ePfLmTDrm4GoClPLI1WyZ+cP0TJRM+X32iU4tv2gwfxPKTeK2gSQ60pmkROtRoV2W5AxDDl1
07WjELr99cHf0OGU62M7o3EOzjD+3mu1uqUsBq7ylZmoSRrd8CM1ODXfhByeaxvOKnyt9JzNtWTH
aVrH639yBWYtW9X58BhryWRdfYSwgTtlM5jTlcMiK88j6PY/dPhZr2OtqjIWLiAKcU99LgpGsyFm
IFfc4AQz5BhmrAS9c5JidAfepZ80Fo8UpJO+2uIlRwwGNY1JaPTlxj2zHdwaY9O6YOwrDHlUiTXU
nY/Ck/Kyx1pf39/4XhvUU6Mo0hehSXvIOgjUy0VX9DZKWoQz+vvO+Tuc9wPgGsggO1oWlYheQ/jA
unzWa/guXgtdMT+wEpdtnr1AOM5ytko0/XgpWE4/ruWprbNTNJcdZU464QNfHFHeew09cqO1ECyz
9hFoHlJ2BpN4wP4NgQlVI/ZZ/43+FmPiY4VsDvWnQ6U9ae72RX+YcIDd9q34z/2mUtAakkIPjRW2
wQDdv2/W9/BOolEctwfaGY0L6sOqH2KT+Wf/OQmMxqlubk///mKZRemWzkq1RnPzON/halAAZDBH
lmtBDO3LEqHmDS5nQVQjZaDK39KvVbEgc2ZGnzR1Z1/QOX4h/f4CCrVVvddA4tDm96E1+1Z2Lhim
rREsHFEybPwjb9/JGxWF97bmVY9Q/7Xi91Xe96FId1YZ1HFdSZdJ3r1bX9u5Dp+fPQww8fvdMWYs
2bAxrog2mHgUaR81EClS1gudBwipajg7rjD9NdrmZ3tuVAAoYycK6VGVku8Y7Lsn3sS9Y301UHS1
DA54FbpTkymeIikSA0NH/gfsftichAcNfBr7S/YQOmFVGgATGyWqAhucEJYSWIOozztHBCvpToNk
7G+znEzGL7QzGTlkAcfpuNirizQOSHB0kni0OYW0JbX8LOXF3Rq6lw2SFbBUpt/HIChSbmBq0ejx
804d6EZoEERuyfzpCaIoS8mmYjUSMrZmLO+8mFx8joDofTzao947wm/bjjONE3VS491YLMwXFNSa
jAigllVLoLoc8VgqEwgJpN0HqKFWx5oaz2PIkD0QGtYobvw4VryCcLnY6VAdeyi2KWEr+8R+oYqy
tN0yNEhK5P6GimnTFrHXLTwMdeoJXqZCZBUWcfNX+Uchqv3+gn2h6KpFDZRNQFmzZXQx0o0btVDO
WgQ4dH6C7GALIq54D8tWJIl3cZUyotg0Wj2JVz8HErQWLeqmidubeeBF0vEfM9gWg2zDF+bIMKHZ
ZSs0OxG2smSzJtvpqlyYdmvQlJVN3KAN9nRR3n6V5ed8ITqv1bo78MscNe+EvChKXDsPehZbG9Y2
I/PYmq7+hoGkpqTboOj239JCrjbm+S9/dEs/V1yiFQtUZ0grgvwpvswvp15BWszLpMvDhXGUBiYd
7rno/f5vmysQDjnH2pQLIlocWEHZhRgxhdShriPznAsIqHxB9ecsf45F7VQmHwaC7ttuk49kJQEw
6jxm8U6RR5Q+Lh5jIT1zR9IFZMU6N/fhtRCrmGnhXV5opcImjp+YAyUa211tBn1Z8XDuti/J0+i3
Xhmqsk9krfDatzfjZdsymLt07mNVLJb4qUy05+33cbIZmgTkdCKUVOUGAiWJlGMde3s07QvLVtOr
J18iLw/zvefp495NdombMg3QmAk62re/IH/XpgtTtjVXnjmAx6PGOPF384jq+ylIJLIqzT8qFAPB
7cYpeJim1+fL/VB0vK7khrOxYtPOdrLbYST1mCLqjxNYuDQ9yDTSOEnVL0T+zESh0gbzi7mraRq/
F6OiaTsmss4KW5RmZDyzsWPDe3LpKl0KTk9vaITiuxww27RBNEfff1QlWgaE764hof+l2CmCBB8Z
VH44WIddpmGuQbwpz3to5Box8xPneJ8D5CTTXfAh/Tv9dFg8A+8L8/7p9sauwuwe+LLy451VzGHV
sICPq8hzLQgCKFUkqYx6N4tbW2qASA+4MiKauhGkrNQmT0PAY+OCAZB/l07YKRWSZ021evkUIUEB
oAxW0wmJSxJZsq6z9KNDFrHl7gYeW3CWMMkA6VWq07YZTNzjWMjG8/PPWWj/fA39nw4GDHmnhaPo
BRWOpx6shYl5aoiueKpdvRteIGzDtUHo2IbxCgU/RFdyNXZ43y6+D/doYr1CiWxlW6Rx2g7HzpJj
tx7Kf/G6GaJUhQAYIZqwkxUndpKWwm3x09N9sS2/79+iAVdSfSvuwJzFW6xNDV3ESX+G4/20tkQX
vz304DwIaSoBcDkOdDQ57roHZYJH8Av9eL2wXGH8nexWh7dZ35WmJ8muBIe2c6q4x9GHeX+8j4CA
yZm/qA7RuNjcGifZWaHzU1e00JtEGPQX1jPdPlgd4kb69i2gVdqxiRheTJKZTbQpi9kk6vMn36y4
MWpN+pTATz2eKyxeY+4/9/q5Janok02ItIukngwJMKHIsKN3ts1VJeeYh8KqWHuiOvQDf+T8Z+0X
sMPbJcRdpSb9pi5J8lS/oOCepA7OfxjIFLQNPVTqdA1mnMHdozr267WQ8n1OvPswYgOafxXfmjQ2
2wbzSwPknD1S3onMpnQcBlVbhPic4+8lx6aZ0kT4iin+/akpKhst2HvzEMAXYigeiGgWzOi9Xaor
wrsehV71kUSuwM7sd2dKs38ecyIMNw2tkyFnh4ZqRUKBYaIY0jO0vl+xYqWwRjhRuHnVhYUbE/96
8BLZpTAG7MgeDuv0Gd31GZKc06gwemak1/yK2nrPLV4pzOW/c//MM0vomnm0XtePpRzzbqx7G6Sw
zKbK14shjeuxi7iPvzwNdbAOqYuKoQ5j1xIiwax3FRm6cRG9NFD0lOIC2QU9+iCzfzuEGeU0R+6v
/EhinVJoHYZWwaHUo3BhQa3SqFOqsJzEHQ6RB2Bsv4B538nszJIJ1npPfnCGK3bO6pfqzZEH28GU
zBeh52iDOBjOpaOaGKEclKTO2hXPiju2BYOKIaEDY+L7Pf+GaRf/H/jcEGEyAMzWY3wMu72Pz+g7
Jvpb8Lhva2kZQOVLNxEDeW5rwI5zX3wSv0OfhkIJCIBTe4ckGAbYRSsCymAWAQ31BP1VV0MZ120B
eVblezxAGBJ+Lk6Ae2bh9Prxnd28qVVH/pshTgIH+nAUsssrjofoaXxxK0Ie9SDr0GE45orObA6w
edyP09NLEFw8maOeAkDxOGH32LElNgvOLjEVLJX/3RIJYdICWlpo3ApN+SyYAVDDM5mvUygrkzMt
QnV8aLDd+JbHZPeknuUhRo2z6302rJg7g4+nVPjd2z3HZ1b6maZh0oEpIlXQx+Hy73ybico44NAb
hnDTkXkyHgDZCbshlk8NN5qSTpK4thbOM5pQkf8CjflEcv8VIgCoEL3HO+ORMEkAf3wAEQbKVVHI
9LgQiVtBGgOFkkuYh8XQFKrj7+1TuEtYRfw3w+Ld2faDy4PkMZl8DXrYjSU0/lnZby4qDx5Ub1bk
5B63MpMdEfom1J/3HC/fBh/SCar8Tmv7WskPxtcXZxj4LhgBQH6scRAuOVuuribDOnOwFoV7xyGw
0BB+4aUZE0MMnYFNZRO/AZ9Y387Dl2NUodzWgrQPheZzHe4JSucHKs/0n+zLQ9oBNehUm/YuNq8G
SN0gEmSbU6obUBoPSmbgHc0p8vEzIM6aEwUTjZy/xZy8J5fXKwhRLkdSmiM+nV/uIbwtTTrSPv/+
8EsEPKqtybECl/NuPhuJhVaCyWAQCCjFBLwnsCNxyzmfTINSiJqiIHAbiWkW5sKcD+L08MzF8/ze
xTAdVH/4aTt0A3Kk8O2RBi742mvXR4yHn843qBHVHXSYw8/xY9fEKkcMquNVXFSN5sovvPFs/ZEQ
cJMeEPDhHHeFDWMQ4e3s3jNMkMhbDik8Tg9uno+bRBB5M1cFMKaSpfjxuUT0Fd1CuRii+dLVb1Os
iGUdA96SY/9e20xFpBeCu7g+Bk492lIC2J2Kg/83ZU4BkJn4b/XYVyFIBibuZVTWR7KqeVc7pqLP
b17nIls8j4QJLaKJmnHRF5c8ZrKbJ/hckpKpHhtThQrFYf9VZ2aqsdjSs9fhoL2Sy3ZNJNUORO7a
rGORPfOXp0a7secPAq8RnGLO546t5akWZFAZj54w4PzkcEnXTp5TVgXJIDwaU/uaOwAMdB1Asg/M
5G/J/ZGkY04SiIM3hX6FUZ3XqS9ry5cSbfx1O+nYQ0KnX3WbLW0Yf4HTn0RYlNTuPGrwR5d/QZ0O
Mx5JSpjZRaLYxFUjVqC9EM9qaeN1Un9mJc8mho4wPeQLQD+sXTPf6+wsedLLVmqSBLvwyrBYvd/E
bzXCiltYHMVBWf7XKKAO4TrAu87GLiDrbgB6A1U3rBgkCJc3AtlNw7gkwezkoRlHsvMj4o9VR0Ii
FhsBJ0THMW/A+ulc/t8Ozgv91xutxmbW80KWK5nXJpCs3anK3MWPVX5h32NVNOBw452+w2ZyIv0z
iqZN0AEoFG2ZnQXtmQhbEvRM9JwYUfvEvqmvq4KM9KPQByVtgmdVwWXAfTpdmIjrNZ0QnU4LEmoU
OytRSx3grByJFMTm2Zuq/CsppCb3Et9Pln1/v9GvNLcigGIamjin6ERmoE1CbjCgOmhieXH9Z5ks
7NqB29VYvi18Dp+MHjunDpmvXs0rXcw95jGG5TN4YqeZQi/Wv+MD6B2frGtx+xwFD/RYNezH1FFU
5eIEKLgzEdXMSnOQ5167mjr6W5WaOS2C91BceMj15LPT2CVhJsEZYGQp/t2sxFG0Yrf8YFWOczpC
QW4vmFX2yQ44ZnpQBCo/P/dC8d7164St+dNLERz65Lqu91ebmPKl0L26oPGB33PHAK6xiDsW2iyI
7DrUBVNg0pdT2aFkZ2MbbU6EPOYqfR7U/8Smx8tScQKUoIWFtJD3kfiKzXbkbrDookPpgEymwFee
kbsKh2xooUCP5dQf1wQVZnJlOZ/Lc2t5wwNKoTTqbfKcrRrPrS8nIUyJ34/2SgO9eLt+dsLORma3
4IkQw029qCxOMy/5Jj5TClMKt0w4Z4CgtfEOelTz68kZ2Zy6BxL/dTS/gE1lGc2+PYQRyJ2lVCqx
qNHS7J8fEZLQvNeN9hsw5LSrEnxrTNx/Xv4CfeXCNRVUMaft7CLrkV9VSJfQKqY+ZSeHf7TPXROL
O7dhHZ7+6boiypIon17Yl29qCP4+1kxknFsscS0w/xw10k1pWgTY2MAoQAYLcnNPlI+tWvtuwgh3
09vou2VgYIb6DYZwh1AIjlN6KoyDxZJjx0fHTDJTkR/DnXdX8oKlw38+vNsyJZV/IxhdK5v63Yfx
TxwRIlwPeOTQPOLe0uHIC9EbMMv8e2fYCIn/KBg7PIJf2UMFMXmhncaynVEaOMPh7s/ma9ebr+At
ahc+uIzstthRzKQrI/ulP1YUUYZGnIo6egKo63CnfJbF2377xkp2VoIMAuwY5dfJjkadX01K4Zdq
Zuzjacr0J80aBtj7w7sqSkK8LVdpEqQdkgDtjydEkkOz/Yr3ldyfKLLru51+fWKRbUNWHn1FOLNI
9R/TF/qX+0mIkdbAAy/7zpm1T/tj3RL5oJfcJyLG5/8GR/Jh1Ne9LAlneGQRxDVwItrMA1hjIszX
6ovj1F9CRcUywmmckJ/RC/rLT3OMuv86aJK2hDjJTegYPpZ/H2LGcs2NzDe4B6xR9b8DcWiXfY8w
P0Sknj5a6DRy1Ed3PiwDG+PGYtN2/8bg3axRPOb4oxo0zrjMXB5Iqp4vheT18uXTOKGF3blJ8aYj
dxfHnVHKQsFYpORIrEY4SJngzXAZCiQnv3FDYdXNMiOXKC7xxMSJC1uUHWXQHCImC8LzwOhdTGvb
+6p4AaUqQ6XW1Bw1vEGkVHbxmTQ3JKAlrOP43Sn1xcyJEiq79gz27XQYJttAEr+MfYwiQk4Ylbx1
eZbC+rZhOPEL+Drv5yj/XtpNF1m6/WzHNr4yoxQznHP6wlStD7YkQpZG7+pOTZcDVcYylGa2lK2d
X1WInBDMR13MfwAoT9FVKL6hQOAHyEAVPcL3Fn/6DYIYW6YRr9xu0z8W1kzK3q6z/eZHmti/G6LA
T1MMQoQdL7akC10Q/l7ubvGGh/ZKl+W1SnExWEOfyTqwPjQTdLEjc5IYdH2Jgbn1QjMw+TcDnkUC
gIuYHvegAARYg7tcSyp5m4BGmOjZq5aavO9/kEyj3DVUdOWtltsHYtF7UhrcPiFfAnIStnxMJ7wx
vh2ysz1Tijbb4gn1Cqy5WiDAMpubKk1XPl6R47L8zweZXPAIwuydAg7np3o2Sgss+Y+eVfQZkW4F
5x6PVY30GomY8AD/bDZZgUiQHYqdHwmnW8kgeDKxLps9Q1E0o+Ih8qrMT2ABRYgQ11Ztk5DucEQr
uFa9npkP/DgDpNi1SHYRBEoGLYhqUhX5CXeK6s3I4niFkU+9j5Fq3ZP0PG4QsrNgdMoUeo7xz6Ct
IDj8btgVYZCJPT20S2b03MF8xaImAGFDVYHr2MM/syblTE4tUhJifDkP34m/E5cAGWBlpeuL8F5C
W79qTkXR1DfDYizbCSY/11qF65Y+Qm6SJ0Rm1KHLPWScxBU+BKgtHffVktxY/ntbHxQrJzsSs/Pd
cKLZM9NIo84+7QhOWfNaYqxZXbXSWH3lv3fWqa9fLKhoSMqgkGICrTZItq9vxEG4S+WEGaMpeyp8
zv23JmBJRyuZzebTG7OZNl+A+v+paxVtW5REKAV8GDne6v837RUSej9an0e4JIl9HfvhLUyI7DHM
vhv8QdACi5qeHgteHxfs1yFEDQUyjzde2fjoSEcV9fznvfQZdymeXiIKWzqVwxDuzOCz/7qKc4kA
7Q28txmJHF7xTq+ARkVAQ5H72hqyXM/V6AvNHUiM1xaMJKigQu3idvM5Qbl31vtYuhw6+Ki3r5PC
EQriYB6qPdM5y2HmQIJ3QdTEiS8ekUTnq5VAFXjLkW0JIdeHayilWhPO4/XD+M4I+8UUwyNI76wp
hwSdg9jIP9e7AnrV1DgtIw5ZbiKuoYFOWpOxAT8SzX/pL6HImVphmG8YEsEaAiYkpa6WbYVHOIx5
P9cIAhQ0QTDiyzJHl2xVkgcE51Z8of0R79LEWPEmbrsi2qQaPSIng1MJJHLOeNX4V0zSgIwkzU4L
1++rJhQiDbdc53uCf2+tqEUzlUtBeK5SXRdpmNetqHGy3EK2ZM0CwW2LQHNgRDMJ9XF8gnWTX5RH
7fIgsfYOKgwKviMJQtOyDH1v20NZ6IcnOpHW0u8Wusqb0CaA1GQi/2p14/0tc0ec83mxU4WtVLI9
GwOs0WxUJp0LvRbpxr3GX7nl0P/ZgIdG4huehaXwAcHZmzZ0MERDHU5wMcLzFypdKAX1taUijh7+
3VIXNdyTQ6emnRLOPzFHrFp5fEJ0gF7plCYgBE1sM77ug3IOo49Efz/LVfb5H4TGEXec/lfzz3vh
2h6jv5s0hoHh87udx8wgkYhlLVfIy3DLjO4hZ9y1h+Ca9ArodIFaiOM2ntR79GhUTR8InbvULQQG
n06E/+pRjUriyaPW1LS+YAVhSSLCRrz8NNPNzxzLiFEGw9vUbSOXJVwU8UwlcAXovKa2AGjSV1uJ
AsJxdDY3e88Bizifz0x8/0mHnnOtQB48ZXB79vNDLS8/Vux+eTdCMBLCdI6CqQXKhkk7JHEN8Pa4
x41EfAAhl/qq6kpMjGmh1X4XvgEwfChYfjyFpdWkzfllg55F0XVTXtnM1pwE4a4xkk+SfD2raQ3E
RnvJhrIRFXHsqP/t8peI3+dyOzSaW2EFPacDmiYavJYcIoCIdaxjzbgd/S1imRjaWIPmcfDTPzyw
2Uwvtb83uYUfgOs1oMBrV6LefjLYa1zDsf3ZjY9wQQT4b5XPKraVAU6QVipSC6SxQzq6baXi01sq
KpzoG93zexCKtClIYYuWCDEP8mBV8zot1H8oqbRco6DqGa33P27PQzz6b+M4nXt+AJD6A61EEzzD
om6hBBXEcSN01bAJFNekls0snh6NScfMLBsvisp04W8S/Wik0ypY57UPfq7owdQyis46SP5pGp+2
30pp8BFGnfqtYnS6qTIQWDPc+0EokxZSjXvBXe1vND8dmkbq1A2Vsf/NQTqfP7ylu2ZXgvucPQYG
Wf6n9yM8JyBTVg7hjmoF/KWyK56DYh5FCmDjuGgIpKZnCnaQRPdhiEEKqzdmml5YznHD/uMrTGMJ
IFi87uhxbSb90bmjFJaHxQi3cT/JIcJfygbUYn012FncHWAOQ5oTEJYKFdpSpHvZ6etSJg75t3pp
Nh7gUgXOLHA311Ph61FjlccGHcbrVVJ9w7+dtghqpSFtt09uUrnHT4upvlwCNH6UJ+6ratYOuk5o
JhkbnNRRM8OvCYEEAqDPbKTH0FMWiBYnq4f+4na1dluHTWRuMwsGbM+Dd6tPz8CFbSKD5gH7GucJ
ZvLR9UhurWBJCUt9IWo9TKIdBoORmzrKiaaSimxIxkOCQtLnWukI/JYZZRZO+Z7u1uVfCNTG8n9D
Q+q8XV8AIr6a7W+9BfksIsw9QPFblGzKkfkgHc7RtpbOSXAScIGmYJGp+02GG67CudLZG4beEy8j
7eGwT96moEq53R+/ISvYwVGoeJSr3wemX469eGf0hGueY4k8CmfSQC+SEsoA4+iJjR/tNlWDK01z
nenn3M/QVgUFVjVBTqJGspvnhMEXlaDpTK5NN09W1ZEmx4gLleG3+W50SbzULYYFRcTLtU/YCkpW
9PbwNel0Ucgev6jSHW+VR8wrJahyXC8+swivE5e6++RjUrFGpOrU+slOgJgc9HKpok9I31CEe7Qi
tgto8U51UewqPihZ02tkhyySYgR4HLTsVdZ17ZjICWNhbgf6stQ6Pp+D8bg+FfoEM3qM0KsoufA+
m/fQmZmuTK5ZQrd4gD0Oc5ZJeIdBjvQ1a0KVbdmXn6peEQKF+GT42x3CaHqNYPsD6zATSy93mn0t
IZ9QSI70/MN4h/iOx7YEBTpWtVW9u22TvAUY9RLVIMzBDCdLoeAduL0zJK5hn04vfXEhSN0CBOXB
kGkrmqyLfvBZ6g6NpNLsvBJqUH+9dRmIsQ0aause+lteSlyDEdP/C+HcFKeBcIyQ7makWHyX/lBX
EDCY5HTsQ0iHxq4/TafIv15BHdgpSk0glXaGfziAikqQOV5HeuhEvEKnnrq1GYmucGfuKqbrUdFB
9TN+hODpX0SQwrZOt2ZzHee8XnMfZvPphXJHTKi1kvwTuotNbzkwb+pMytLlyaDkcGAhxq7O64jU
dOzlW8crOGdEk8/r5JwphfhjB33NNHv1zfWOEhL+ZNvEJQOspjbx8054IjgSRWLyn/BpY/5l2SK+
gMm//xhMM2fWPgujdlInp71VhNUAR21nTwaaJ4d+Xs9wiWO2PBpaLDK7wW5X77OUuu3Loj1SsCRj
28+h+23JK4JcKqhIAC1zrtdz5i69Aov/QRnhW2qa8dkPvOXfRP5uPSP5/ff5C75wJscEAXkvGgul
LrtTpHQTFB4AEO5sMZ5YPjtyBiEqofIFAKliS6cz0u26Aj3TSLoFhAh4bR3Q4Sx2XAkl3iyzl8Wx
KwaN7sDZdR6BnNnvMnXzGqlOxp1kxkS3WGO7r1CcSAy5YGKPOdVFiACfiQsCjPXth/BCLCXmbMWV
3FrPmQ8IoUJ/47WkSqrUMHTKLVBFXDezt/diA5hsW5Wt3tGORIckpjrZ3Pkv4Z6vyu9ctB3rHAYM
WUmRfTSXjc9u+ynDaaY7YeGtSY63nGNhqnuW0MbjcGk+wb6UJKs+B5HESilB4fSpkXlbPJNaXfxo
gaCkXnhj08paXEEAOeMk03uGCx0H9cDl5/nlkl+vdqgOMPfYwJ6jk4uq6mmOUxyhHiJ0bJvhKrYN
2xgQYxmC/Imq2rdOtnuMRUj/MM+2ej8RUbE/yXAjDdhSth8RGb+y07bnxACe3GgSOsbSToVtjvYp
tJJMnmo9biBVVZY6fMoEH/x3tQ8e3RP0Vj9KvMjkTUKMEuaFTdZDtQfQrtov/Wxx3Nh+YR72w/Rt
wNKjO+hnxvY4hbH8gwCALjOD6BrBaOdeE0gwiRa+HwJqljFeXAaBQhvTkvALae44dhb8NFKTiiMi
3QMa2Wgof3JkZ+F1g4zIbZqq/zeGCacfBwZtFEGH8bRcsYU1OTa6SouvYDYRy6BdKJNQkCygW3qB
ybK18n24dKNXGgvbZrvzzZ+VWYu7XCBMc6SpcZguFMDdoMevJODY3L/EsYK2HKCqQVz8jlQvfYoj
qcmhkqO+zEBwYxxypyCe0BWUc4psdpiJyDkMZBI+IJ6iQxBAoBmsVMVmkEwygaZsxcMUQ+PXLHNV
CVVbws+lGprR9Jxmi/G6IQ4LLyBItOuLIBMLdedandbWlousmWz5LQUazg2hWUkBVx/Gs0KPnAkZ
NfDMTKl6BdXND9vDJ2rER/TlReJ05o+eeQ61I0W8dBotKmX4tLrjf7RyRVI2P5AyVX8+rwKNpr+Z
FvSZk4F081I+fugTjkGTrmqr5b/E/e0McmjXOhqeJyE7GoozAAk1WDUJ4YIv8g/WW+YhN9ZaEDVX
X+mwDV7kN/cgNuaQJXN+ZQJIHjPf0YmNkgwFeSUE5PTfzOargiq3uqzTFQKwRVuAgaiP1sgu5S1o
VqhQOiw/KTKwvgr81zS5T2MXE+mXsBz0evv98Wnp8EZmtSpmMJHD+YxMBuzEVXP6+fC9ww4fzsco
iDrRw5OVLfEjdlLs8xKVANiHRFyJn6/tUwZTFsBrzFiriSif/EgxgSWqBd80L7oBZEk8SjeyhVdm
w3SBUVarC23FbBTZ6jn6kI1MuuDpOVcm7eGhpMDVhp1w2I2ZJcLlxbJkUQSfn6i1ON3KRjMhmB9O
jp+mGejcYoWT8ga0TKeZqdpoxw/mZSXqncFdCqwWGtC1/UktVsMleJWvkVEVuSIEaftbscX3wea1
ZD1S4+LUH7WgtaOZjAZnYyxfQ1ZlIg2jOdXGKaC422ufcNK9/PlziNvbKWMLy3WnYwK34p1Arncl
uUxKPw/h9kEsQdXzzeNW7JlfELzIEubHmyhAjDfRCqBhNTgSTRwyFXxe4LbxvQGHi25L8sp1gk0m
shojDMRHU6cJhHAxVfb8aDg+zXAgOMBSqMTqFlUeLveSVYUzj8iGt1wnqEaW7/AD4pU/xiAAzO2c
fh+q+cm6vakJ/4/tjY5uVfQNv2rju1XRGGldcRK7bvktXVjDylpx5idlOUg6CofgcrPjpO4/ijHW
9Ob/93PGnePu3D8uD4an2rMWMZkJqm/Dy5nnBQTjPvl5qGN4Sg/pgQ3mA/3X9n4i2OPnJNKZcjZM
5god+ranbjEVfrV/rfU7x3FhK+iLz2Cu8yXlJ5WjAYnSzx4uURt5mb3HMqQaa7nSj++tIodgjhqB
2ohcCaknTFt6fgDQh6GP/BHWyUC6NEu5eModnGTx0Nj8Ic9ucZH2b1HuWYWB0QkFxVJIAsL5GeB8
9Rdgie3jsy9wsK7s4CMXpDGEw+B7mxJ0CEsms0n9euWeziOH2M+CJyIZ0PCVQV53ePIIFy5I1rfB
yyLbgKaTUX1LdcLwaWw7usYXrEqLUuFVUjLbkk1vTrQKR7rXIOwWJWQpOTmZbbjrhV2OH1NAOz8g
cTJpI2H5cjr7bOlmyizAIPuaEMVeNEMOYEy/rKasRgxKUmK7fE+X25iR88z12URMtBtpkQ9eGRhE
sHksp3vQp7ZFTKjnrusLF+PKFr5ijGVUhGETT4mM4/C5keKW6EBsmnEXVIjKdOC826O+PFOXLqJu
DUwAKPvBIDehAL65n1lIwB9iW2c+b7xMZQ+0MnekGxPLC9lEHw9RSSXm/uc4UiCi1KQugx29R51y
SKBaZlOCvWI2W54V9Hx1v5NxZ6X1Z7jQ5XmQ+etKiJi+jy2OB7WGyiT3o61PcafvhxskTkJg0eTh
Uf8KbUaMZKMQnHbDEGnPAtx1RZeWog2pij4FUJSUNgdbhG20OnVBSFi+Zz56Y1+1EH9rFMvPbrf4
1Ca7Wfgzu3Rax4e66kl+gO4v4NuR4txpdL+EMwsI8nxTOxYxFVms8QwtfHn8IntNeEmeLhtmQe68
/viLlazVgfLdTfgIxvH+S3vRL7qhspRa6UbB5G0ZWeoKSl1BGn2BpLFqMw/sC42HkYSiiMs3JUoR
cro4U/VcVU0WebBxe/xG4z098kogTpBgdZlWYnbzp8P+VFA5FLEo5BgrumKBlpwrik1J69EyGjlt
BehUNHNRQ5q4QFz38xDG4cHA2Yrri00yVscDftdkD+o/rX4irxvWWRW7UBGw5uw++hWA4Of6t4uS
aQmOC3NCjWnUrogqdQ2bpB6Ezn6QRY2C1tqHK9wo+cQ4Em17zV94JsXrnIC6YXI35mFBevhXfugj
VACDXjlqH1huErGxm9stv81COcmM1HoAgkQu1UNMEBQuAxK3HTXaim6zbg4MdAfXrg1fzfkmmn62
QYuAupyvayrIEpGKCWHrhbvzDlcs7PtPqu/lx3SvM70wOV7CVfxBwn0GK0ZKJ57lZM8FfJ0BISAU
AkukJe27F8hqz2BRAtDDmZpS7PVRFuKU2RPb0/KFcG9fMptdBTziTKaIt7m1F7QQSEu29bqUmgtM
IXiSFgBU/uqhZqlvOs4G+ykOGqIAsKMunipFCcH4hL3h1OA6hdWEZXKcPD3T9SQltV7vReQ/k27X
G4P4eTfmDwufQPcsdPpIGscZ+vT1KFOrZlm5lSB7BCpQdiVVU+WF0SWX/U+Ax9WF72RlouxnJSu0
IERnkVy4bR3l5a22TCTUxci5LFHfg0HjOUHvBpytDU2eFqi2jg3jDkgJbKLI0hsZ+Hv6bEE2FaBJ
j+fPDDWyDjKHhbqSik0wiszk2c2fgWUD2pl27lT/U6K8afe29ZCvkDkXHvfMz7scYPIz2UDDq1us
8NEPTe3nrjOPTIjDshDewpXNibWuWMx+kEEHFUQm3meRyw0kYgzvsZS8tsRXUrPacraXmvI+B8sL
nnYnGBwnRqMeb7FbGdvRTg0DlciWpbo0u89PSHbO2+6l/cfVJyDhm3dx1J3kIqRTt6FRln8GawTI
EtI9zJtPRg9dd/rbvd+jCQjeCmr1SIjsPEQsxf6SJB9scV9pvBIjRwEpZxbtBS1HDDz48EcUvqk0
wTorpL9PpgrtFm7dk/9r/aTLt0Pm+LFRLTGW+Bs0RV2PPqYEwjOP+YKpFhyU7dBabrkqNwUjN9OV
cBHU33WVOBS0UdI0rzyt61WM0qdW//RmXnbDKF5tRMSVTDK4uPbRS6Q/5q3Rwp+cQzTEf68dxmRS
xGmMP/0ah9wlKNhui2j1bkAn1zMCTS9+X1qG4STCZLiYoHa+PvviMp2ePVX8+HwDXTyXM/aLlH6+
dNr2f5CYrADLX2tQ6CzB5nZm+BtmDCORBO+jjQ8IUxYmL57uXRCtNntnha3MK/ypkt5F0UWoVMVK
lp9wwhCjkdMD+vdhs5ohrcOl+0/4+Sh7iC6IzEeHeafPMzvY7TqMJprR008pBJ6SVnvUCwGha2L0
HxutubyM827bhcaw4IG8tnkdrIZczv9fWLzrbo9O7uCtc3oa85pT867k1VWdQmSO4PR/3+DKTy8i
Zx9PSGd/UTbePetkEnrgfdLpTImvZXCUm8bDME/A+9HCI2Rauxptw+TaJt//X2QFhYEwQ5vufATN
ND7VH0mHbyhP7Md0uR0JQS/ArlYtpXJDQc5qhqpBDPYb9fe6wqanxMyq+kXsJA2OsT4hVMhW/D60
tegmiLXyZl5+vscjTlZXjq8dj3hYgL3s6JJYitOOEmhKFuJcsW3JuCEXUTcXUKWXB2ny5upQdnyS
gilp+wFXj9jE4TcKezvhd7l/fYFita8HIpyRKazOEXT/LI9JHUszT/RjhHjzhm/odWI8VEo6+o37
jGOFUqyQn+4r7rlYwn/Ef6wspi84Sx28s5wVPo+GeqIQVEO6eKjvSaFQO5FrZ893yj/gMHGM67lg
9pcLx7Z7sy1Qf4wKTtrR/k1jWjB8sK16HGwoO8UMHSHecjJxlnEE3jJLXLSA17dYu93g+pvdqWoM
OydKli3QkMmUFlzwA28soCGV3fpChhCcVgE9pUaPNdqelY/bzwSInwcKNrisNLrLlIcc6EWkgDPe
/yLXsJuY00nNIPBxC3OzgODrVvM0bNEtxJ9H0AKu9Fc85Rs+HMQpYeEIDcV5ef6uabxmU0wCXJiQ
yRrKjazJCzpoHpTl8UpfyiaWFuGN3yja1SPOA+gRPryOyocVTRHS6BparnoJQAPPEf6ViYrcdzdx
hLIG99I6jc2p8iYUx8PeKmAriAxO2SZOTFXqKkzlJaG2bP0OWsoxkO0pd4kVbWWZ56Vr401OZFaS
enGAMsvx5xAxMeZetcmIRPOOdCwwzcVTWanfhgMQmYlJL3Lt+kbG0+V1Ng3LPlaD+in5xhwE1g7u
Xom9ojZzGttQneW+uqOUCrZEkLJ/FE2ZlzR4xOw5EeRyhyli9T/1VXbCV8jnUgZtSuZJ9NWs0vgm
Evuyieg2CukqmbwGOJ14EzCWnHty+w82v/5C3YmNldkgJqiBNzEBzKgH0NYHSux7tEvVJDWxer7d
Z0hsbRYNtbmm7TmMg+M5sI+hCaTyT9L4ywLTzQh6RM2UVMSm8YxsSNekN8beXG86zJXSHb3+LFjA
/N3euVhmpUuepBgNClFjqtPuFHHKfBzOshGJJ+PjWWxda0lpIRg4srbDFy5Do6TVmTQs9iV+iWNc
Q2byIPvjaTAR4y8fzzaKRHOgM/flk9j/H9I0zzY31SJHtQEqmS/+Hp0ugpReJ0HS8KVkkXQcFK9J
x0EDE2lCua1DwYfYZ+0ogNULS7iHDVlNutmLzQOTNG89LA6GnyFaQUOCDYiLndyq66fZupE+ddYJ
fTmGxg2IqwtHr7EvlbRGLfeePzshjpDe6cVmA8oIqYRcy8Sm7JmkqMdICushgXqC5UHwm3k3Lbgn
VZEh8QRfkyLvQAoDDoO0b1O+RXXqRMZ5mdgr0pShx9ZPynczG/YhAmkI1LvWv9inDd6xH1kfe9yE
ulA3QM5fJNx8ILmmQU74o5T/t7yVQLsrrHRX0lJRSCMIA/LCy9SxBjzuGJfFKPuF/2qgZZRXzYXq
jvRo27eO2OKFw2UmTxIRGCdTT5dquGvZgNFUa2nVPQG73ho2p7cTCwzJwgFuCIeTde7q73Ma4lMF
4mtxGMUVPMs4+U2C+ufxrje8BTvZ/sW9NClc9IRUTFY7RoRlMArUZynTM2tzQOBlg7ZHSplNMXaA
ACmg1dgTUGANvusL2H/hchJoAotzbJW0L+dIHETOMp7TSb8Se8G7hraerinf7mUZ0rNeE8Kdtu7G
/FzxoiY1iJOdu80l5bCkd9Gl1yjZZ5BfvCDxF2D5t4t8Pc7+k+YP8CCNzYgh61jFYmBZfx6YmH/1
59YiDhrC53ypu0SLGz2LUgN0sAN2vWvy+2SHSbQVVpddI9j4f979XQaA+HXOIPhN2a0tYUj0jcDT
hAMpo3zILiF0GPmNEeqRl+IwepD6XnJbLepFn51wPrV1C8YSlQiIHsTbOHr2bi0KUIGLYxd0CbBI
3RPXmcure/wHTdotoCvkYW3eaJHC8jOfr7dbxujCXAf4er3k2oCsC7SjyZd+I+vvEMTc8qEVoZ4R
2OBwt4qTzk9UiNaRqr6iJl+f9QZtDz/q/fyg6hgSbEU5CI+XdU+hI7csfGyHnxe2x7fIv3oYkzsp
q+yPC0S95flTParhAv3rA5FRAuN0GxB7qyPrEvtn05z9WA5B5a9MrlPki02bbUvacb2hrv4Qazpv
yqjDp9uNYtQYI03UAA6xPQ99lhv0ur3TVwRuyL8+IQ9kXTnMLTqmN9PLH8PtdT4tVSPDCs3am4kN
KmOl/fBGoD2cuuwAjMeEKYzN/s24gEonz0sD3vqpvsCmi00Is8QA/nSISyCtBTPhWTdVmoPvd78L
x+jSIztRwnjdMVxKxgsltaouJUzL+0cysR0/tNn5+FpxHf7xQ83JA5COs0bkSrbgGuP3TmZuP1C/
BXo55GNgrXQjkPa2ep30hexaebZaqpWwlCkzu0qv/C7nvAV+i4IPM3+X3ojMzYcDLM8kxUe8MF59
4sAYW/X2p4j4RA0h+4RCL/IJuC/Haf2J83YYhG6xlt7eWSBk5Ii7NCVSSQTI3lv2+iOmJMmmGFb0
47BKXEaHdskWQ56k12yFbNTveAd3Hx5VmE3ZJshhz/g/O4xRygeXpcr5nuFOMiS9pjRFpZcbg8WY
TxWkPVQRAt+sp+ZpgdhyFCn+rx8eF2OOYH+IMY6F59TiXUivPg1IkcLbtVBVvFUUaxroSzoiHpyS
jEbun28u6TkTUNonEE7P/vBohhKO7bX6jA5B45A1hD/BI0FuPV29rpNQlEgn7lCzDSMnZjR4QWEc
ZvcjKLlYoHrww9pNIqW2G8XCtLzkHYQGjo2fM5Vx218WeWH0elAL7R657iDHCxhoTF8aAvYci+NV
igxfIrxzB5MjpO3YwlkeTzqfSMMm2F5Mfh3nGBsw0PjLuPEooTRQr5yiKMidbRpVdvxxpPgbLy+S
Y8ztU/DnJ3LuHPwxBVYSjEexOEamJqrcbH/Vbpj2q+HF/vTlhk7POzRWjlYFkQcqOY69AlIljz8r
ULXbLOHR8KE5EuRdpI34AHNZAdtJWHgnUm8jhZuFOPSVyHaSo5q8QaIj9yy08q7Hy9otwXPSEoDr
KtOBYhLwyGFCNuqMffa003OQGk4L+yjJRKHcwA9Ir+Md64o1UX6BFfe3g7vleMZyMRRwL6hgQCWp
9/qMEE6rN9C270gh/T83kNEtB+Sf9dsieWORRgGlkWeoC/xK8fAoHRoa8DW9In4POmKEk5/d6RpB
jHiiux1qbQ7Z3sWnReCyDWT9Zktxj+Ss4Qs2rlJ2ta5OXjs7fgkllb7EHU/HHpake0SZitPsNCMn
cQLQfKTw1MI1jUsouL9wKUrN8X43lmgqtqzQz/1LD7qrUCVNU4KUrMA6DiOKchFwWh+CAD/JAy3C
5GVmwbbBwcQ54bfLf8KM+EhVGqY49UGaxEr3KcXoJrBfAY7x1B1f4wHK0iR5/0Yu/z7AmHuMJpPW
0G4P3ajGdVUxzzVoPVtAeAetOpHBo98Ll0Wt0wQrv6o4fd71W1zK6YJvhqsh4Suiojzj1w8EjSmP
SjcpAsoncAahWReq0MBS83S/YZ87M9RbASgSYUCvMMB5YXzKg6/p6lidnPfomOf1zeVirR1ddmBB
g9W0GnD+B90GTSR6tbWKo1VAOEc/qIdV8LuIdXC0Uz6mUdGImPsr+yqzfw0YmGw/Gm9g35hKOpZq
ePv6SogSVFW1Y/9PEd7nb13d/cxyVg5E0A4EVkhobouedGbCqF6NxdgG6f3p/R31TB4CrY/ip3Ik
ENtrMV5/YHF1+5b4icHCdbcga2XZyJJ58zRA0Ed5z7Tu39XlEVBKPBNb7dEFhLOMV+9dfKde+clc
CVhLyw27YvYq34dGYsnDFErEH/o6D3iQD2Fad1dej2071AJLQl7XqX4e7UyaZ01X7+1dG3VNHoOg
T+dlxolO3DSx68kkSukTsXZdaz+xDAivO53k6XSGvRawQZkA5a0iuVRWwSGVqBkOO8r2oEDrUAY/
jsjEGswbrYTyXhp2tdMSzqbZNWnQosGpxxx+NtrLhnYjKsUJImZAV+WXyuQ0h/5c1moOkVYnz9sB
TSPziG6x6GgQUrRolSteQllZGgujmIxEYjC3C8Poq428dNS3Oqs3Uajy0LC0OB4tA/x+O2vsGAOG
0ydkKRV+miRixXZA2QoWm47ovuYIHq5+6MfFUMdf6N4YhdjAuMbVOl3UYKjdQUVfYqsjT5pqWU+Q
fC/U1687hM/6N1t0ft1YocWlbktvjyuZyx650BAWci8i5GBHMMEfXn4qvXCpoctE2vYW63QQ6WzB
nQ0K48ZIHPCXecy6W6VN9W3w2+zEeStggkZpcKFTeYe6/hnvZMzkZ8oX5VWLzjlSWhpg+R3sloR6
YgFqO2keaKH0zWsy9pJu+guVBfpsVfOvGCJcTSjXhg/rc1gyAL3X6OKzqNN01rIEk7yPqDOcUj9E
eDa9o0pNC5hZ9Dj9MyqDcfVN5uZCpsGZ4RWnf5GMCA7XhicSqRibY1e1qznx3cS2mfMdsc0HeoYK
0INRMv8EYMDj/55aXP0jTvzwIFjWGnDP7b4GpD/fGIVvuwmFZSDqYXQk/SXy1ef4e5S6BfBj5U79
933vlvRPaC/J6V+YdagQ2zj4xhf28ijy3Sw/1tmL5nOpQcTeD3p21A0e8uxArFTQAftvQVk6cQ2y
BWua7l5d/QoFW4DhG36YzkFmNMoJtIToXCgOIR52aTPRzRXiY2omYF8URK6d7zA6Y/ZmIvofAIPd
YZqRJkurtK4RZhTe/ybTPQ0D8lv4IZcjCPRiWLxQ1XegUHQ2M0877sjpRhGeq2RXAerW8ZTz6QHk
sOchavyV/38BdL0qpW4T0sjv08pvh/o3gym/TT8fjxcB0hX4vpJi0jzqbK95VJ9uIUtRxPVDid3L
kRG+t1z0vvXvmjCtpqqa+ElGR3RE23mIG7qRrtr0WArMV5D2dNgudKNW+Q9Q/a5S5IjMqRDSnKwG
+8iMt5qkYhWAyKyGbubNnYY09R3loGQvjvt7eQBieDpXf+uP2sl1urve50oyoclFmOx3Jy2haZ6E
Tf1+HROB30G1TGYyRIYijivobh0X9uI7jfWa3UOGGaWPOIrRtwAlpbemjQo+72jupEf9MJgx1vzD
hm+Xqrhm5ZdVDWN0zotmTGhtbzFwXpMB5bO7r23Z6BAomDVvYnt0JZF+KcThwIXFvYogb5TvJ97B
wZdSQ/75P24BlvNCmuRhHs+RiDocNBWJtr39MMPIajDsI7DPmR+HXmpn2SSBRBYGkfrLVtynG5IE
VePiRcsnDXD7TBAijxM81y+yIXqswHCiC49tzQ1HfuMhWFB9jkoBfxfo4cd5xUheEk9L7FeXDh/g
r82BiPEePikE43pk2PeOeGVUEhzm3jRz3gZP7rnnZSZwAUQJqeC6VgU8uUK+Dv2cr4e6LSmQyNrX
NzzncokoAKdhE4lUgpk+ZCDP+DYc56Yan3nLsSY1GqGRo6DWjDYTMKQqAlyIAX5SGFN1HtUwSoRb
s0fFu6WWzLZ0NjVb9ApkSrotJ+NZsG+ru7YwT5gtggN/c7CLhCKCJic68+0uMLnWZIGJ/OXofTJf
lXTU3Q4mJblDtHLEOaUkcuTXqvf52WTteI8qZfZAGISZPZ002zfxnt2vu44KcVPjSLpNDnJHeofk
AohkKvQAr79vHekNwqIw+cTwqpYMfqrM/RHmGzE+wH3uuVvKoILkCuLZY8ko/yQ04pqMZCADePPn
1cBMlkNdOrWL8N5mhgF5Rc57vFopxqxS6B+ZFfW47/OV9msFbos4lWZhC/O3hQkT77clPKB2kgff
5SzO5Xci2Y79w5QByekZvePyiM6VlNOybMccxDKCcD+e98YYPehfqDIh4Ajc5cznHcz/EMwUEwpx
6bjCGPe6a4dpQVQ4sz/iPdlWPkPsz7BQxfjpSwvsbwgWnw6Hw9s1Udm/JiRRM8QLEn/IjvCNmJT+
HgcrcrYzn725Dg3PXWfYJvWzijbGEz+MzmJcqk9DjFvC9w3SYe9bHXdG6DN+dEfcgd6DVp4Lp4U3
8hdGwUs4q6Ez1aFXXyKmwgLpMYlzJ0JDXbi5ymcFPckFYAKWm5hpoQxaKLqfpA9Zgj8Z0jJlg+nZ
DUP1j8okqYYuy+7htHLGmNPKbVB5PnpJ8v0QMgsEaGlIkLcZldrA1I1vqfB4GtLnfEal2ZxVJOdT
MgtrEytRxuVAMkPH5SYe+vlHDjJxF63ratb60DzN5K2zt6MzckCGACkEM0tOhOh1huxSSxBSoABg
p3tJBpk254J8Q3s5ZCvEp2nHWA2EtowUF19RtpVEMCTOYWICS/pc5nwIQF/R33Dj9YI5xwX9WydK
5VnSvBPRzn2CXcn8aaQoTbwqHfXCaMsNDE8+7su6q5gAB1bzfNplwqm7WluzpGCcjasQwlhgiwzY
zBnPnPNe/WxiphKejktsdagj69uLRlTO3TVceu4hPof8+7svnCUXP9XC2wTVreTs6eeb1ibuJmaA
exJiP8+/4VXqGjvLleAywm5kO8KNi1hQxyTuPfuWy5IuimfBqS43XO4FccELejWVsWYZDf5jGa9R
bpuiCKCE8+D6Ga/jVlo4gsB4YKBLBJTiCvzZxiVGs0VkEcFDHbZk2aSYZ1sdOcpABiyhhSyO4RpH
yfDuJ9JTBiQ/cGrzO2jBQ+7CrYIPAszo8cD/GLzDabsgIHtGu7lwRl0Lmpgw+44le6owUKkyJQaF
C+zvLwDbGCPwH2ShZGJMRYqwv3TPY+HLUh/R0p0WfV288lZuwab/oUjhlsBcNH94hpTRya2zngyg
UoJeieyaNzy+l2hqjejWjbH812nE6T+j18ckqNKv+CQEmdHCHDajSwq/39TaTz9JUd9Z1Mycvh93
Z5OHIB8QXKCsqXimFbH/O1CI0LNMHK29zZFhQ8eANkb8l/gHzNjcFW5t5sXBZogi2KXDRSif4otg
xWz/oioSZiabyERedqwQirlYWH3SMbJ5h8zpewBg52I/RtgzOA9otJzyqOHhXmCW3QrHyCMMGaZx
5Kw+b5Qshb+hy5/9On+MJGHJuibJ5b/whPJdkIdr5Qa58ifb5gEjuRBFdFYbbJbrIqrnFQkOWRlU
0VWvTb8u3rg4GHDBIx0FwU4OGL8O7aSD3rqnyayx0sH2r83m/EhVeRw/RYqxTZ3yMibbw0NCkiDq
VJm0z0b4YSMi2IIh+jpCxQVCOjDr8s/6ZOttVcO+mKfHlB/X+nCLwFVDS6EvbYhn8vyxJPWMVqeq
4EHyTMhtFhDMyaBDDK78w1+8LBK7RadWq19mclRMCE2qB04jwX8linHzlvjrM5Uw4B4bfGlXI0hi
6yrQD9B8C2sQKGz0BK5/H1Ira2u/7u3AZ4+TaTMK0c+QMMrM/8WyKqtJtOCHnA2Dk5EuMJXS0xfb
GILe198R3NG4l5CuzqEIW7L28gwfoZnvsxj3/NcR/u1k0VkUdwdV3PNi5l0p5J+LLgfVM2VKNIVA
1h+JVa3gRuTryl4zDyOxgnMoYI+YtTc8z/ZVpD6jsTAiSJnQCmkO995G0qFrcVePdgNjp8iNay/t
v+vUkOO7ySWbCNc8KwEGi45XUtQQv+PU3duQy6s3IcIcmEzF7HiJWMx23sDrQ0XFvgdMlqLzwSJa
wGoeTbuioGej5xiCK+SHbbkxXPkQeVkr7V7uDuIEtKR0XeNH2EMnXBSj4fPT0iY7jgXXsuTXYXWk
jUXhxpGRIVsEiuf3FV15mOc0P+kOX3Lezq2Xhfs3qPpdRBtPGznstDVcSeci8S8RoB2t1X2IUigh
7sBCTR73YW+yba+L149jV4FI3FxdPzF6aJsPjPCy+7jFMH4v631qagjMxcBkTZUXyJiBInQVzfZN
E09+Nx+XwQi1nEkcYBD+ZHy1m8k2pcrnI38X6UlcB3MDg/tGPe8Vrr3yvoIjvwJ1OWjkDTatlh/a
lgZ84KfWJaX2KQhDSgff1RdcLZihp/j41c5kOgZ95ZfghDBgxFDenypNImUlShSnfWv3KgGLzo9q
SSrZB4ImgCoBnalQjaaJ/JobhfCZ6NC2YOUaojPOtofVno6ZYXui4uKzs60/WqLgAOHy6lKsPXhK
1BBR5gNrAYkkjXWqhn0zL0Lj9MafpEupr4lMNczhyOrxhMtRWQJo7cJXmYQQ4yb39GWUzs1jXRpY
bGpuOJPIR8ckvqiz20t4UmUB7JYd2mRD1Of+I78KT4WIyTmohNl1diGFim7ZEYeyiJpFepbDgoua
hELxewOilBiK12SQVLZRO9Dyx0+xWN3Cm6uVqLmNiMCyZv01smE17gFDr9G9FTtmnDj5vcLr8mog
+B1n4y/b8frxK/fNV4ScKdStVg2laE6+DfeXIuSjd5mFJapprmGdJvRQLZodxjJrD21hWQS0h8Dx
BNoXdlFNiaP5YCxJnlTSSKLkuk15h2hX6M/wmzpfZ9ys8FIxnVcQd93e2auZ62S45PgBaKJaEgMu
bU65qXwezqeUtSCGavfdTOEGo/aOu2p9/1h/MVvPuwz30KsR+v24lQwdO7U48Nf4OQeAEc7SMVPH
a2wRUlweJe5H8J3Nrojhxe2GL4qH+yWFUiGJJgOmnhiGnSbcNAl87HCWoZM/hrpBMxyfjO4bKQDh
zui9Dap9gS2x+2+pAwbTTWapy1yHtATlKON1CkGRTFJRN9ZNfKSsKerJJYvLW8K4T7G3Be91bNn8
E6ON8i36KovnurgE6n1uwHILKYYwryldntJg2qpMfzJvStjolbEVEJQ15LeTsk87ZhyYdkSTI0jd
z3rhmQFiYne04K7/MnFEco/VGjmTjzTBABjh79tWUO6srEnVuvZnMRJswCfdGcJcGSHiy1S/ad51
WXw3TLu8Wh60h0wVSeK1/KQyaibydJZNs1QkJ78DqbvcAeHEY6Zlh/95AhcXeod3xlCO0efMhSGy
4MALpZaA70PIyG4MInlCYXH3oUOAUzrWllIck37gubODKVZKorwHTqPUxCAPclkIYz8KoXS90zbk
gtc6Eb72Db4EjoqHaHfDqRYLhIlHl+gg75/NC80Jn6dvgzcarua1zvc/IzStwfC1crQTOrZu79S+
4zdiH37qZgWnFLvK1uto+24rxrcCqW4tutO/ppLQKjKpPYptx+lxrzZomIeMLUAu7mPga+ukny6d
phhWCydLzTacidcJC1E2t0yZzIQZTtJf/r/n0HS2wcrXfxEQ2mlu6tny7HgCDob39e+kA+hnruom
sb/4wmKMn8Ht2H2pHUJwcejKs6wKcDN2ZrxrS6m/fkIuWHSiOGFhBMT6dHuZ4iD/hAcWLpbHw6R+
JTqLqMQQuV+o4rxZj1XNzarmUXwAqvvsswFo4KOMnvgMpKvpYjmtwliamDFTUsFAqMzd0KkKFuwI
oE57ImLFgkVNCALIakZM+Fcks3NbWlYIjQHe4sfCeaENE2BTB9MOFSx1b88ojinkIGX0duNCcqL1
EX7u0cUFNXJeuJ1qi9z8bHfCtaXIa/gx+LhIREj5OxtnnoqSimstnI+AcAoBxByuhICam0l1XsXT
nvQAYd05/d/85rX1AV3Ed1hL7enRp1s9+HvdSJig1sfc4/IbzOJJqT/ThVJ1m0GBbuWioPnlKl/r
T9CxQ5BnAY1lYEvZAfyJogDxddbSZ72BgIW9vybplNGJFwpJVQPmFVgTqzn3QiWEsqgAipLsZZ3S
wjZZy05Y8zOLud8sH0C5HvtOOOsubzlGAB17AEAh5yZfok6PAUl7G89BXPPV5ASkAcoefvKuTUwb
+jBgaRxHyu3E/UNyOmHyHHa2sn0adVmFjCjAjycrzyNn2R8AOWI5bgTOU5ABqeM0xbpxOAbKBReW
yew0jfegpZ9MbGGHFHxdvZIAFwDH9jdUoh35jv6uyRX3JAAQbjfEmjdtwlmvVfDIIcHM/wsFe3MR
WYz44389wd65kdAgFKqj+JWIrBCSv/QlYtTCYlwdABPLr8dIo8VSNWuNaNYo7VEXjX6dUJk5m+yz
5LGRbdnZ18HMKB132RS0CDreu5ImrVy/KpV0rxHJ41sC9k9/HDleSCgBApvInjcCJ513OWa7QeUR
aMDHWUPL+L5XoQJgu1xP8GGjXD5pxybVfOCaMsCUI8fZBAPWj5+6h7oXDoLF6DF/S6cFypJLRrZk
5A58WlyyapQWiQh+xh506h6ehChRvcFw7EznHSmga6nYDzdG5171P0EJlJcTUkdFj5V8ZNbjV34F
AChlFunhp/5JpHT+ZLNJTyrreKM4WnajQH5lu1km54sNPXTLLmm2IFtxcf9WbsEK2s8J5x8QcgXM
RrL+cjln66dIBHbWtd/SUtAttbOHFP9hp5KYE54oyBkcj2hNXKvnpnlr2CHzwVXmOTFv88f4yijV
ublvHHXW/LD9td+LVBo85WzVxV3LJOGmMhQPXzB0UPwrCeJ0JE+RMJyoQmFhidaXG7dDYyD5tlZ+
hk+PgFFFHwF1qNBTh7jWdyb41VYdJhpIGgj4VoemHZOQgDDE2CyJLKeW3Ksrltiw0sqZYstlUTF0
Es9O1aCul9B3fBzRvYVc/UpcIzLJYcxSXx2Mc0MzIO6AOst7GWa6cT3J4c/NVxRAm5czjdx/FiVo
LuE99W+MGehRrRSMcQDqOIj/KVUFoiTsu8j8O0JSTWgg/AjPQGqglMLFSdeS/3flZARxh9YEvsKx
gmbxBUpP7idEwb/+AxMIvGO5+GHIDmMQApnPIrREEGPNseobfQx1pF6unYqBIqu+3jpL7lSQ+rWS
S1vE7tcTCVOL6U5D3rQoHPOsL6+rSBrGmlE6SnTeWMW53e5xJ8RApBmK+GDKG2a4jBq1H6oPcrYg
6MHK3jbovzjFcd1OYLcNK1Vf81YqyyzFvsN4f8O6Dnoa0sKkLgMKOa2gVIRdN+Vbfidl6ipRdpTK
EQPNpKfBPmIqdOrBOjBYi5Rh7gVJjQRChMcH/cnyzz+USzPobFybAEwvK96byzk8DmY0oMEhxxct
7QOFScUlE8iuH6sqFhamcuj7poShIAmATzzc1I15HsRSTBtlBp1maUkg5aOCctgAeyBVAMwsQA6c
h1hNMB+5xO5/IjK4gB6NYIb/xzRQvO/rNswtr6mPBQSZ/HRBYvWjXiyNslOuEHDQeXx0tDkTVe2J
9q0KSlTozh0S2zEp9sekXKaOffYkgZ3ZJ9zHXQaANwaB+AmjRt2KbV1k8MyRIeUhMQDnA/fjN/Uf
j+DpDoWxdWTpYED8VAOBAIyo1f2ZoUgxwQ9Oi1LPIYoGvvAxADeke5PjQTK24iDwfzL6Z18Tip70
fmPszVJeDb3D4MfGTbgm/35/ILfB3njhSb1KIG6GPdj4uDSBGaasgjVU56TL6t2/1oNBy00t4417
Wg/DA7dmP5yq/tjjP4HFD7WxiK4a4bvuK1WoWlMyDIA7l0BFQqfMuvtcYHIKdU4HJcYCybfKoHFM
sDagACvAEj60CcR5Y4Qp2ExxontXBGePSGBnQ8XnUHh87mXn/m9SCiVzY9/PbjyfsaQAXU1V4O73
0x+swKr02z/L/KL65lQWU7eijSQONqRmpOc6Ztiek89eqm8IbmV8sU1m/ub3/C//k0OKvIsbwHGt
UiLwFGazSnrxD6XQSfLQfUk2+SkadxIyLvjUGY1YSkdniJYTa1pDuIB9+H8W49P8Vn1UJ2ob4xHr
eZ6nUHoK0P4mNA52cST1JhQVAB9xbOahH80gJKeh2PYKRc7csT88GQ2cc2IKfq4BudXziIta+b2X
18oUIqohKNEojQ4PccK7P9fazBcdVYrVno2uySB0uT96H8DVTuRoF4PFyUAw039kGk4tNTaYhse9
zhHfXhwwvOa5HBZxwIk//T8v7BuxScoOei8KmH0LgOxd9rNf9MwgQO/+Eja41mbQZpjoSRWe3JqU
zos0hI5IWTeaj2x3xZgY/427YAt7ewZFf+0eRBm/uMOvjyAJpXbNs7XDGHmiGe4nZmAbZec6VoWG
ugFV/kXoDUrE6pmFPokNLKEuzJcnMo5X4EBHGsvab/5dRw9aXPAcfJj99aTNdK5uPwCz24h40HsR
qnp2jdELZ/fBXuHURSPIhxSWV7N8dsxiJSr/cNEkZKu9g4xrMITarbGUkzuUHgJECU4hD0ZEHD38
SecMqdgkZGO2HSzuNyAgOjibutNzZXJVWU0B94PBH7yvhs4oI5mLUOlhWZyymOtKE3fkrRWCcRAf
l+OQmw9BSVwqRUS+B1PnqJaIrHZHgb4OLKXryd71G/o/phEn6GU4xceJz/ZWsuyPL1uPppGy8653
XjWfd2Vg8E1CoO6tmGDKJIUyiIJNsjH2sUnndc+EN2bLncj0hZb/4hgLnuXY5MxjK6e3UQWwjTEV
2OiA4Kce1+gdk47cRhp9Y5lrSS+FBxaAPnBwft5VbxO33lQul5kSNsPgG1maMBypQJReuvSXVD9G
tZRXYWJSyqQd8XLOVSJMvSHpcLELZ0po23AHfhqAAdRKlLfp8oZbQc+Ith4e5gxt0PTht4LlYmhM
8BiHsgA8qprwM6lgWKerpNmA9kOgXFouzDEbrvhJhIEywjC0pwmedxKXutA4lFx69hT6yKgD4MbG
hQH0Qw1Mnw/l1BUyku89c2QtoJWJlkzqFU5UgSz9i56V06VpVMrDjbR76zQZhn9aMBX4V4UwwgnO
m2zE0U1jDFIsaCHz1BZlMWUkXGcWxlAk9t6Ilg8+RhZZMnJyYShLjSnvCnTZCvoDpnZA8QhnX5U0
T8oEOuSzX/8wCd9QxZIiDuwb9JC01OVD2W1RhqjFkSdMj4ogdGbI1N1v1ze0c2oUVH/1GoNBI4pG
VZolQtfToyPx2CHXy4t7lrs43OqskI9MbHK65zok7YDr+HereOpaU+F9rfwjSPIYnWev832E68Jg
RxfvcqCGP7bDKntc5pbrGOa/3iWxeSSAQXldUzZak1IgT99L2HpcZYARwwa5iL9Kil0r4Ht5dOFp
93jAE9q0u6GEEVMOUA5uAiab4c/+Cx9TZ8WqG1qfxJWz/gdZ9pvvgY4RITadXkNZs+neVtcT7DIM
YPJt04m4Rjw/zDsBmmYua6uQryJ+TZtNyOf6J/rIn3NPM5grsDmCW5sKRgC7Us30GS8jj1UgxgZ/
5mv5vQVZYDFSCpOzwj7hvmbpzvhC6ude3y4tFc7GX+Dg4cr04DOZHNSb6PULBpx/atQsV6eIwdC1
Kq1eiFgncTk1pxqRvOBmjhZZf969QnRSK0Ucsq+VUBkTKhjzcrMUpaUzFaRF/0bm/mmu/WG2ym1y
m8i5CbhGNeGDSyBDz70NcPlA0GOl3YnM5lM1fIgBf2YJLQbbfWtdo91JpXGA+K/CdPFj4Piie00S
rk8BNePCGgQlE/nQSwdh2y/jjUfVDHCr3ksspVlWMm0KCgSaldMMghOs/WWI9mreE8K9MWQqZuoE
uxWFnAMplZpXOHSYIQxe/J8BgpxQozyjM1AaVaYxWTObXTV2WYSQFFbPloJlhI2B4+HXnS2Zuvv8
pXfjOjn5mtmykXPEF+8rez+byJZMHU7BvZrZSsw+Y9M++ob+KIHpY0YrtM/yLQdLF+4gWIJtRcBv
3Ort59nel1gTBZfPDg8Wf6EFfYeIEGQjbWkalL57o4aIS3oBzW7O/CnzrWX4YRnYchN2cMjCq6Hu
JSolAnTUk803zSvSdbcihPqdMu7ENB0jZhzMuveS5qJNkAGCvsC1+QmaUi0UC/ocKF5snxWh7EEj
7FpYYd5zCwF3ebGt0c0smZb3Sf74NBNOV1HG0NW6NxDGHYKWyx5+dKBKPSooACtrVQ/L54chrqFI
7r1q9NS02xU6xmcCb+tuVCHUM0isJr5KhKj42rZ/ozpRKyBP9p5hmbNb6g44DKucGQ4BdwId7y7l
ngAKc2tD7pWZE+5Agh6qsMIEl/TrjfSx/gBpShhCUD8PbPzUqFVgk87uGGzPaDQm8q0SpbYLUj87
SWzwHye/IGSJJyfh9II/dEALz+LiGeQy79q0y+CM9UQ+d9EvCXJdmRIyY0ru6nxelhAqbUnDMEEY
YEcBCJLpk8tUn45ahMy8gQeMCFudsy9c9kbxi4yG3w9v49eBP9rjO5lCr3nHNWI1/EvVS2Z/pcXo
Mwaw6wljQrbUc5l8UJEkTHg3Ur15JIXqhbsQaiV2JNVZNHczFTgcNWfU/VxWlXyJKtpQUXnJ69Zi
kLwpdXyEN4XbWOpopvEIxvwkGC0yl/N1aGfPmcrbE3hqU3KXhgNFiiSVU0oXLfWindoJJWx4KHqc
O0wcnAIfTL6/kNpLifPJ0Knlrv8w8xnD5pa0M6isH2PqyHaS79U7vFdoZfvsazg7CuWh4r/dc4/t
uiAdlbeFCcP2B2O2CyCatHOFV5mUjxudHJUfcRtgEBJuSJTczU4btDxKZYCFOTMZF92lSEnB3n13
JHzXQQQoHTCuYKroQbnq3Yi5yXMt9d/gkOh4CCP8g27POjOarVmffDNSLeQixLuEwYPjOdUPrvu8
ReYPD4Wng5lXrdMcCtMkjGPuSO1DmzyMqJoYUhMXYQNytOIn/VGrU22TUDW9f8K0Pi59SwXJQX70
uid4QI2Ryb4i/jp1WN2d73aV3Km4ZX6M2/30gwL3ctMSjDLTpRwiq1RfGNS5HO2kjuMi2PAM0FsA
t5Si0zudXMPVBSPi5xC9wciPA2tfYLmMZQmrQkndp5cDMk7oG8M4O8TOiGV8kP+xu3mhmMhPu+yn
F0ibKuAtO0xwOtA6w9DJMyjUb1bJVi5NVHY87w6RszKne4okvJSacIKTYcIzVcE+XidUqsD8ieUb
V/4W38eF2+Fd9lzeJWX+2XDp49JT47hST5ZAcC+ddCKwkV/qg3xXuWxwh++cP9RQx/eURdqxzYk5
g030Lb9qnUPNJl5pMaXLdmKGp1oYMtxb6OJzEJtjTxuSm/YJuQJldYXMmyrmOk4JKfyPMip5uAev
JjuQFUp2fCaqT3e/26Z55efG5V5QDIRWjIrdOWFTOr4pJL3TZACQuMls5k2tC2Dxl03Usa7lCEj3
gcSGPL9ObE6Nb/EfV9Ui6EjbTM5zsI08I8aN2J0EjQQpkRHVsUEsUhggUfjo3Y2i9HAQPWThiilC
4Lno4GBNrUA2CQh2jBq7v6LOiyfwpiflOjtIa9gQ11SWLElJZAjY2nlZlCfR5RI6HpfH3tMwyKHI
XM+mhbBveENy+0gtb71tJLb9TiTxiIbwrd+NmR+1i5d2k3GUHl/k1scUy/gOdzcfcqmO6d4fcLhy
ZooEt7HtANC6gPo3tN3MenckxjNQgBu1Ee+OT6jLiG0INHgWMfHiI11IzHbr1MkrT20OmYF1OHKv
d51k9YagPAD+yZ2QAlG++67CVejoVLu5SMYX3kiEXprQ+QG0EcXTchdJXCPttYOTwDcoF0xbX0LP
HkFZas9bthGesHIP/28K57A6d1WxJufDZv0Mfw8b6DLssysUYQoxcX6QAKUIrRSfGzjzVDv2aBPv
6aGYtHi6H/1rF8r+i0YbWNEIXyRg9A3JYJNYpD+jMMnIfGVaIpv4f/vITdzeb5TFp4bpuxKsOvx5
GEMe6LzdsfHZfE83hQS7WkLkzB6haOiBcu3W7TEyRq4CR0a5QbxqeT0XBPc2TVuJ+jeO/DFasJoM
yMAUdG9uAyGBJvrXIFH3fm73+zzuF3+Zf7ZOnkyJ+BTilKul+rURvYvwcgIIklH/ym/AzXlkucZD
ZN5joz3Jw54FNC+z30N/mNm7l9JyS3lyFkz5oiZQ87kuRS/gWTgRouMvRtOoX1mFQs4//mxwnE36
6NkqnN3+jHxcp6DSukIWlEUgh9j7klFMhP1iatF3tkV1ecl1LIG28rxCWVh0YI0Gy4ivWHcuebMq
FSr+UWn2hJbCWLqClYmMAebP3z3lRR85JFq1FlYosG4tVBPXcf7/6aJrgXQP2xfeYPHBgoCq8+dH
a9YpYMq4qOWtR6RjIm7F4qG9uXIUtbq/3R+84bKTJCbDESyJ1pI04/YllfaNeVsi96t5wLLunn8U
KK7yrclnVfgtpC2cKqGjrR3k0o7RQrZwY52PB3c48ZrPMWNB6e5xOZ/dyxHlXr/QcUGGcS4C0wnr
S9pZmbozifHMWTMKtZuDbEkWFPfmJo4jSgjUW7fy4jtMp4sVMCr4oGHGUOphq1HZlX2ebZwZKVmO
Ns0+Jqt8l34524GxbF7XM3MPfpCrPWCb6wOAF2zs6AfSiYI5fH1e7hkXygKVTrXw5YbGxes///bS
2XXZqDx2V077mxVcbUYWcDgPfmbMchzDdsC2RWWzw9DBWiZ8SND+oFN5WJR4yp6OIP/NtoOGuFTV
ey1T28+FEgX5cN8L+U6PvXjWp0QrziY/OUZzXOm4cIk/ZxxExINMLh6IbkFufw7sMoYSecxv44Al
OpVPknv6ix029Zo61AYa54WIR0uHKn8CUdAKpwkmKGFXhTgXxpZx1RUtFPvP33ovKDdWFGtkEDa3
QajQMdKMLlVLnla42PcEJt6JwCaa0XxMmlBO51RJW36mxGU+/eWAI2tQOFcm2yAvmbVIg2lOyaAs
bakBAea2Hjs7x7NvoKcdLhqLnAXe3t0UV/gqu0J2T63zvDTQBtFVhKrWl/57HLIgP723eR9nJQAN
JKi/oaGpWWpAALyKy4cFIOMFMouvvI1kh8KCo6WMsUsAVrmJaZUSY7lqXOo+fzQI+jW+6H4DwAXj
FQJWNNEqEYzGfSC5xQrK4OggyEOyU9v1rdTgF2vv0kvRSUA8Ix9EI8aVh1YDMOKjGOnS+OO5CaoW
AtNZZldEhqAvd57NIa3Xulwtajly7R3Ai914fwYhljgebkPfwLhdXs87l5AeFy0dF0QsHm5hmvq8
ny6wRuNbfrm5inFH3SIaQMvFRjUfs3Jg+KK1zy8xXQrlVYAvsmeqvOhg8fxRWFHXEtks3YgekUFf
UX1sxcnMQDCBWfi6oprApE8NRegGgU2tDERMb6DUgly/BIW6sJz/stu+salAc9XArA8z/8V8ZXH9
Ssy8SbZTfeppMwwj0WZPPmlGk7UF3Z/bSsZh+FF/8zgD6xFheAfH7K9ZJ3QvOWE60HJ60TKcATg9
h/8I6xIJZrCA2d3VfV4GfOJV8wTBVpXPUD8CRNUZHZ+yvOxnKqGzu0P1L4/st3PvUro+/CTO5ilo
KS60mgGqbh36Fdmeg9AOuWkNPnzPm2JmloDyPQe9cz1zlbGya5Sg1lFnvVbuoU2O5UPlfsP9iBgu
ZvgwTowLpz5rSYrmqCzArawckHY92cSb1Tm+++wCqmxsYq9XZOUp71abIyu17PWpu49vSDi3zvu8
Bhhwt+QBz4xtyjkN4NQcxIqeyMpL3tHAZhTjwTvpsj3+Mnn557b5eJ4efS/vZc0cTL4mJQMLjJR5
oLNBByXDOy0aKZ1g9IPUn1lo6NWkVwncmY84TNrJ3Ks7M358Lv58oqTGPBJIZp0sWKWo9OvA7gb8
6BeLaGbCEuLwuX8BBw3N/fW3ezd0zKWnJI33f9qPKkEMbmHn5yd8rlul2T963F/TMC4yItyyXCzV
C28+6B53zXMEQcnMwBUKYKFXm1nbjD3CDsTlAM9Qgka5MFua+qVPSZgCHSLO9NSVySWtaAv2L+xC
N64yMi/SvlQzmoheo9w3GWxtJPOaL9Dyv4Lv0kKFjAlvoLzSFHPhAdBFgXHwhPnQy/4p+fjcaTHr
Z+HKPxPoW/YHkrsxYzzpZdv+AGKkgMMrjnnrAOTp37TptxN/14oFmeMWKGnqVQoBqjbw9ArhA3K0
gBef4tbCFnJYjI+MFm6aQEXUy1fT95krwL2jKmq7rYB+EnT7oc4AXI6ZQYXhiDtRk453emHYlXFA
kH4x8bV9xnDx6ePHofspZChKm98F9nOvEPR+KHRMwXMFOvA8R2ftzHZOXlEjUtbQN8CsHzTCI42w
bySd+v6y9lD/OpxC0iU3DzpCShwqqsWg8CYP/iY7G+CvbpOst1vYiZQkospIMeMV31pNHba+5ISp
WMQPA9HpyL8kZCjR8TEwzexTyAhYVT2FSySIleSgNohrodlA+wtAWEUM7Avt6bsbMjkyA+eHcfoW
G+97pGqgyGUOptiZnHL06tPIRPfqyZfYbl2+tCG1yYQpD/A8OTU3PeFioubvKWsN70Ed1IvPvLgd
c1v/XvvkhboIvkpAinkGTfKtNgIyT1OXryZSSQ03caxkZ+ekMYrAyqxT/+BbDMuP5YifoXiZ1x4J
7e0VXev7NwD5xIo02b+bzthAbRHqVu63rehVqtgdmpQbenqJ9KhGTvJTJWSXeXnsAcStsF9lIjh/
Eurd7dPERkEerd+lranCM1WuIYgYWszf6kc7V5493SyulqbBy/ds8G/b0+yw4PzvO2aatmXIEZSy
v6a22Vs8hYYHbXG2gSDjyrErQTBe+hO1oLt9GK/RYm471FBQOs/dWK7OvwgQ9z3gT0tIsYo/f4BD
JVmEH8DMOcWK+86ZAlqdN+iOyacYKnvGQIWkAAiciBjzMkClfUulA5KhaDQDXklCxgtYeW0HxGeB
/pVBOivOHwUU+rPYCNXXOPbMXLZ3KbY4MsufXpZyPoPLhZz61oCIebY7O9ZjqDdKXOP5prwyIYWb
cNpWZdlWSmUDJ87w27VgFdpPIyjd/o3WaTjxVn5U3bXQ1fi5gWxZ2s1xpm39QPc2DVP4RU/EtEnE
VTExSUwq5ldnp93UtvCNmpy40GmcDeRTefhZQn6VBfXJJL1JKvnIOTnsF7Gx2sKOYhOeBTZ5U/WV
YWopMD+3ZXQsnPQd7y1YwzxWJHMY/kt31lFalnESdXzBukqV0Uxg4Yg+XfNiJ9UYhK09SX4e9h9x
6jUXbAlxgUdzzqq72d6f8rL0QeFO9y2cCSw8t+wsgjT4HLQzqA1LUJ7oYnMJl4HUoxGcwZNUPHRl
90/j9CzI9ZKt61nt1wVytxrigggMWucFnGAda1nW5YAhuZrBn2KwGpkErdqA5mgMO1xXlE2RIQVQ
Wi6AYAlPIWMOPD1bHQcp2xEKmbuTI+zWJE0JFqFBTzK+ktPC7rcIl+jf0Slo7HYHAc5Of3fSUMsi
vVhGwLex6i5YBxBCATJGkS7MPHC4Zi2RQjpqjwVOwATBS1Q/WdQJjUR8Nw+NQLA1oarEugn3q42i
FYULCq3BriCt9Cw6RjXgG/WG0yBjWlf9+sz5ksW52PwSydUSmMFsjB/QeEPsvNI7H0ySMdDWSA84
iZYM49fjjZjWfTyqZb5Mzt5KLzL4FMBB+7fSN/dcEo9LKxyHIGU+4j8oEuMWHbxAg3+sQt7RnqTt
64ovcU9pL1pfsoDqkQL7y/L1P8vV7yjnxdUnXCE62+WikqF6RRjDgVB6aNMU4FWY3bN//lXE/X1L
AIzfR9IH/TpOYuJI6gH9Gd8gdXlXmmDjAh9NX3t2cPGMq93cA2Ni7CUoXc2dSTTzHEX5miRV0mF7
A03SS9goE+DTyOzEtRsB5gGtc5XOPixoz7eBCpwzr9PEK3T1SH7qZ71kiiy4cDICOV/XqILXBSrZ
E5QJ9ZyRkQ2JzqP3IS109GhslHdt0m7WfhN+8p6ZvFUFHcLqt2+HsFJqEYGRrpcnAWvsiTE6pMpa
FmmfBtfIsWrkHxvLClO7/ffYLvpLjIqCefKT6esIsPeNXIDBzh5+Ad03F/+mjge8NRwJzi3iUEVC
l390bwQ9YnRxDJDylv/d26UBmjlznlo4CoWgkKY+U7PgXi+qTjgWGVGxc3lrzlDBVSntw6aIS1IE
YNhPXQ3s9qJbznRV6KptRC3xeDjFxmP0jIzSfpF/i90f+gywukVAim8u7s87rwDyJ8Aj2rw3QtuG
HVCGLuSomf56KUI9nNloMajVGYHaAfwDF/5do4lgSl3t6ju/C0IwuNGSuTtADdG89z9CbFsHqJXP
7gnVahGUfrpUi/HsPuvwSBgK8NapN6HL36kEFzqMEF8epEelVoMmYqE7tEhc3G3Jf94e3wvYdKBa
VTyiutN6ODF3bofKy9PYec3serUSNoA59F+eEt01+l8hyTKiCNklYOi/8ejpV7Xy0rJW7i/Vuf1k
azylYCeW2IEUiB4rTvaUGKo4VCbs1bevELGZ6sYywKbNruRv56Gy8ij8Xtfb9sXz9RtEf+rCPoUQ
/82aKrZxxjUdmCgXOh9Ib3jq4LmnmNchgcHeMJQoRuQJy8q5TdVvHxV8s5tRI+rB0ij0j6gII1k7
PpO4fCjPPPfjsBifbCrslicIr3C3CW+EuxSCP1OOWdXR8nn7Qoc5gz9zNvzHw6b+p1/WD0wxAbvC
I3OnQj/egMi7rq5d4A4a2H24IZNPo8UFCVf6XIcdRQaSluKb1jtTo8oPX+HoTbw4YOSI1/3hJuUP
WA/BuehYfeP374HhoFJorEvRqjaDB40MMGcoaRfYF94rXUepqkv6yqYQqcgh2OaJReaHc4xYw7+C
mYWsaotrGJsqDcVvgHVhxnLQAnRd5rZLfliLr5bUpWUgYSjGtiEO4WlFOVp4nij81KCn9RFISjIm
Y6/sW7lVEfL5hjd3PQk7XJwn5Hm3I1yrbiMq/Q4xv1a71oqSZhwdCaaNKjJd7Sj+VxZwG3PBZwiH
b4WbMZ6rXZi0jGkWQXglP7/tuUERKsanhFH2Gt2OKJyPMdU52RxsO6FNYXf3VOG+hefW/BWemnX9
gZJ5ZuzvNQEpCMO65cn2+AaeN/1dPcglu1McER1Piy44v4tnRI6dtxbWdcDEntHcX1s2w1QcyuPJ
bgKD9IF+o6pKDyu1XsWMAfVY9clX3EbfMGBrVLwTsD/+iPGzAdOXqPQ41GM7wyXhg9TSC9lwWcnH
SoHQ7aptLr7R2bkaM/ofYsWlrVVH/4PH+LJig3vSPWFm951hii+teW9DfZey58bFgajvzVT8ur7x
auuQRmBm8KQn8Hw21LJNxwyVWpPr8bUAmX/cvR6xH0iMz7A6PMC/1IKhKzbIsUJNwrh7UMdvALe7
f9TqAxBQRgHWPw11y1rx6mS88xuathmK9zgf8QsxmK60aCPDpac3Qjt6ca5bFe6zbSINXtDiQRW7
0IY/E733uX0ZN59AFhgnjYThbS4wIYLD/Wtb7m63uTHo+erEz/Wdk4ekJ0LfAMCZFUHKJi3Ua+/n
iRPGvJQdfE9ao+u+1cru408xmnQwPpqZDLsZWi5Ow2wYiUFBCSA8fk5haMV2JTECj/GIVVtmPxTI
dcadS6mVa44xbpOfLvwynUHhrtTvtNkvygP2kF0bo6MffBFpDPLqulc0164Pn8H2q+Ea757t3pAe
HoeSUtHQCnbhwVJPsuQB1QUlMcrWi9T5FIFrw6e0NqfeFEpCrcY50cQs9gt4gsoyb4Hyt61U87Gk
OEOHfJJl4hEb6oWlm9qcEsXXYxl9wgO5yLol4l+a9SedEI15VH8asd88lWTIpEVDkxTayK/oOumA
ErtxZ57uHVoeUY3N4J5CpstFrGJQJTzg44ehO2LAooKrV15sjm+Pz5mCnREdH3jtv3EuH/WJFsSA
uCuhrdy4reUNHUnfpm4r/sRwRvmMEhkexL968qsIgMutSKykzMcjWE5X5MUlu3a6Q7TEdzYPsnQW
bR2I/K0yKeWe3rcOTVf3X7aLDliiBokqiRjSyBqPIjGa6VDYp5hd1+ky4wLlVrOyRNTkrR/2jugF
bURkgr/nJnbEQRxeck2HCnQuxiNNvIAe5oI0BDWr3ZO9SCvnqlWZLutliEKwfeBh4n+CVq83UHQ6
4b4mDcc+TkssS546CSH/5wR2cbO9Xjh1kf7BvTvUZlvdv2CCMsATWeKnu5tRuuRM4ECkK2RHV74c
x9sRs8O64bmQ3IrfwB72YAJ0wSCkam0Qisi7QW+bA+68rAl2tinRx/TYtQstfn5mJyU5/Rf+v/h0
x4qBPQomOTD1Yc+q2iBlqCioGu68wqfEyNjep/qnm8TmZpr1eW2v2qWhDwRWpzO3PZsRfWywpQ79
xL2mazWVRt9cuOCAqAQ1ncX+oiTDdG5Tbn4o2vq44TxgNPldVHa6poPQBlJIagEdSItiofywzyeG
lmyjDW0VZhR57UNW9w/Zae+JuE2O7ItoVsVFwklYJU5bmBbsQz0MdnkHR85VjWHNyk9js4UB4Xhp
GTmFk7F1/IiKhVGsHGGEBnoiLCorvB5BD/lS6prFFjiMY2Hf0Tp1wHvJnXe5s5JQrvo0gIN6MyMU
n6UCQm2n/ZiCSm3qES0iIl1qzldBf77MlUWlI87N+0NqYJOHWSAi720IJSzGZAL+EJLANbBAUodV
EpEHSwPJzmsy94ClVztgzFKkIOmaXKgbz/hZ2qqO1y0GfuwJp83oPGcqR8R0DOi2V2ufAMb6wnn7
wyLqUuuPNmVtrVWN1fo/k/yCjt8y7Wo/iUIpkgBp3G473OJiUAcUUQVFrjbow8+jQeI4UAliyugj
Wsn1C+kfKklExcdVLKgTNn1iUIt0bJsBBgVxUwZCQHMzDTclZu/jpNmbBdj0GdjDslgOWHD4eY6D
K/fdpyMYgjRuoMRJ/XGJhVYITrta1Lle6cfcBS7SYiD67FpflQjuTJMzPV72RBCGmYbgZOAdI9g/
Bq6+CW7eZgccfUnBc65xncIkdfSChBvK9pmaWgxTXDsXpZikqge30+SKzrWUnl00nZXzXQxIvBD0
HKqZPhh9++bEJU8VMJAVVVvFrJkt1D8SI+6r6PlWhOC/qxlv/u9U71SxSpU0hbv8fHSfkODcuxSx
/lDF9paTqVxTBz4ca5AuXVmxO20dSPV7kju1yv8UwRrGR00v61zDxSy03zVIrHxsFsbRNqtSXfG6
mQqGDZ9J3OnGF8LHtJh3r5SgOV+BsaoyipeC0J8LvkkuR1CN3kNLTO3hYLdewOnOoa14SLe+GQM7
9hFqIM8loG4e2dz9Q8/mEj7nw6XsTzpVMFXYmfQM+ye6AW/Z2nP31eNEGHxz4wxd0jPsVsTFaCUH
KvF39phGg+1Or0SN5TuwNJGVwHew7zwKxXaa50d4pp1DD2iTCf+lmkpZMPVUVLyiv3reYBAbJhja
vpGeYF/3x1OT7p6A83KGVbJeMFCAvahNYWhh54KvOUVk/4R02Y/eITo9C5rgoprqqwv3z9ZA8SOA
noxyNOq9mAVo8r6A77nLA5Y84ImnMI+c9rNbhB+3NX7DgwIuTYnm73pfoaQBfz1aTXiO4oER40Ve
dT82ps5jhhZ1+af0LOnFZx9Gnm1i8HlOO+f5QbEV1zXmBx/E+bZoQ36EewhTha5+K7e6J3dQQV4/
qQLL5AObH3w+jjhulja/bgo82A699Ry3ohR+i5615PsltbpEZQ7RtjkQJsNso6/HVAdD/NE/8V6U
Gd/ZiQ9dS9zfhnSXvYDVK8EVSx89acE7iNxv2qzrB9rmrDK+VJA32HtePXCRIMPeKEzcGM3/pd8O
RCtDfjd81tqHBaGQKXbyEbt0FlTGtmCubqNpcwiq20kD9BHQ0pHfkVYUa3SP6pp66v75dTAVj1WD
1y9hCX6tHMGbB2g4rk4SZaUT6qVbl463DA3kJEf7mdJlO6JbIGZehSRhwLrAfNpS3CnKX0yzbV5m
8AilGvt/nYAVK0Ns4Hjp3CT7rDrJ7pkKRLFiqRiHLuj+y0o3hLrO0KpNrZxUDeEw0C40f84f23T0
ZWeYmPPcoZgKfAmXHTtWg7/TsCXcWFF51QVVlpd7TYhcWV7wJGnJij6RRn3kXK8B1MeH/WZ0QAdl
KKwE+S5oLD6wZp1XCoO+08VukJG0Oww9XQnDW9tJo6wyRpvQn0NrdF10n+Zkwx6jlXNCUaGSHckY
BJyZ1fZW2emwP98ulGYmtAX+O+e8qxySm7G9Nx5Ym266PGIQUgqB0686onUbo8MEcm43V7pwOP3W
MstuZ06a6mRUYxcTvlGnUpI2tRSykp016eoIge4gLbsdSMBGavzwa8gz3gYjQnujDGuIDDyRptrc
vBjI2TP9Mo70p0bibPx89Ec+NsP58g2iWp29yIfmYiZ18IAb5eZQr0/7D0sQ7fYvYnyeTunDs9gU
KKDuxDOsDAt0BPeQJsJmoh0fryTY1FoloXNrArixk2HG6jAGCLJSjT7aXacuFTOufatd7owgL3rR
gE9I+BSndg4tGDMWRO2XPWet4K+n14dmLqJgEdC1wRKsExOLTSo6z1FFJ6aSTeZBJgLsmWPA/8Pm
ugSbuZe+U/xgevipTBjxDtUTF31aDp4m24NNG2TOQ0570E2OKc05MjtOO4w9bD7JpvxNp9GL9yI+
3unAH1fHTVfDoGF3cBfy5hsRvfpKMQ4eNiDngFhuksGXxS55SsSnp3d7MGW2W4cIbhNYonjRw4zy
Tg70w7fr3ZdOZEpaDe3DlORItzVKvmE9sQGV5PG2tFyvRsyjSe68DvVDhtheoXre6miq1O5+/J+P
swK9XsDuQw2eMgoYqiv1LMp+6DMtg6LMzTVaA8SwT+D8m92FOtbEDgIQc+kCwtxc3ZH9R35aSiDH
I0xEnYZ7vPO85QN1b08EGQxC3jdg48vpG15mjBKBlJrGjF3YOQURTvIQhJqKUb/JQAEMzD4BLpjR
1EzjMMX6t5ZI28S0tCLQBdExSUwuV3GvT9FR2UnxwfMV8555VEeek30yxRgz3o0mQgi+LU1x3QvW
8P7QcHnrh0Zdemzy+mUdetie//B99m7ilRcLPjZVhQOymDGmX+TGk7vuxZnZcYhpTE+Hv0D90rI7
g/ca4M6Om6Fj1+AJQ079HWqH5z7rEVPc7fnOl+IwR0AVaT6cw/rRGy993ayxN5fg5jUwlSOjxiYE
csLyLhqBoyiHJSj6wTlQFavvH6K05/Z3Kxv1u7aIS2EENVQVFJELxGexpPVAEQkTyDNj0R7M+33W
8nBNIQG3ZJzjnqsyck6fpdpmKoSah23Q1WG7v6iAc5Ssx1eunjc4zBdRsaOWXHoJIoYBBUAZu8VJ
Jqx+qc34pDzFYje5KfK+2j3qEv3a84L2CqQJpqAJ67eFEGGdjngJYHsvZuGXmybiw7jpahtGipwB
3g4MJ/4nO7BE7wNm7wETMsiPUTDhKMMXnDNLSbptrYBuxmxXLIxk/S10JcvY3593gyP3G1Xk/TlS
vZFK1GWnlkaBnTi38Qts3xCjZTCFsH1HxRVA/8arulgCgi2DSJf40JsxwsuWXijvluM+o6eIoVpS
D4fP6y/jDlCGJNF+pZJdK3GQ6yLm8PSNARxVm3/KDSNkAy5m9lgWE27vUruNU2SZ3pIQZwOQcKsW
qYQ1uJcpIX7i8CKPZe7r6PD433k1G3lym82Y5jlAZHbK4epVxmF+QYGCjXZYyF6EByGVwC+Nna9V
jucyzylYJfMVXE0r1cy1OnqVGiG3fJurlJsPc8gmwa0AT6L6Hq7fummaP1nxSgg0KvKkG2xgAFFt
acOfuUaaaqLq3u5m75/DvqPH+AUSWoorfSh/vqZINlEPGbCHX6GIILWrw6e0T5k+p+GFD+qO+3cm
kSXAA6G5hJCAVowuvbcxRGCn8QPzZF6lUKC+x9TjWssKA04rpC7pgeN7w6WZfXU4v+aKNQy7B9ON
/ycVE+tL+K4YuQowfJP6AWgEAY6kjROUrNFDPMxI2R4j+sOvImGkwfYNE8D1MGwiL97Qto+9cxpa
Jr0kk2390U1ZNLHxQ0eoNYejrppMvnRBcfPPiDGbiEPcrJR3LAmmDMPGJEMngIXahKBjcL8EB5o4
5WHlGhsrZ5/aLlHtAcaHvK8ITupbqx0H/Vb/4lfindwEnspkVKDdUzSmWskoqlB5PMJUVKkXrI9G
vCBcZO/YEKp7NUzAhfUhsklUdvIDrZx+LD/+q8pTuRYJRz7Efsj/pHCEzJvExgm2HjuYG/M94Tia
+Thkw4+iphBdDVyjGEyUV4gavlHF2+Y4DczDgezzO99bzCHYo1IUW0FuN5aX0AKoAtCpqmFedf66
iVGqUBPwOvoXRxim6moGMeAnUCrHDL0V8IbN+X85G2O7cXfq/4sMK0GusuEsJ66hFWEBbDzuaNIM
AoqrZ/XZXqPK6azu9bY5WcBHzp70k0MNH3djp7wIrLZsNdmdSQsoaFjHFXfBnETtL0pVAFhbvwq0
Cj3Mqk8LOBwUIRaOdAGrtAz1IYMidXsnRKYtHVr1sXK0UWgU5TH1oHEeQiVwlOCyZL4VkPU59Jx5
wM//yJWAN+MeLWDOR4RwQx4sPPSUN2fAlfOnacu0FG0haMKJULpAMKtZIIkP8tyqJfo8hWuVog94
w5TuD5BcwJYCZzBZ9tZH70NbO3iRdH6x3L4K3tBEuwTLZPdaVqbMYhQEU/wzo0aQERbOmZhGBIwf
KZhe8weDZewvY1+9VeI4Ufy226Tt464OopbWv9T+11tM+BhK7sXloebZz/uT8lnaiuRA+fGPsRRs
n9pQSNDhw86iwk/f/L4/V7Qwcwn/zsUfzWD4eDgekpKRJphZJyDIDYQHXzhnop7C+JwbPARphuwm
oUvImcBS6Hv3r9x+YUhStMIO06TrUAOcloAGPLa+64vsIZ1Ga4WHvh4KXTdrl4Hjx1z+FMcfRUV5
EFdbjiEOpHV09QNh/lWXxoYrwwCcx/5tBD7p1YkIRZt6fOGlRMQ/K6BUrvtO8M4EUt8Xl3SefyC9
M8y7gprq0sc1+sEZ50A+Pwieqxn8aUFmuAlGTbi3bEhTtiZ+DOpJchErcmeDjkZGgkRxg5YzOp4l
CKOICUxlNLCMLXRyhKRNzAbXeU/VCtb7uCC0vTVw0FqfCvhSmPHcCrqC/42YVi59FkFuKYUmdXz/
Rhot3vBImASgqsJxIymvrDqNtFhDqhIzvCgDbuP/X0jL+u+Hl57yTLTC6DuPKqN8TxD4tSps0NZg
t8O4vzY5ZftO3dRphlEQQWpOt0kE9telWgN86/mctNgBsvO+kR5RvFdAN6GmIHMkToPpHEzBXYZn
MR1mah1aEA+03v0BUMw4Lfm6Q7Bum26hcKTLdtEeozDpjMJ4PO0MBVopvcnFaB79ZNB55AMubtQN
XLfbNyvYwJ46yUqGRdbufplrIp0UDY5xCvlh2fHhgyJnLuauHiU93Rx77Fz/BqJQPbB32+OYWDy6
WUCF6uLpQSlu26hX+lAcXVHconLuOSJdIBkoHHNadLFf6xq8a7e81zSmcWL5M0VNFLE/dP1QFgzT
k7jB+lkpreF8qdLQNQlu/OrEWC3TsauGtyGOmVaa5y8xhCJp35xJgMNM3bJ6SsXq0EStmeWvV6gr
LJGIuXq0Dz1oIH06SPh2W0oC6yWihelfsA9j2nPattjYjDKOp0ogNG34W9ZjGLCHsIw5CEFj37t+
NhoBXWdMJGgOss1XFb0hwTc5vIhMwZcPRJUcNblqcWgmkt9MVlcvtCodrRSQhOSZKQfTYXed9ecz
C2Wbx31KMkwBferJOtT2CkGdQ6owMvssg66XnuUW2WhVVvEPwX+Q4OPcnTPHABNjE2KT6CH/qiYC
wYl2sUEH7WAKocyoTzOo6LHw0rzbIInfk3pwdA6lzTMKeJ1JoFArEP4QWj6CxNiR4PaOaKV+rz1n
LFTDg9QjR+08GyqxYX85BBAEGHpLnKqCjYNwpvv3cuCTW3Ds25PuRp4VW3xP++QVvyRf8Xg0yVhy
M6zFKmN9UvEU++rCZVeAOLSoijZt28AzvDs5Os/p7jgDIIaaQonuoi1pQPkWnBA9TZYATmMfmSHl
9H4a+Lzxt4cBCarygIb4BwhEPrvcn0VDvPvuwYXbl5B8by0K7sBTuHRlGmY3llzDXkOA7brbSS9p
xpdDeF7El1k2MsAZYek/p1jBSgWebyqWE1XA1ItOKsEfKpfMjVn7B5/p/yX83sy76lDiSsXTgjmo
f/GYXncy5jYID0ud1e6kXQAYQq3BOshSrztBNao76JHvQdYzMQnvGGv63/pjmGGwv+EglgrxpyzJ
jpHUYtPM5AyHoGml2OHIYVzmXd6l8ShRGQTlS1wr2QZhIiwZkWdS4+3y/l5jJ2Xi1I3yJwNFw8aO
BTY+87EXLTRab+3H3q/BEqT5BMrUxzsRQshS02JD2dQ+WexMm4a2RxmXVoTR6AP99tJHgHaPRNqS
tJ4NdQu69hBxqa9y3fwCfBHaJ9RSaY5B622W1thfsoHXmklvVCzKyLX7T5j4SmvS26UZjsuSMuVk
CYw/u8hjXwshjpxjbNZtRELgzuI13BvCaa9+U46TYkw+aH20izFQ09xZ6q/z3OCQ51BRG5PA0TBu
cLWjVlbWGifAq0nGWYtJr5DtZouBGy2m5OoeTnfvbH20erz7LiA7IgugAA+eHFvLwKeHEcKFs5Q6
6NbX3wS+DIMX8UT3GyLrYS7Nefi5yhfsLanlEQQDzXPZJTEIum514WLMr8LPVAl2FrMcNjTCmtCc
hEWCIb5nV2IItjHnNBK+w+daoppDDkh3yyEgLq+3c92qrNHfFtqnrbyua+Df8ywJFDnUyhTFzLCx
2/RwkiXi/6bmg96F9m2YxAwHI3dndIN3Au7Bdj8qwH4WBJcPca7nAIhMP2pELtirWNxVtaMZyT/k
BJd5RabrIU3CNrMbZ9pNJiNIqGQJjrnHGWZrk1319hyv05kmVXfJRxS+zpArfdQ1vd1PkxKdt2xE
mhdcNRMEqaDDnF3yZFGMSX48kSkinvl1agK3+CQL7RVg1sCL6wRB5iI/fNPbqeP4MxqN4ifLBYyx
2YL6+6+RI23ZCJ9IacPCJW7jlgOCn5TyoM3ohhhkb3J5EpTTyx/Zrpr/Y92eV1vdXgBD1g9/HHK0
IBxz+GhLBgqsNYcu8DwueLMCqBhAzgG9H+9ZhlO19pcvcPRvn6kAmuGzaCyv338dv5oYyMJIcFQC
Rplqqc0UWKY/18a91jZ3zK3xZA7ej2EfyILzMUJGvsMKzF27Zpi5ZjWQhTMzODysCtaVRURTqIX/
X0aaLrmP2OxZkP4sIMxjI6x/cCYYSwbNgJ8U53JcRft/RpOQlPFKnyco3gKY+JCFNc5SWb+aCrX9
9X7SH1xq00ZEpT3rEfPPL9kTtLQXTeZqEzlmLS99Lk9jrbPwDxOjDlinFHZh7TL26pajLpaCFilw
hwT/A++euGp4udjKEsyPiao6hFJniN2qUw4/mm1QffyIhu1yebzMprW5g/UMJY3XgTcM5mEXkMh1
yGC8i09fpl0bYcrDQYLKUISj1AHmeM7Fngh+Rlhwnn8bi48hL3ZT8vu+XOiWDoK0abi7jy4KxLj6
t1oGRb3yCl8/yrS1T1Jv0ukeonXZTNuUOXIBjLFtXo6VbZBzbRW6yi/wDvmyK+TZ0hfyjg8d9aWG
EM1xnYudifb9dXPCgIUvMZntk1DfMeV2w7Tx8L74Rexlm8J6Z2piazrhupWUfhphxt6QXtds5d0n
mK0UN6DjIluQ+Byb87d+s//BECOdIqDYcvsQjk0COuckUDPxOC2YnyypGu9rmAiiigPZNIcrcCst
2MmZz1m7HmZRvxSZrKglEUJ3UzNBBbxAwK8A4VceeX2vPy9HFRfqi2eDfkT9rOQ7b4knUIVswK1x
JWhHfpHcWV7nTrX5ToI964XKI6FaEGqX+rRPbO+jVYx5O4vHTmeaD02S01P3w8SRXK7/mIDm9Nj3
pVJkRC04OlkuaHYZ5BDTjnaZJtVRreZgsl0J/vCjFYF1IkSWtjA2Tfqvp2JUnGwzJDtQzrDUQA7P
P3xrDxqGKrI4p78cmZJrfYSChXcW9MRH3b/EvhAqmkUXzWAmpG47HJKCbTspCUVz6sUIuRXDJa0X
y5Eij946YEBlP3lA/9JvX5yOugBeGvziF7rzWoRtNCr24TRZ3kBPQpxVrKp8zUraC1iHV6G2jq+l
pKaEHhbQ0Yt1rmhhb/SDe6dBKnhzV2ehMY8YmwKf85askc/7eHy2isoNhG1qfByXEaZ7tP99vlV8
XneEak1pNu3KTTgdvfYryb/mZe4TQksuabNu4snRpPSKErSWrKU84IOSc5WEbGLObqPdwrFkeLGg
yz0/5uMMkz4IyYU1FMhWti4zUcmy+4E12PF4NtZSgVD+SOKLgbvbLGJeOlABV4nVH7Malr/RtPVP
OHREb2rSH/wvI5ldn7fawBnkTmmQsRTYXszfYkAC3IJaXaDohsBDbDi4PpprfwxcCdk0chDfbUU6
g5knwDa/9PifEjIsxQKl2PlIN/YGRoXMJXuBB8jRVaryD1/+yA1nDCTmEJcpk8eFPLpNgi8NzT/9
eUiDLb8kWJXzX0iE/0ZZGtDXpOzzQK32Ea2+qDfEeYzvubApsEwR3VBx101AvfudKiU0t7Y6STjU
+fKvcXku00/vSnPt7qENoF2c8Iw7xujqLt+EnnSXaIl9r+wIy0+wxrLD7fiapx5tdvYewh1V49Mb
Na1qUMg2/VbtfzsNtq0vX6xnWqj7MxdcBIiIg2fcMtqYdxCvqWmnmYd84R+oX3U3PIZclLXUPitZ
iScCLF6lIBnB2CqHKQFQC+HlgPM2vcLcnG5jlF03N9deH2yG6xNGphJDgKA7FRqKTemlM5Qlf8eM
EKdTctvUOGe9wsdTYtsy+k8zMAtSzSEgpPUG9NmHWp4k+NNo3zI3Kt7sBitLOwqUTp/N5yYETMqA
T0LsQJ7UYnOqXIAv9iNoxI/U0Wp1V11vUXjdnKlf+/gf+0S1X2E90MkOcIum+rF0fVARqwK49egX
sd349x4z3YzXlMhFyrgZAAU3GU+t7RK1yAfyM3iZmBJE5azs2zRrtJx49xCI88v5GVYLZMGLjQt6
1QPznjPuKQDY5ohykowlPny22QNomG+cKq9Uko16Gv1GmPl11LYSUEtXsyXwrcRTxpI6oET9eL/R
1jL85qoC8HUyGIE3KD4OLRRF/+oLCOv1ngjaRFHH2HP/VyTQ9O1QtR/FOXyLOP4v3IymC9sH6jTb
dwaIcfqBbAstS6aaSERuft6D25fKUdrszqBCPAhMAUggG0+h3xYnmAkPgvsL4uyXIHZkmgBv2E5Q
PQfhmulGFDfSzOtGBlMAQyRxEF36mPJNwzyFfpSNU0MgGn/2DVBy21dXLDaZwTnu9X/Dmz5Xvsb2
bbcbayuqeirtZDU1o+eUm050g2L3bMU/NJ9k4eMDV6c9IchGDOw4wGZCq6iL5Ty22zr9UCjKpd1b
TUZ0zoEhp6plv/rf3w0N5GzAIprbF1vIhykB0ehBDTq2deCP4Z5HMsC9WwT/FnTR+JRWa7T/27nU
vC6e3WSu/Ky+FYBw7PsD2bj/Z37R4w0UQF4hgJHxyU7V2+V3dfGDJv/T/95/o4TybtydQVG5Z3YK
u0SifnQAycRvlMeSS+ILmYBq5YQU52xJEH7Rrwl2VvgSef/cNicXahJGKijOfM2UXam6yPGYxWQD
8nJaktQ0hR/WNiuWbaIMOjrsSssRZ5G5MlT7SscUSdWYr2PaJof4w/CJ7VyGxhn8EOoa1bY+Pc7d
RKlXkvRcLe/NhPteMFZdcMbicd4lQ0Tmi5J3UzTUax+7Fdb9NaHn0Wy3QPZ//l06Dc1/NqH+O1xC
OrdglLsUy5+i+mLzz1mA3cj2HO2fXoDVFHr+STxjlggwrXUORvE6fpbm4UWImIgwpBWq76ij0Blk
FH46WTrUtpBCw9IActWs4ScMZKTSzagQiyBNOH4TbvE/Se6oAUSUKfXNMTKjYgadvYb6w17+BXb9
Nf0RUL+WQzNxt1bujr3BN/iudcN1aFIWRkZpSztQl9GCddwsiy9GJlrPH1LV+CNz9hfMfJQAFEbz
uRlDziSYY9oIUuimLn53w2REuWrCeQhg5gSgCE62Jh/WnBLkTNTWcDjrtvR6XRnYPFvsWuyGJWdd
bujZtTnQQqw8iFsb7lVlwjOuOmG6osLdS8bwVNTmZafiaujkve8hRj2aIH8uFaKhNk5AtPQkTTFD
xZp/XV+5lkUil9f8lno4avgAUovl/s5mMIynkNHRkfK4L5KPShIWO6FNHpdhigCh2wpedVuCe+F5
5QsmS08X+8J0CN/R6GZANuNCXZdMvPQpRhOIb0+U3FI0Rr2q19qjmwdcWtFW0SjtCHj2wYEJgjcU
3GnBJy5cO9ui8tfnTab32GNuq4o2QmWi1w7RE0J/KmYoURx81VEMbEUbFDXkFVlJdYocjY8fyLIH
3KQW/MZZQD747G5o10dus7ANnN3bVP1uO7AX7hPyJEoQVekGww6CkhORiu0gIfpeI26X6a9fgu6g
1yB3p7vMmw76upyPlQqsaaQGgFRf/oYvNelxCxh92epdi058FU+Kmc3/APaLZpRtcwA3qCvh+XvD
mB2QV8/qgaxVsxG2102j/hKp4TB1DNVHS5Bx0LMWOevBVbOELvIeAWawft5G90o+mUkXsSs+OpUk
orQ1r7eVMP3e3DGDFovDenmI24r2oXxGqb7f17c20Ql9ZHRZWiJz9EeuvciOhVRhTD0YyDrTMDB0
lo1nyCV5Dix7lzeBrE8wPw04VQq8EEL0Q4Bp86IgQUfNgxQbmN8KfgUJXIXS3/POF3NvWu3eas62
Og9gLJejRW/IcI2uL5JSGfoulCPlvYhrIMsI0NmZN0NK/nU4jReOBzTQqjAtsKx1zYmbHYEySzj7
TauWaC0bskBmW3EdM4LI+rseuqxa+NOLn/j5NlneGKwvGJBnxReHGJqhr1MhP1cCp4nczqVrZP6V
Evq5e79YMrnlT0nvm+Emb5ZNQhnarbLcIdYeGXURgqgiIsjBZRKQlBaOL+vsq2AtuVZUlLn6kbWE
LSfAri8Y/imXOQadJ78iSha0C1Cb7x7gtonSHpS9SFOtDo2WiLZ+634PR+fwZVax58u1tnm0cEQC
R364+QVrQjvHBOb3nkOvSty3OKkaVngPm52FTa8mwuxw7ESQ8a5VT98RV+TW2b7pe4ov4tIdddIZ
TiT3IFB9MmULDy/SGyR9NSDICEErzuJ4XCon518byrKuJEMK8sPln8pQUZwvY2JKRgBBmSvNeKed
OPMQ1d8hJIXrxqR7FwXUByK6rUYGW3GjewGyxOUV7ItRlREt8Vtjf5kwFKve7Dlxcj7y/chVLqWn
0fpWf0jf8EALyATzBu1Gr9Gc8TX/vhwAfhcJKFUaLmVrrIBQ0bWhwSafOtG9qIpDldMqz3o6PhL5
1axGgN5moJadFIqwUdRIIysWmeuIjnKsXKpAVeMhiAac0faOJqVLUexMrB10BL6/USxL/4ix/yvZ
Djph/vEzA9EeMRy7vYjW3td/Zg7WJiLjPEL1eWF0ZGTySdBj2gIcAX/efsrqjnvrIHJmac+h2mCB
VaYf40zLTwgRbhfY7xXxvGW5gCj8LNzg4ZCEliJ+mr1uey9KsPFvniVHXb7xyUXqCqoa+zLbkMiN
nw5IdAz92ZwqawfwTbI0Pk6Y7LfcMkW03c71WGP7RmLsypMThOqWfNnynfpuBXjZLZ+T/pM3eo6E
jAjkMJX7xxAR9wTPeWOM1Hg/v2lAuU8iOg6UO66WreRCbekRATHZ1hNdVZ2eSqiJ75vnoKxBJP1u
o8IFARr2EHJUoprdJOjQfgUyGDGvqQN95LOFscavJghg9//RrLsCdRuV/m9+KuIjcQfZGgO9/GA0
lm+uXeEUZubCcrVm6GBMVyuenLV3u7Av5obf6eTGDwQZfbByVJssZ5Pq5EY2UGf4tmJnVUQTB6B6
b4YLbTR3u6pkEo+jF/HwRmT4+s+SvupYwS0fPwjBQOVBcDTBbZZkZ4LYSyBclaUQXWlA3RNzfBQL
ddBDlejoKYfmJ+QPmvJEfYvIcNVCiCU26f5RBkT1ExkHZncDuEiTxbYQqdY64kDnJKJ6t8yY39Hi
aevzhzf/sLHZClaHGVL0OEe4XxilvqJrdpEx0IiEm1gcAamr/9ityfembjk3DFUkuKC/I/yKInpL
hSmJUJYtg2aoS681/7bs1PMz4YLcb/mBpoHAqHN8588YeApGfwN2MTEzNJjg0ez6iGIwG28eWFym
uBOLauY5GfXe1Jc6usc7vLIbPadkMVekDAmWIx+EmA0UVQMPuX2XIGWY+esIuroTWZuiwETqRInc
qjo+EN+z/UCXu1JrbNiKFjia9cgPmy29OkYzrZlFy4lWWWANedyzhp0SUB2nOh2sjVW4k2rbNdZ0
U5FzG/lWJj/kI7NT6ED61oRqHV0G2v/adr5Ghzb5H25XeRkvSyAFABQDU22ZVEYYGJ3Nthw2CBQl
4wQB787RhNir3yhJrBCzTSd7MW9za9IyCxzfHK5SP0/4aXVyifKcvx7luKzEuzzVSx06iXlBMwE5
jzoJbt6AZBwkBI/XKeL11zJ+KclcZzRIQEMbqP3ezk747rLx5x0uy/C35dgNUdlG84S8PO9oKZ3J
1UOv3ix2Py3hOLA8yPbdAoOmD92LT6HGQaIxbdBmylRljNwEvmRI9FTr5leCB23mmcmC+J8dgr++
w648WzBWq8tfBUdyUHJyekuD5K3THL+lYk2prNBie0LWIIBQhdWbWCF8QQ7C1LZNIq4BYYIw83pQ
HkQtAfQpq2JM74WgRKBNMmrDYCWby6MRIbpMQQksAfSVa5kKnH8Ora5mb6bNriOhcZMfqO7rnIKR
WsbQ0gw3ePD++QBynFNhYkaJShR+NOAAsNx3AcGTpdQRSjmwEfxoM/32JT68tw82JSnuOglg1aj7
K9pKHEN+gCJgrq1o1rhz+PjVdpoxbsprtML24El7usONBoJMa1Zo3QbAVWyJZtADyxEC6GNrMLsL
52FOLbz6xh23i2WHu+1jBnNsj5QJDWRxn0AVT1zYFcfL1AbP1eF0b//luHfivWh9gwuPGiYsTOBK
pd7e8aQ0XlV6r1P4HfPLW3wgzVA7+ZAmKAbVAYwuOYFR2qmjwLS5dc5QJtBLTByjQuPjLJs3mVdr
4VIVSeSiGJulCEZ5D+YpD/I5iAD+OTyIQvaQSswckD/ofmF3NZLSYs+906Mh2L38PcanuTKpZvGw
VfDtOfl3XzcY5LxWzRugVPTT5FsRhkCx0xvMrBsUh+RBLJR2gNZrgqNsH9IbCpjZrO1cC/QRN1r1
qsrVxYR8jvV5Bh5H7osYeJ0AM+vu9eg79IzPpH1lpEGNsQDQyjHTvYeYY9GP2cp089W7pgz1BoPk
C/bDukbEzi8ehSGv300+1mwMLZpzjPtuubPIDFJHDXtZ/bhcIY1zV9JeB2dU8jGHsaSdp8ekOc80
k0wVRhAG5GikbLMOeXRJb0d3gFYVAAyGnRQgKNauDe+XT8CnZdKe4HxSDujGI5Scpjkx0lkkZm6Y
AI5J2qeadZalFwMsHY+pT5O1yGM58iQsSJ66Cd03SVv6EPSgrugXaRkGEEj50JFHSaVXtqHfVS5f
Bb/MzPQBuImb6RnE30spNOyZ5jTE2q8ABECLcg5qy6RT1tyKRWpO+cBXVXBGoCDB57AgE4A99crB
NqYsbp/PytgM6gnkxuQlmBZ8mASAJhvmVgAaOM1MgG5lu4mALuiBWzg2uRbXszhhhA+k15+g18Vg
MpdQoXpwXwS9/PKvNX39STO9AKF7IwGdStFMI1pJO3MDKWvOAmyJkBTJUJmi4Xl46AO8iNrf9mSp
TJ+6WPZbHxWK6PJC8LFPdqCggYVpl29kPpNyDeOxRpm3nofWJANubXNbhbYyauzG+824NHNp52Mn
N66ckwzaAC5nLMKTTuS9ACmXdRHEUI2YmyX95a/7ah4qy9I64eiikjWD5HBQ2NiE6eIGMjVEqt+A
F2S4Uc0WDidHrfQprVCBT9Sac/mTGgaOAVMNPCukYFVVSBkc7P8ohPakItR2qZcCKWt2Fs/KZ0Pc
z7+gOTPRrjtA1qoG0dFliF1OxFWyGEiX8pgYb+W6Ln9DaQ6BBkNGQNP7asen33/WSFDBBwJ2tKnZ
Wwr9KTjqnMPvhSz0jrTK0xdOif+sfdFefHNcz03rGveocxJT537pgpoVQjh0HqhIDRowNLBDKRiX
pUMwErhxzSxkh+s63e+bP7uG2Ta2jUBGNOqFuXzXaiYDHKNw6v14K8kHvftmxIjoOABWVklQOOVg
0fYYnMH6YpTT56upWIXE7tbIlqPU7gGPLvpv59xACaZIusiIMUGzRNf7Yq5rjJnJIUKJd6aVmV3f
ZofipZYdzuQwHYKNjuiJMZapbuz9bDwc9BbE48TvXCbqWt39E5QsAv5cjGqY5SWCi3ile3qpqQX0
w+AirIMP/hbZvDsKrhoebvii9OGCjwYMzEppqjl6VHBr7z6yMYvxM6RYR1ikDhfheycE3FzrhXeT
OBNb/qJDqUA7xi8apXx1cF7KS8hOfG+QKYQVdcIjy5IY9GzULnXmsRz8fHv3cpHfC7KANawojRhy
oZqmKHjz+jYu74R16pwpKxPmMvvODUqAhvm4R/lw0QV5Lu2VYBKGhiOBAbz2MQe2ji8O0YK0w+OE
AwpgwHfHPgFxfN5eFETzYFNR30SubJsKgOqrf3isuPl1AK+kCz8ae7SU77SgbX4k6hx7GR8Ep/QM
06zcXZ6+fCZY4Y6/9DEJsBV8L6HGTgrl4BUpfUyszuxakj7BTukJeMhTxfvZ9D/w9ac61r+gIJiq
/S7ho3yONUws9PPLbaQJ7/iI6q5FP4GOtNr5MYz50X1QFFFMcKIr/nvmiSY/oAvExTYuFZitb1x7
f0Q/KshbuYbgzK5e4SCDN7JNd6K3RDqhXhR/EUNoiNvV84+nIGL7xZFX03FB6uI3hfyy7S5twdF5
AESglA34QSbtbxsKQchzdHIQz+JvXcjAeTLTWIv3AT7j3Ewn58alz7qIWYawDo2eeGOflkt8qNId
u9jDNuUsfeBCkhMHGgdCAIhdtfIDGsE2aRDXDk3+pTn9mhEgBwM1YxJ+uoW48s/Nw4j6sRTZx+oJ
W34raw65RrdRmx48mlFFMYUPlX3lxlamDQQaKms3mOgajTxd7G/akSNNBxs4jfvAap2O0dwdqDAw
cN6F5LXlr3BhxsXkMM+D0rHR8ANF6CH9BiHU3eO5eb7ryWX9/zv3ceEOYixLxExq7H2+fKjqGJSg
YhBQ39jUwuT7dnvd6lo5XzAxy5vdXe23ekEDuHcLTU6qBWy1Mxtzk+3ZQpkCrwzZl3Tq4bh8gDKv
hturOpPj3I2NtSonik9NCQqX4jX+P+FaV12xwJh5khwhx4QKqiMBGTcC/HeXatkDtcxnwswhV0UH
lerZSpqMJeCq2k8qnz89WQoiexmXg9CW9KbobWVvpiop3zb7E5cpV9clRuZq3Z28Mfij97uSyoFk
gokz/7WkQlyomBHdo7FizBjyCRe4QGuyuFX3rph6BtofAcL0GC9zEObViyd63Ke9mpx8D4l53JNX
8ZDMYawkUj9021/Q7pBXtPMBuAXTrJEa65c8YZS8b/YSTCV49Mxh7qSeutBRxdtOsJv02jKkcXK+
QO4BLLDPBtITpG0DxAWrj1we0Y3T8XoBjDHAbaX9IMGXlT95zD0D5wfCVLN/WaDxFdeavbH4ZzMy
nCVY1mYwpKQE7cNH0a3alLSvN+pciHP0dbgsndhW2dNpkBI/GFnIP9ExXN/5znSUFWOMgzoidlzw
Jp17qfPneFrpWY7AaFXmURojmMaFW7CYfNYSfsWG0JZD716u9XlorkOaVQ0bX7HpS7/PgSgiwSTM
wIeTMPKjDl/OeDY1QAyifUZxdC4LGfDnjoTOqFkIFVWKhkuYBO1EItHryjvtcW0HMm9XiVSi7Kzb
f90cc1jI9at2ZeuayTDPGs0C/o2az612A7kdup5eo2fOY1ynZcH4hwXmgVFC/BQ3xOnU4QNXd45O
+S1apTpekunhnbcSheyGc4Wae7WhIG6H6qz6DhVrNEU3SGWJ448kA6VG1XpdUbuGTqwVbU+ZMpzN
R4BqykXgr1O2ZSgJ7p0SW3Os/+ByvkYTMDU6mUoTrPSdCsnI71NjCWUYLmXUJeSGFGh4KZw9nEvQ
LMLQCfS/ZT5UqKjCpoHmM8M6FQnJUea8akf9hhLqyvQUb1rx1daFFFyPgSUxDTCZZ02YU2q95WUA
/nnSnMSObcRxEn8ZsUOp8rCw28vIVz7tnlv4aUNBpuUgsGPISzMJeyTk6EGm8Nau0hVYF8Vruz/1
kcMv9XDgDhGUkM1hyRCYj70ERZz4HRYZ5CJhvta7DkoRPaZkaK6obOqLy6m3EUnMPK+fEcUjRdSN
YVp+PFeLMakMNrlsJ7OVigdTyMasMUaLBxRAa0Ap5IJyM4S3Q9rT+tZ9/zGuUFlp/iNHol2OMWo5
8Lx6yATiSkfqZrPn8a/gAJ4GVtDu4nMlTx3RjM2b8topcOhWntN4oUUsIhgHx8udHL1x243flDHN
5602TMO6nC6MijirPknbvlBV0HyWaF/PzhICGjZJqx6N77jRsI2XCXQfT5R5Ahc9YOyxc/moGN0g
GETxsLhWlxAlht7ujkVjfWtFFZFV9KcCaDOotqcwrgs/hAE3eVLM+vG8GUW1JErG/EW6eLCdpzp5
pXkY2VcGO72K6EXJ8GcxCNhqKDsn0lUQO7QDke5g6h/xA4EuiCZ4zA2RUJ0l5r7/ugl8u6y+F3vr
cNMBWL/jAh/91h3A02jWyk7R7vzOcNNsIFyz7nZ8YNJUv0lzU1E+KxR/MsFtvn8PhYDrVtFm4Aeo
TS+lNErzlsquaEnBEH7M+io2Fyb+PHCW2tAFU5HgXT1rRD18vU/CfdJc33xEbmIf+DERJfbtljsV
JLoqp7SSSbEHJHL4iu7CErrAtcAJ8dndDED8V18BjjAV2UYJd5DMeOUDC+eo8jajFSgAUk36OjRH
8IHmlo3hw+PH1sZRm9O93iccTU6Dl14/TkupeiFcFGlrAUMmrCCQ7AhTHbUKL2vL8HH8wDs4dwoE
lp5rGWhMzVAJBICGEHEAF7BGprAqaQMHDyJnBXsytCbbuvIVLZ6YL1YK6gAtcKmLYPnuJI0GWVXV
IhKd6HdRyoVfzu1zn+IQJHkrcrJE8jyCoSP5rKjPEDbTJ1sNTsVe8BKh62oHCUhRNgsn33zAM4tf
/li8pgdkIRb8bKoNWaM9KlQBvfRROHIFcrMY9eetq/b/FtZcYz7FtsEytqOH6/IMNjESqm964CPu
Wsp2DsAKpuaWbsSo6Ou9iI8HxgKEBqxA6IOGivAhDXJLEXKxU1n4cZvAxwJ8YuH1e/gF5HsL+hg+
cX+MbvxCSXj62vx9hjSVJb8GBuTWyP7qOD+tnVHDctLYS+RD0Xd1uO5ARHPVsa+mWppeTy9IjvVu
vgznKn7sffiHiWcAS+ZsGtttcS1hbgTumA5ob6MOaH6rk/BJZl2tfAvkJchr7rOpjou8SES/qJ5A
4PJUbEMnRSy87WQQtMfb7/LxwzyPAEr/G7Fp6ANyBfpnqYsyqUh2o32fbUuSpvEblFG00AVKT8qZ
zFFcsCRq6XX3ZhetCD2gCrQk/JN2qWOCR9MJTDgTB0yqOcT8prJCKc7bxFnZTe70Bcro9K22SoOi
DjHG0fNRhFKjbu3qgCRfzaOwfD/a+xXxB9lWVqpT8Q9gw95x1nRhS2RnrprwSYWh1k+M3+frkz8z
klZ6AkTVE838E0itplfaPKkUEv3FvFT5sRpMjyj306WFLebwSVkJUiOa+4iTsGUgzILypc7vwyQV
DJFR6w5UWppVFGRlGoG7vgxMMCR3jZiU5+P4JPXR/jmHMWbBcYWFi4ZtjzxSyasSwq+9SugGsy4M
jJGVzxMXBUUYM6eejgAbdIPvHxXmQ9hlAju6wCGTCanjYLP5fVhWIQv5K8sRnhp4yl/T06YTYUIM
s4jIWO6lVgWXstwgpDjgrVrJeqSGplf+rZMnr6XXYCIhQjfSRfmeCzPOKO8PC/41q4mxntPsqrbB
4enE/rrE+gQ11/2CVwik27/KSlbzj4NbxOzypg7H1sqB+SqZfwc75+ELtvfU96BsjxZou0OKsTVI
KsSCXWo+si7jbNnDZr5wMA6U5NEXcp293nE4gA8HhLhAolrrLI3ceXQ5qqXD1rRfyhCurt4wbcTP
EdnnbXyziBRajWo3Cm7Fco2Fbqh3lT88A+e8cIxC4FAJ+B4HWsWxTWDb7ZCd2fCxlnJ/H5iciWvI
verxxs5Ct/H4q+K+dk6KnMbE5gL7hxXySVdoYqj5ePNGQi/aIj2pxTBANGuBjc1daubKN2YLmRmV
MA6WJPoU7iwkBrByrpQaA6g759YoBG+Q41PvApiVBqRCWWt47knQ7AxRWiSl7+5pW2CYYOssI4sa
7o7SIay+bN2K61nxP6Cs8OwgiQhiON2gVwIyLHXpuDY9kZ/AMxqY2S5ID9+ZCaGl4Ok1OK8OTw/a
o+LxL1tHgDfvoZbjY6WumJ5EENQ1QwtcPf1DnvlxIAVguwQD7D+mm2CTi3Cv5LkqaSbLhWQQ8IKe
lJLHM+mtivBdwJvG9+AgDLD74vSrGVuDIlSShevfmhp4M9mUwFQtYOvLO1VOcehxGjFqD/daH0o3
hC3TeX9aXz7oHW4jRg5mcOps7Dw1ylwsaA1AL2Ba4qW1JsMvdGD3vEn9RmdQfGg4NEfBTqgw4p5f
B6NKpDUvPSZppwATpiT+WFqINxjOPRt+W6kWexJzHE0uU+JNJt0VFnbXL9ZZtj82y5DUCRrUdRbL
opzGVg6Dsq4cmY9pzM5iNQav0EicyhP2n/HL4uREPOzrGBxLU6y6Nz6tizSXcDfJ/nTMyAFPeCDJ
myNYZASVkhobT1a5QVXq43al/xxorvL9AwoC0JI9KOmvW6HIQS5zsE6ItdraKR8mp0xxU5//Tfmt
t4s8dgNUanMphRDYj7XMMzcgXrvOxZ8crgm4OFrYhWADFBNi4TGApFhkjHzuILDnmOX/axSr1Dwj
+FrAgz+k3poLDdoQX/Piivo4FZXSMBTdCymF/FjiMZKWEQCoUyEzBDm+7lBK1nIy/dAxfqWdI1sO
i4dYPg4tWW2PGBzrs+FwUMmfcobUrfTgm5D2eApM/W5vqxuhectep6R+7OJnz1dJJpmMgAvVYvkN
fyB3zNyraxJMCnSJ248t5x2bPqteF5EmiMJwf+mXrQzOy272xfsfOqiaZyFIZntDkVyOXotWCn91
ir9xA4FY1u6Gf/TDYzpnz1BCKlngGXy0RogeFrbuyPbX7h5e78iaSCpPbzGplp9gjZGgIGJVp6sj
4u8glalfpigq/RckBpFMaXvPlkrSkbfRYjuFHmLBk2Cdh3vRjDu05kaPUk8jZNi8t8FiCROicnZt
PbTrfzcYjATM0rqWJV5c61tbBEsT/KltLzm0Kj1zHpRIVNjIPm/Jhh0miuRtREmya2jyfOU8qLJi
1LqPmfMvXQjz9mOgk9+tmz5K2vhQ/Tb8evb269Q3roxSOz7ah+QIpoijKAergcr4h+2NXeFwd4Z0
cxNaPKM76jGrDz272FJkMtD9QM50sRChS56A0j1+tgogeZEstFxLU3q2UKsawXTcKBNN3yOShriI
ZcqiHePhR2sb+d0DHDIn4tn2+UT5hCZWYSvfm7efpqy4kottfNZ0YeFlGFOKO+6R6oPlDkknDizD
6FgAkD0dSmF9PVbL3IiE0QN0e+WVRHAYk1770yMiWubHvZXUyugBintXOY08S7/KhW2xIs0+KFYP
+MV9bkbGMB8rnREBrPQ+7JnQr6gq+I+DGCl2ohoseMvTctVXBOhpAwOohxOx2sK0Ptr9mj1o1Nrt
pirsmAQ61Yomm4EyY2z/TqrpJz066OjiRmXxi+HeKNku4W2mUU2AoIBc6zlw7XgIEnZDgZovT+OJ
XddCUs7CYPF9lRKbprtS77crKiyHo/ZTif/Rn/potMn2pXnK1iAD9g03DNsbrhoESOfrQoJ/SvUV
aB7yetQ+uZO73A0UkiqTKHnfKio/ghksr0mdeLEjxOq39rAARbhRCXdGl6Q2EcY/1Pr3c1ZQ/Q6h
X3RVi/rzUG3pElKOSaKESGGk1UNu/04EXIQ9jlApckZUO/qXcCPcSujuHOVp2wxZxG+fpX7dn5p0
TUsMSJB+4aIER4j5oERlLLVZQz5DqdWauKcg7TQ/IniHNKSjSFcxDj2FkG+TWcSR4oJ5EQvE8+QI
dUoHa2knzI3Umve2zydDl1nlLuN9K1JvLVNUGFzHeh8FqF1zqacAQiAtn9qtUJZ+3XL56I7S16gN
NAAl4r8TpLMKofWVAfqhrkon1fI/LpN9rIILlfrScqRKribrJBTwxALvrbPnfSj8fEzd4FfEhfVu
SiKWK4BBMBXbDKe2qaJ+25Wb/wzIBbqESnh5DtZDqBtE/4SJ7+EZozqF62aKXEURClUf6Nqd1Umm
kCexgFmd891+m6gS16I5JR+ableid91ADZNaU2IAVBIizvv8Oi7J99RqX7q145dDA/iKdAnvAZRc
GRCZI3//YIO3Ctr2aYAROQKHqc8kkeVk4JaRHSlIrToZfTu/G4rG2oztgv0/joMAlV16AqaY0JPI
tWjpl1LTV8bRWo1fEGvQaaH0jg++nOm64a6w3bDLosjnK12AfRi7Z25xl7i9dSih5xDtMwOFhl7B
sABTKYUCLb70oBCrdCj5ECiQlEie542pTRylcolxXoS7bfej1JRKSL2T8MCMaCOnQP+al11p1oJK
IxxoS6ccQHi5PmqDeXBrrwTuuzmdUWliixdjbM+Z+nxDY4ofJKiYU93895BuXPVOpfhSYkLZkRu0
RLht54ye9N+q0SKlM399bhRsiBtgRdawa4695QTvFCEeZZeZjiswc+6jBYc7+ti8LBGOX2RyxbCo
XjnQXexFiUzAxmG6T/kqq0U/GwSY+V9zKLMjFvWeE7WU2Cu/43wlChhF0baVPtrpNmAx8T+FJFx9
6Rsjsv+yC2ZXrSBXT8tA0BY/bMu9kmsOMzzpcYG+Qnac7TvygTKM/Nt31aeK5LMUttqPdYDqyRFf
GALgtFxAW8F/AxqT/4+0s4PS0xCe7J3eVu9pdqlefKdWnUXowrVmguBrHMLepiH11FHOl7kF9e+N
Gz5UDTVkkwasdHSDmER7kfbD5wE+ZMTLr+7S7KbwAnNAfhwEls9vUH86MisKBg0NbUFlxSmfYj2e
/9jmfHLHjeoY1B8eV7ppxXgXtkNwA+4Nb0/EdNcYCruewV+hgAOd3gjmFdepfXXMuWpBqSsVkGCJ
wZGjUujkThVr9q2Z+6U8iCwlBLi8mnPYb/hFver05vfH18GWvqfRiYPVWPrwNLGkiTaEMSQMVm1h
5yeUzC8CBoOO1E1UCRon8uGGmw/zQIhROEorEvY8YFR0HxxySb1eYMIsuUQycQtOou1Ogci6I2+v
X8/qNknzkT2i3L9vpxjhjoFUFBa90YWnXrYXQ6VFS+kOZdMSKCzrg+DBc1rHrQX24JO8352oeaAh
W3n/oeo2cFHYeBSTpEvsL8K1jvt/grdFOM6l72nUU3j4cc5aEycqfrqIvtQgxEo8h2jPWKr0Lr0V
/mT+GlFPJnjalnEKtyCYELzkxfArZnrYLt2pGsTH3yD1vEyfj7c2BX69Af3SiSnC1SHtCkQjGe//
6EBQEnexeA0TdcMJkj/YBRf5EHp8cm58yTNTDUin/E4sXkmHCUBf2e30VDnVAkljzBR6ubJWqFXh
WUVFI26DNEkZwos8lK4YSs0eeqn0+7nAC2ES7BuGKZW4NmO2w8IEQeok7KMR6/MSCueC860OH76p
u94J/m3r1TH1Q9WhGJHASecs6JKzSA42dd2PPhPi/ZSDqnToweTkIaGEird61VSHasI74vhIwdSu
+KsMlsliOtdt8curx7W0JP9Syz+m+Zp3RsAV+SFO+3L7tp2o/xNONBo/tFFAYKPPqLcWIbMLp59i
Aa18UPs/pP9Gz1Nbw3DmSyEG6L4pZhofMRA6Y75my889lG/kfceppXGiGfFVe3VBO/RBcrM3ddD0
+J+LcmYOZ5Rrw/VnlBAxVxQPBYdjaPZHgYOYDryov+BkizEymRlrl8Zh07caVv4glnGY3Dr7bdu/
/OgDinLDMx+8CgtJhw3cSPb50R+EOQ6qzJdvvlkMhUI+IN3d3IkaaANfmTJa9E1PQg6ifjpDhYur
fapEqAoyJm0D0ZYOsIhOP1LHpp9wBAqc55rYiMyA1hYe6r1lvCOJoguGi6vei60iVdKxK/JKfyD2
QzOIsZscYxJq7i3B0oPQJ3bCSO/71owSOrhx+oF6SDqQmVOwYhuiLZGYE43cjh5w3Yqi7/PuVsR7
hZGNegz7Q6cxSR/fLh1C5lrgfRlVOFb5nDFsMKKFT19fPMBD0TgJs9ZIeYbwCK0ANwlSL4AaXLoE
kqUILABpIa93K/BcAsvOYvm/REoYwZZTeV1afUKROlsjQ4MA6Fr4PKM2UepokkzAFjAgBSuc5OUN
MoCBWMJeK9dvoX03CwUCXfVnCoj3ML9G/Dmop1WqqUzs1Pmwwu9a5UZgvrOH0jvDozUOKqI6D4es
/fgugbUEnCt3HHpKNMNIIckslYHLAw+r2sZ1mLduiiyntHSRe5XdcvrH4x3jZ0ZXk3rmkxgsToOj
VbuDlxt8YkXHBF7pxFCIwnLaYjADowhISveGpQQmBhB336RjPKf15HkfjgdrXSyHLRbwyc3hICuk
aG8H1CnkjTl1Vi7QAJNyUOpDpKQ8A8NEcE2sxSadCEXxa+r3aUzPuObimus7iOaEHGgLHJ81Icpl
UF6riAdj54e9GWGqdBTPm26vcGFLlInNaug3g8XaaOequ9ypwabKvp/cOvodcPtEymyJ3VsToO95
FqHdfeat9swGe2z2kwcuzqnSgaIqH3KmNOJD5bP6vXu4ahWQoH0TspfaJWZS2mjyQy1tEtf6PMDv
GNMrpJdca7WpcDATdbQ/8zAcnvqS65kjKljJxPZy4iaHDtuUiFG/F3cTuKfQxZD9w1pYsXVazATi
zTPkltP1njsEFBHNHCOaBBLt+l4moPKS4sPE4Plvf1/HeWraPGRYjSxvdfn/QCwg3vJDYv7/wIv1
t/HZW93bSaN4isDo5k8PHQykKGR6c5NFXlW5b+d+UFKSC4klfFNbBICxxpYUWE/nFaDL2HCtgIwe
c2VbOWTnxbRGXrh58n9sNr8Gull+EtOAFdxQUL+ojuftQT17Gr/D9IpKLu/v1GcTVUEb8/4+c4Ni
kZX9dWgoyfZVniNIGHITVSTM5kz5g9N6FoS8BlxPMlBVJYHnfPY3Ay6ong0q4YoBoib4Fu5xEYsK
3cChpCCQUPsyXatLEFwppzhB/pVzr8cLM5BipRP5LMWy1pN+wyOh1nLVj3fsqzYVWcubEjOG0EhS
vDr3emEMnBGlFluhW2dZKWqAUEPXapdzAIWqH9gqb85WC4ysEMjEnQBgNY6NwpwQ+xcXU2W/hFYv
JdodKdAnL1FcX7BUt5pEtPlSl5IyqUC7BYiFDQKtxNAims1R1bqufD9a02rmEidrx1XiHddoFdTv
XMvrObR2QdI9ecKXPGwQasj5i7yC9SerHA36dX7UgppGqD4KEBYHawCutRdF806nJ/JDK5Rafgni
YAxFwKLl4hgu9yxdCqQHE1/YNAq9OB3zejf8DneyKCv9ML3i5Rb2GpIVYXGSvLmgmfCnCfSohsae
TG3Zhuiv1B9Rl60DTTZM6GL4Hlv6AEpd1WxcqBzzDNc7Xb3WktZL6nKIrUnxIhWnwZ3xByWdGq5e
ZnCtE32ADO1M5PFUfnkU8GUhy1WWpxEQUlNoCYKT8YncwAyD39y9CbR9540Yna+4QFn4YdGUs3s8
J9eoH9IHMIr7gbpfdHio2UWilqGXsBiyKo03gTLDK+Mxmau4Nq8yKqk7o1W8kCwyFbq/QQORn+fD
8TiawmsG9izDE/7hcp576PD5aeVLv0/tOo42GXXV7axu8RdFr5Dh7mLBL4IU/Pv290jBVQ9iXuxI
zHnKZSmNfoJpoQMJqDmcW3ySBJ6ktOo9mMfA/0gl10HZr+6P31Ii+1bTI9EOHrqzM7adBW+8DY38
LndnKFe8LORUJ5vkoKDDdAZSADhUUJowM6QTww/Yjck9nbD/C4vXbSM0sM/HaSJtaZe8Q2Bj5CLS
oqp3eAynllAJAxS1uFxH1mO+Y2krzPOFdzFo4N56N/L6bHK/7wuaPz1g+E5bfLxSD3Ur6ZRKJzth
DsMlQ2AzgDSr5enzvXhfZcRwDFalYDQlncOulUi+XJ3a0gIMspjOYZj425Ik7p56GwTBf3VlHp+7
aVCC9AXNXzkb03+WtTe/A5fqVfqQQLdTZVAQBEC7HXnGJZ8+Tpk20/b6zSWFEXI4ARFX9eO+pQPD
QOlz1fitKEupOXi7i53mvikywGXMW/LvBA9e8sxexe5i4F8dZY50E+j+KECI3nM9p4XV4lN/Kwlk
tokgbz7UCk2WfBupyAVGYpjWT52kJKH1vgr5Ulq8gpdA7oMhqgIyMyF7GTrGPC+M7VvlKnjv39tm
eDnxrvlCUe6ol/eaj4ASrUqsFsHD2FprhocBF4ZwKIZY9tExc8iWTYSLpCJ1fi1plBOBy+cpB7Tm
8OVkRRuJQn33iNTmqYooMcOjQxHcEBSbjX+uOTK0/3aQBifVgnCvYSkD2mM3WG9NC3h3H04oeJ58
wbO38/D/mT3ffIFcXwmDaeF3HmX++Wg/gvgird2AJyx46ozTzknmNKCUGWDfmmLar76AJgfJ5UmN
WnG5Wfk+F+moGqMT3Tal0EpU43oWO3f1ZGD6qqz15p1VYDu0e4NlbCtp7FYiIk42B6tPO9Y3cKjV
Aaf9ccH5dZ9aK0LiQ06CYlp3Y9FT4r+MerYi5nFcN9mpQZwR7Mk8jyFWV2NHwgzGvrH+fXo5IFMR
lvr45Xe3aZi6+LrMjjc4uwVoHwaZGa4Ay7ARIohVfQkXxk5RGVNfLikucFqrSdCPikYlfcxBFSqX
HA9pvdk5Mar3dRU3A0X2NH8rqZKdOk1jhKZrO8ID0VtXF9tqS3P7CusJl4zbp6HrrXbxnVT1hMxf
2Wmfv1MMXVs6YLyJigooOQuGzh/c3Oft2l13q8+57SVkU5eZl/5V4heW+dou4vSPGCOAfvPxmav/
tjd8IRZJeUI4NRHh0fEPYdtYufRWIImZkzFAhoq01h52C7Y//o37QlB8l8ZPyAc1t0slqQtRyy/a
etShjX7wt+jiKCQFhlNSV1a/YhD92G+dD/DU1JdVXqZqHKtZ0oHolc857DuhdCOBmlMprxB1z+AR
dDEmJN6p6xoUxL2HiRUI/GQxadSrRSpKyFOyfTVyrQzh2kDj/43X1+AdLHfeBCgzDsEgzpqkmMt9
40kaZcygcJwxXcMGT6ot1A6cyetyq782w1121ylbG6Nu3nyNk+91OGQnJIZm6x6KEnbjDZiqwN2t
qK8waDiBhUH1N5VDRreylVgAvHa9g9zAknRsI/bcCNUKGtbauMcywi5Mgaxrr73CMaJfld8RYUgw
JqGezmKdiMxX5G+CIWwMxfWlQjf6zlAN9nnySjGP6M1w6v/kxNkQJxKztcYH0gcHsgRNHRpWgkNg
FtDe4yv4orlal2oeTlHCjbFwnogFPX8tJgMQinChWNANqUKfhhB31m8xOyQPaTKUhL3DYpZdDGyg
XEq3uOW7airmtJzm7rVfXvMZV8NHjNPXmxLq5UcqZn1TBfwKb3zpT+XkruR1VJvI7LHY6aVqsUQ4
wAPFHoxOuXkup0SSt3Iunwx07OXXnqGjrlQoEMSZ0shVAUAT2IazSPf552kkRWOeNyv8GF4F37/p
dZGB34s4YQbeeFvCkNrifWBYgyj6yKPdoSJOm/Zj3EN8vtzpVtA1aNG7GIKBdaHAD9S+S9+jAt4E
H/lKCjHw9GrtkpO69c9+MZVnmQ6yg4xQNOXxrAlPZEbON2wGtbPzzlWsuavFLh9JH2qY3wyAlnaO
8rwzlQGYbToQGOB7hKeg93RVrzYfCQ3ga3J5vfSDmm8KrkVv28vyyyw49WURaP08WuESIhKQdcbs
SuY25qlz1x1NS6z6uJ5FWadEEPpY/fRL/vImUBSa34pJssRt/tZpWbS9X1Z9wq4mEboCJqpziQxw
fI+qe3n6f5I7YpMDM12cMxyHgvIhkEfIRcC/tbaBRKP5+ofrlx/wpHguLi5T0xs0kVuqgOxVBvMu
lfXxiOoOXIeh7zgYImWyLC2XBgkQgCwEzh959MSRJ4+0w3iuZc4gSyYJgcvfaRlm09713vudPuf8
Yj8MlJV+oMDu08R/EYUq+/ImWVymD+496brvGQiZg1d6Wc2EIPosRvUsfdwamhJWvf1HD5D0KbcE
oh+7q9LYSDNF8f1ARIrD1SqJUUeUpU6EUyN9oYXnSDTL2dj/UYYmOzPFQe61iTxYwOocF1pUv2ML
TmFgkUBjrsb15drjeGY1StUL0bhBpnWpDPkeFPk5dRMQCZHIaqiEYregaLS2MEF4af3a8p14Eauc
EZ6dKFD+IVVrF8feT1VVZ7mge/X2Fd3RmHjYEnhLf3wB+GMo31zIW2iVeyVYufkye6szCDgvcgFp
wzUcQVGuHVDUBjQII06GMuLddLns8JvUhpHOUUOLodp9lmi3ZnH70NftXuN8ADVycIeT3mwZkaIN
eDl8j1NLLROXh4oFj7u/gOoSzDNBv0vJwDJG1ffZ9FPF0ZwZ34j3vHaCC4Ywp7zvscXgmLi6z3WT
8H2admcdiNATDObJ+QSMoneoS6PkTDjXrkygR3d5OVFj35OxzyDJ0vAbgqVVtMfW5LEMItPX/qt6
1HTSx/SByf4CT1UD57id28PrfT9bt/57Vw7YtfS82QQ5o1GnpwseoGFZrEyDynfxy/069u+/qU/1
LctIqlyAjQa2sylz5JYwDVKgw/7u2KapG1ZXB72ciHOFs0WUZ0mtmOCcAkGU5ZztXxS0CI7v8IZz
tNodINOOMQ5eUrq9S2drbo233M326odYenmAKCGzp7HwEJSJWHVErmd1+mnI/9MY7cLIYtxw4Bqm
FuJqI0DZc5aXonMSqBWKTykkLqT0lXGNtDPZyNqgAaAikEP4vSq86pc/guGEkqrpRn94XsFqXkJM
ReCH3jpxFJI5qmC1/xvwsBRfCezmJAYpn6p0eaY3cuS+misrjGJ6Yg3tMu8HccTiM+427RIZdf7l
m6HnoWYmHMZ3r2mhqZrpBazqTkrmmJs0aIkFvILKWOwc9tQQX5mzmCoWQv594joIrAVxSgDHAuAa
rqLuRLr1Wr/qG/H3BbfkwZDP8jFgKbBl9ru3RSXDSM3h3vPJGpoUKe/vnGVtNRChh1pVvBRjyDZN
lSQHYeMQeQEPGSShEh1Q4fUDnHiPjclMFARj7jlxrq5+6ybPXQSKC/vxeU+DF/3MD2fYvqtZDuHb
Jk84RPykcwHvYuJBGsWkgX1u5kBPS0/Ph0GBdfEOOh540kfUN/sr4lL1rVrnFP8eb+BwE03bhVmF
QzwV/55+CZ89tIrJ1eaS16K/Qq4cJcP1SlwyYFJ/Sv5SuInEr09JDCXBOB8cmYR21FZzmNQ/U8us
UeISgCOjSJJNzOpGBvcZULW+/LUYXabTK+duRsCJob0Wb+72JENVBtjO62JIJd+gXUNUGlXO/3HZ
TdZ8O8CxpAMBZ8NVGRKOGX2dQFrqUMrW7tWi48EhQFqf/9VGE9qFbcvyuasMudwHMuS6EtSjnLKW
e+cuPdZus3atVI5rE8ksIWaAQn2xluAwANznk+HLqcYUYGfJrqNiYE4GqT/jIMMf/gjmJBLb30uG
TtDum+32H+Zms6okox2jpMH6trexp0JHtpkfcOUHtWOZfFsRFYECeIZICB85TLT/f34yfEo/PnKN
4jjNEWzdS81ZCtzlW1aO5TBqQ4yzxlfpBKQYbUEQc48/cSCyDnp6Y+YFBVagofEB7K3c+/G9cV8p
ktaTWXOkV7KnN9CJoUlnXTiceX4jy39+LvpwcpS/iQmmMNN27n7+Ar16/YrjMJUNXxHHK8zTSn1k
YA41V0HiuuUEZtL7DF3b3rV8vhRnqkoX4P6emylendIyLW0gANaAR+qKbBLQpi3/hM+gOflmBxAK
8wM5OkV+Fa006KM7DkSiUkzUjoLxBfzXhlPwPXeLcyPlC0nQg6Ok5GtGFRrYCP/zUhagcR+EviWu
luCQ1Lsd7KHOaHabRID44IfAQG2EoGm8rtfQOneS0i7kVDeoZ7wO6i/dAIaSZgVxWhxfcjzNG6r+
vnvTE/rbEYmaHFypeOaXZV9SCIIAVUNrW60G2P6HYZ5rva4R+at7XnfTTbi1RztzF6yz4VspejcA
b6It388l4+S2uawEw1/qBbeAimARLYv3rmxCpEuRkuIo+HrSXQL3pEJ5C8avy+Tg3VngzMwWjIej
ynj6H1sU+ndCH0LiOcVmLrK2thT6R3EFgtrYgyw9+qjVu0TygU/ujOL0KL7mdDsfWhvqa+C/RnXV
5Xx2TiONhMe9hosLV+wiGamrf2S5MKTm62GmQ6/J5mDIQX06dlkmBvHdqIziXVxKmXSwxKeGoD7V
NSXgtSQvqCy5hQm2ZyzHJ3dGCfpfqhizd0cU2fqApZgN8asoT8dtV48yzqbl98JcOIL5JIl6BVDJ
9a33yryKarinN2UCxL/xR1LG47HNHiJ4kcNsvlUcFT+rpPZjM0amVwLh7XXt93xZ+TQJ1NNoFKcs
vpSGQNGfI4Mcw3cSmPp270ZgNSU2JAiPW6HZzEvK0gVOhdUdS8D3MgdWJYKRKhAy1V1AVg/PI/C9
arsXyh80Lz+hfHjkpHBFomkjBNfpm/EGJ3yy6v6CLbvYkLUeMAIlV+YEmJXzzvLWKna7PE4Mddyi
RVqMP3UyZKEC029VPhHzqt0Jn6bjJ/nEiaPp8DfpCZLXQx0L7qtsaeE4JlIUiDeV3qDBL4lb9Xod
MLrMz4qmoZ8oIM/tNuxppWwI3eWjG/gAprYWYULTTORhY62+6b5MaTVawd+ItZSqPJxxG7SeXhUJ
W6gTmqG2j8p6a4MYzRj67cJqOPSw5OkVHziiT6bvdxhL3DY9zZ10R4u+R65BHMpfcy4D91MUkDEt
6RWL4cc3ZEXmLRCG1lnVe4Jfmn5fia3JJEVK5x/qC0LN2zXLV3HLOHVz88ACopqB0t9etivW5lnZ
v01iuMMKI9TdgLZzB8HvJ4ejBUI1s+37OqPVa9zGUaUhWqwbjuWvBWoBg7Y6sHrnWa88MwtUtV7r
qehBsHnFuqw6fxU5P9cc1eeSz6CLqph+yhgyZbzJCjK//ErzCRwbqx/d9VfQ5pIzl37/zN7XmVsA
NDhAHPmEHUuKm8GVNfLD6hWJj1VH+W61itGVw4SQZduLOjOV0644GAjwuwc+D6NnARzPWoebm/Pp
0jwmIeJLUrYjCmg4OgFVFiXwgjd1r6QVFB8fY2y3tFGKz6h1sSRa4kiH/kiXD959citloqYzen83
Z+lsv5hp9sY+TXjnnQv6ftEu9+bslVezjD9doMa+hIOLwjrSu/JjgjWC9u49025e9JXes/5Y5F2y
zY4gZkS2oZ6qELXENP2XLOrk/zpdLghqTrEbjLSOeRwT4jYNTBgzNHC0kR2o2EI7P8GEa3J3TmM8
xcs5+uSph3hyiqbeWZ8WjtadUoJ4YBKclUSe3+V3awD+Yzz5oCZWTYIzMxxcA+s9whvKq0k+/LWX
l/NOYHdAsb/tSvq5YAGdaErKeVcNmQgo31XBKEt44TzTzO2tUmDe/KN6r0DbjQ+x0lr8AAvoNmge
mAoEeTCqoIyt4bXQdhTW/TZkALsfnfy/ticiPklOvEuHyuxMHQBK+f+9WGifcSfpYWdnRRlUxnOd
Q4YyHtzwlT093rMe6RyqjPzad8vm4NpqHq52r2ePaKwZ/57H69FNCOe/DK/2uLAyuzy2scSCwvqA
k8ybDIscYEE2IY4CNWManzDfREPfhhJ2RtCR67EM3M1nz21cFPi1d1GNxlAxfSrTv1C9Ryhk85hP
ykHWzAlWx1i0JF15gnNsPWKeSG1rEIQAEatwCgT5vNGzPpwLaajitCgU+1551HeplsMD1kVConxp
ba+Tw3JGyT3CPwzM8tUj3d76NUDIjfVJnAVmX5mdZjm1Yskib2EH5xUr3HWN00z/Lq6Qyz+REZrV
YIuX4YQcEOj123uycYQv5ssX9rriNBFg+454N6Qvbe9IGBW3YbRioCnwt0+jsLXdtJ+x7GfT6gV6
QoaI/s2vT30jQCWXMFiO6wuSbHn9rnxxQ6617AjUTWApmwhM/YLu8Hpn72iTQF/R4+UWwv3A5gFK
m0jnFgCvPRZ0MvkFftGTma9p1YSVHkex/gLVurNIhD4euSLA96Ev3NqEzbxjkxfhmOWmFEwA+4mX
vdkCyY+32q+zgBjQL2QHR3d8nuw2FSklJanWjxbQLVZ8buLguplEvgvCcE+QkLEzSMkpjf6yOyp8
GLdqv54Udgj0KKeQbtkh8yzlA3y6+taoc5BxJXrksDMJUwAu0YJw6WBf5jG7NecUWkkoLFdIR0cT
nfiJ21uJm/PJ2UZOK/v4S3+H+I5fpqShrC3vYTKAsbKhmtiXcdUxiyYOSqYwBUDpmqWnB3ed6yCR
8XnJLi8VvB2CjgusPZNqlQJfc5G+Bkv+gtT5qfRDz282guevM11AB5o1JN4bNm9kit/VQOufofNl
gBq1kCRV9xMSNB/KZkU7E3G+LMYBw+8kYcoB1dAieHFF4AqUPugIvjyWa7q4H2+3vjJRWNe8aCUr
ezaqcQ4u1N0u3D4hpBJ3QsWtGyDKD6bBZ8xd+lYVSBitd14fZ7U/YKHyG4YpJEmYXoKXIRrDWwli
4q1Cyvff5tZrPNdVdL3edc5zxdDkonaWVDp5urAHSnXDZbNBkmQ9MziTio3krNsOvd4qhra4Tu9W
ycozFAwCau7+I8uQj/qbzBA9G7r/l3M/4eyjFBesfs8yBmzJrxhdCYBFrgYbuwKIwbKkwz8IIDiB
Jz4ZdVHFfEzdhNTed9O+2xm//ELTcTJPVh9WnWXiCsndJ4DBDvuawrSiqk+wp9XQRWKwf91ewP/v
Mnwnk19NxNiRrC1M/Nhg0Cnzp/WgcV3K/AgC4Z/JuyrivYePBb99yczawSLx75qRfwjroDx0lfF3
kdZsb2AtcuTQnVo4ROk0eZL0wy6gaaTEVGOfTrgWqBAsWvB9WGGfvp7RGdxA+kGp9ebf8v3cNwQz
5itRSS+yNI8g79KfpWFSYQmdH92sCcCIAL33nigEqhoYZruCe+gcUMOE0uTkWd8wdZ0rHl4BCpYj
XpQmyoncTl1CX4x+P5mniTNFpbyIJMSBnMNXO9pjLMlyh3K7i/WOxw/gnqGlo5qTSeP2NU5/h0Dy
BHC/7xJC8Ftc115QwPJmJbxgtIUhfHuxHcMX/r5m5V3VzScy/qJ3uTUvMJlA1E4EIF9yWbeFo24c
P5NCNZE5j+VPnk7QD3EYzYOTBsUSX7yK9G70E8a/ODkx9vGd2qBZF7Lh+sJB7s5PrHvTfRpOLOkG
l9gW+2Kt0ehBpq7F6QyZf0uzOSsGwlfnf6iK32LUpII/hkMHukrFRncgoJJY6ryzKLhWgGJTY7MV
S1VzIBT2IeJQI+Donq5douaOiC+jS1Oh2wrjbeRhkvnw6dnSnZIZzEdIcJTKM61jo1J0G2iSKx8F
fIcfII0tR7zEW0pSn1SIFEZt9RyRVfE+IPZQbQVv8qwE1X/jZkPDLNnvnxaHm0rbB1d1XWPNpCG3
ia6UKR3ijtCQjH/LJPqrPO0I0wGAj7Rq8v4B6NhH7GqbqHckiQXa//6ccQ9tU1gGmJec6p7jcX8Y
jS/QMkI3Qs9gEFeWPGGnlaaUjDxQsGicEBvrpeW/dOQQUsOPGSO2PriL5sMHkt8Vn9I3RBPHM7U2
1YDmKoeT1iJeRUEm3y8GEGeDvvCOf3SuCbxa6WYFOtHTdjQZF5wjM37qWInXVDPOThpvkke/hzlV
nEmjUbMGfD/c4nIcX+sHGcB2Bh+WL44G+KnGhpWWzlBBL+YmYocMY9tUva/vzdOSo6z0p06oiFvw
OXCrsWA3VKoOvcvc5Qv0+jMqWtNpQx6sA3iFFME9RIfgPnzubJILCoBjEzgKW1eDOPIOLxNk27Al
JOaqLjRtJYJ6n1YEkKVfjuadiwBsi1BH2EZ3BtBrsNln4VFKp91OdIyJOwQtgV56FL6Ysk5gXJOu
5y6PFJduAfOfyeFo3E0lKYnXtf05r8PiM08y1sYPKREl5u8FVtFTXaBCXfkgq7qqRG3iCVHeYSzY
mdb03yok8S6h5lvX8rQTV6QRJ9tVP9qmuaVrGwbOtwJoJU2kUpjW7OgjEED95U2lrmzh5w+Wev2W
wdJVW2qDc8E9BoiiEf0szHr3TKatvVYZG55iVvS3NEEpBd4jAmQknyVQ/q/+g0NtAKnU0dllVf2m
oBzLn1o8y/ploDOUD3Af7yk1XGU8c/hAPa+I+BkF88NlI0q4yLWh5WTldXD5t8CQrktFVy794u0Z
Vj1539w7pmtXXdvrPYrPyOzd4JMmwnshriEeppNYqkClxMYS6FVEwQgU2YzsXVfSmjPl2Z6PlqUn
9181W+KOBPLupxAqUf22LHKze9GNDez3cs0KB+9PANAV38FhiTk9o8h8mlkO/vEZscB0/KU0rGct
fC0ikSCcmGjuZ0BdjTVQTnFa8XBsg3EBxpdLl2E0CFGTzVNvIjux8lFldq16baJrbpX4WOXNtMPF
nUg9hpX+YQMxfWMZ/MghuRFYVuu3Du0yrQrRELI031Pgis7d8OHw5Pa7LWubFzNHIfssjfUVhlqu
74G7Sljpbv9gK8NxJyPjxpkXJoS51TVd8tgCvtKcdSUN8Kh3PDVuCf9qb8i3AQPuhWxpjW6olsTq
P0Bn0+7On6ezrx2AM71pSKLjh5fhm9TuMhbftHU0Ye9yz2pUM6LgpAcy42+LXHJl7er0FU6Sa8kT
OkcyI3lle/ccE3fyOofyu768rBEyTSoLDa+oKwXHwlOT4Jw2gdkI8iJnSNSJPGTRssC4aDFSx/2a
bXTV2wgvG5UUzxLXw3x8+UF05Avrpb5pp0OKwiEGG4XN072ipfe5ENuLZ5tVJHmj2d4e3mqogJ3K
BZGjZApsF0GR7nQWllYZgM7MlzUWZZXRv6l0TW9kXuKGrgEiMUL9HASPUiSHKPaEDXk2QuqtNVdn
BbqLimtfne27738YP7JFqp+Bu4nGhYKOfH2zJH0NoJagZcW0v/a4xeyeARxo+Qw+I+heAg88ozi1
tbn+W8dTC5Mn5VYycb/cRh8w7264l/WO/lhx2XgoBRKWvuESbkikOZiSomdsoqRYAWXhUB8/tWs1
Gv+yakqLT38IXOtxfk5Wo+b95yGQbsdMfh9O8Uszp7sTFxQvom2PEUnhJDgBf7Aa3vkZCXuEUMRG
+NCqwy7aOJ0KKwF3eWT4WtJi4KfPmEZYL57RfQzadk0sdROAEAwXuZ6KhgmqlamdLvdd6mZt49B5
B4jWPIy3zG0JvG9e5RfYguVKviEWy78hydpad4w7dAHA5tdkmuqKoDFK5O1XD0bFYz5D8vOYWkJd
7d7XXc/goqanQ1MJlkMOhpD8pplwp9+skZCXxolAYvNbar4049jKzx+KPnRdF5ulV6EDhgyRV73+
YSfPFiB8ylckVq1GtsVoSEGDIXlopEV94AryeOtcitzLl2kYSqV221ATK/cAF8OmjHkbu6c/ZvCc
yb6IWaNezcCYJXdJHH2mYs/Bt2cg6gQQH48m0k1/rFWhI6N1zUjv3jDZZyUAk+R3NrV2HRr5YH3w
46n+smovl4WqnacVHzwZ3Ae8hJIO0b5iMlcs8Ttqf+fh5NAt1oPXYCNEiC5kWmO0pK1vf0B9hA3g
Uy7ASH08dbAyuO1HE0dknoew4egmP7Bua51j4Q8CfreCi4B/jZAzTNSHBOLsl5y8+B8EcW32dIOy
hpV1EMA36LHk7tbpKG/9y8wyxRBKe4VMtyd3iZ6Jgh0r3S6cHU3rMQwHmY3YrlTu9BUFy+k1HaJL
L5+yg3LmgG+Q/nL+wD3frtbknq9lPnJCUgMjQzL8POUlQknMHAz85gEZMbXyF5pnoaQTZd4vQ9RB
4HuVbfLPioNyzITL/mQr9u6VgRt//HBLh5ZEr3ToWVr4iK6mjTkXWRbzhNFURjv49e6FkKr3Gh0F
s5m0TngvpYDRML694z52JrTsYnId6elqBO2ozlW6TY9jdbIHCCQzE+fB6TUU4Pn/+cgJOug/d/1K
LOg8um/wVW1eyTfI5dfIuRvSXQ6ch7XT3E2ZPnHrOBljJdcpcoR8dWYa0gt3wSFi7KrogvdS5Pj8
Jt8WQJR1DgtWqstNcKtq8ieBD8dWI3FKqR8eos6G4vS/kM+Q4Mkt08rYeI4M0u/jplXNjScUQ96W
8qwobDcnMmGc0ZCXoCBlXpOOHVpyZEv0yNQ4wN1MufFqAEhhoe/eo1TYW0rVR03DplT1RWlPrdsa
m/VEjqRv91/hJ+fW5/taMixm/kpl+At10dfYwHWNvIXdazxL4XXKhHIDk7nvWjl15Vh6DQ4GEPb8
dqCnatAA9VpOSJGxOM19zr9AzRVQ881oBHNBqIPNsXCRWiaJ71LIZ2d0yikp41x9ffzeyCXmeMkO
Hfc6AV4rVBd0HgifrxSCH4Q4IBsk6TuSzeGYuKOvr2b5J0iWkaoaYbuFmjpeBWhAZCA3QNUSIspN
Nqai/zAo65DLIXenT1G4bef01d0aCqQhgz3gOjW81vIgienHpY9htdH/teKRgJ/zHIJVU56GU6sL
bWk38ZqosX3/P/XYSvQ8m1ABLShuruN0sa4VZphu3Ms5+9NLE+XvE891fZ0DaFIHsOFuDTEj8q4O
z/yzg/RvVXIIzF/gBgCbudQVctQAGE20fF1AS1HdFc3yqL6EZ5hQX7dhcDMECogVg/DqWgfqpqJc
GriEn2zqLJulB4DFzr5a++TKY/z88m+7SWYwPbtXsuzHAZmWo+99LMD3S9jUV3OOA7HAMWgVu5fy
2nXxX6EXrD8jIY681JbaHWAYTQb1W8RKYm5IiG+LIRNEPIQ7nPjpqcw5fqNHzTy5iIKY+7BeIyO/
qaK/Sn9WPSCI7pJXjCKWdMN4WN6PGhzA7/67/Ns0TQ+esOIEMFC30KBiIZq4JZzFxGBGz2pFSGp0
3c/zmUV6uFwSNqeZZZmcYmNJ12ij3Ay+pF3arIaliFVtIR5BdnR/bz10OnOzmWBXLb2u7Q0V1jff
mL3u779Tu3R1J9be7bTdpj9gwNJ7rg6AqvD6t8In+odlssLJUqwep/chinX2/C9JyQZA/yNtvgV1
7YuYtKmXLgy+66Fkh/pa61y+P5tsxr3j9pHT06fJE6EGBkgwuAGitNvjRZJiwWuMNqF6JfQMJS0q
W9dDJMUfkYHtF3SpOYb+bT2SWtpFsPvKtcN02CaJF/FPhib4YqD1Si3CdNMrb1IflY/Wpvu+BG6g
7tFLe9YCilWSKmr/Ct0plfkICdK/ob8IjvPC8cJs8/Duk0FnCMa4Nm52nNbfdMYCLHgFZbfaqxeY
6fTCHv3KZ9voFtKmTccFZVEBSQbJ41EEnxyYWrmxLYBntPQzQb/lG9DF0ULu7d6QRZg6X+Qqt6+c
hhnfskO+BH7tIWuoAX0OJ25RF6aDaI0dtUxMyz1xFkuCu49J3GmiRW9fRfiZWtB8GQxdLNemy3wY
dg/UhLLL604Ljr8Jna9hV0O4vCY73Jh+SWRHTUMazMzwtN9x5l798UssrjOf32CGjPnLhFBhbB2e
Ttk17RrbrD5c+leNnSb9Wc9pH2eAJ7KMRKwQD+IwErQTQnmzCRxKNRysLhmBGcxyLn9Ev+o5Jxj6
hPDJ1hK5SE7dF9tqPp4EizLD7u01tlplcbTRzriCIr/vlqgUt9HL3rhHJ4YLTDHFd6Z3vZiojD17
3FJntTu99OTprdMW7tr3i3XEhI0P1Cmkk8EiBEQgEhBSlTVd2K2lRzsJkytMLVrnO7NZH4YfHmSY
Iq8o9JxczSnDSXBlie0AhIlsHZt9W6hPRrLAn69qaI2alhwzW0ojASWYSA25UstDUOLif4F90Vfm
7V9Ok178WznLmjoEV5PDSGTR/8fRrBvQtoVPEt4OPn+C/mgkK78EzxeLQnK+EyOUfAkQzzBcJMct
QF7cQpWXNbR8WcXomAC6vOQvXzPmYHyQF//o5dbjWr0rlELN0ZjHrTE/vohx0029zySvhWb0Xvho
MlqA9ySchlbE0uoGYi2Et2TzLRcxjC74pBdL351UIeYEfsBy9MBBz/5TI2lv35PuYUMmNTvCPyNx
LuoMDlMfSPA6I+zLswNbbytDVFM0qGA1KBuhbvzMBm800ULBnw3fNuic36ZbXcKB01tDkfn/q0HC
KPP7w/2Mr5kgnZBnMkC+7bxhSoJjBdCGDIJUubCRv4X1Yz11ObMPFt1brX+pf8VxstdQVSnwFJVV
Lr9YKp97kOZ234LJPb08qBoFklSxN8kR0t2r/GKbN/tljUNQUKooD6WjAaYldNRAFyWsSu40mXIu
Pts70pn/cinxB7TD/QtiM7Uhn13Ygmyrr9gPU3VUWlgUP1Rl0K32EbGQToRofMt6p5jaWJKvh5v9
m3mdjHaOYv0OHBa9tATWLmFnlX5MxdQp/F6MPuhP8W2V8tFux9ZSa5teh+25sENPycOBZNJ2PBcY
QXFQ72oVXIL7PTDiP5BQLhzHFoVt3RVSGgfq7jytMc2yjOB2SwEc0GbGTGb6DckZmw3eyqjD6vXJ
cN4eoy2OcnqB0oDQrSmyvVCWkJPxse6aIdyXOtDK7loVdNzc79xwCV/+CBvlmc47WK1MN8Z8BdYM
msJoqTDQVQj+r+/qzlC03nd7lJ8aJUEncGBYl3oYsgMWlqfFYZMwV3Fyo7SV7cEigrJox3GIdheQ
cOJXg+o1UK9+maNgdZsmhBXUybUlhjOkrZ9fhUNu1z1/IKyB/5bpna57PvmnZXWgERU7YgKcH56H
klwp9XyZo+Tn0Y2KlEN/ZraO5VXa3rIIvuLXol43nDva/WGndrj7FfFLXolUnLNOXUxt8Hd6L4ol
Myg1fyMxLQtyRH4l7+Ggaa5af3qk8aOCGxKFTgU9qRkw5SVUuJhs8NwzNsKZZpIbUnoPGjj7Ixwd
XzcMibAdZn3NeY5l+xResQBPfi2jRdsCYfC6TmNzdmQeMtLnwEmnJnGsvfrU7lyZhhsmKzfYgiob
gieZ1PwNHsuGaYVxL6N8SluNqP8vng1C3H6n5GV//acR9wxuj24Woh8yaM96IrBUwIhlGgqZ9LyF
U+Qr6mDx9DHLUK03JfP41h6HiRFD6u3ORHRHQv8ZQApRT49j0rDBZ04zdjxYEe1hwFoMTZM2myGG
dNW0DChLTiSIE2r82nY8lOdYa5YDfrZ8zTJ7YQF1SZhM1yE7bE1jGDCUafBehg01SrMoyydS3kWT
Q3qhpiOtUnza+atGW5dzb3Mor77mJINMmQUSyljCnGShfNOcCksWEfblD5/Q8erteFad+rWrn2L+
ZYe/MMUahq58SOXbmc0oHksd1tsNyKlnEjZ3BgM3mdps9JDx4KCT7mugPTfte+66hJvCPkfSJZs8
tzmnyez969dDoKbK11nGKLKllhg1gYm0eCdW19Z0Pr7DVNGH9FGqLJQLn9TfmZzCC2p1+qPub8pj
8x/1h8gln4XUoCiI64ItKVtdu40RqaoTGvhCOSuipS8SqHClkfEtxaao/3pXjTEy9Wup7g9gKord
BEFxUtqxDYVuxegVbg2ngCFpcwrhE0+v0BKl1gE1R6SFdiMxTFe8Ea0Ofspe9oHVlp9hNmfjUVnq
5WS5YBm6yhgsV2ROFUA+43sOPuOSslUiD66T6ttcjTA1mRVscjx7Rw/LoOhE2T70yQCSr0MVoReN
yJH4KeakqJmfI5+/glsYNshrVKsnRiuN8zMoUqJAQ4++BkNroVc7bGwO/QN2sgIQQZL859Ev4MdU
V23A2JHJIHuG1seJkQP7wmYNpkKc/Nkdwj0HUBnCoSzkKK+eQImY5ZSMaZnJ4Gi06meMWRL9sagV
4gVVQMuxLa1EErA+BX9zL8dwp7IpuMNJ6hbGP/TocneBdzAzhDBYoxoWOnEynk/cWGgmj85xq56a
qx/OILRrcd5hPNgv+xaQuMpXgxT9bcVMSlyTXT7vjsIQ1si9SuyYB1bgDruCVoKTrYfmdQnFrSzI
JyOaPjbKRyndTfuUdv5MFONhoEnn5KSLHuhI0XMatjndgYC6jNnyVZ8RFQxuWVU4sMOaOLqhCqPr
wBdk0U6GRG3D1XnAzLOX+LxWenJn2lW89MgQ9EwtKuqLNeXCtfwhaN9SEpotc9hS2/Efqa3f3WWl
1Hmcar5ydtfxjc8DUzRJMvmCoG7x8dNHSlNOeXf+ttwKvzHoq/BDt8eGo7fdrgVVPzxaFOjcEFRt
nmwpJbCO4Hk+6Zv4UEOMNXRbtVvJxgzH8MlvVj6+yKrfcOGmol84AnAFPp6wQNOCzdTW5fr0BTVc
nX5AnZl8eZ7VUYoh7TJmKjtXkm/CpbH0tzSxepoALCnG1wB6u/lpxndbwOI4HH21YwaPt3l4RUpL
b32vjVEAW5DUtrNp48qtnyNDfJ0Jsi4XD8paD7pPZNk/vdfDdAwdCVe47e0/qzRtxnTpCrDOq3Jc
0S9ZL84Lp+8PR741s0wNFFv9NTYcNQA1cZaImpMH04OUI+cM2CUlnNca0ukxvcB2mvhH9nrBUTpB
HtbZmF2FWlQ9yElxb0n3h/gj7u4GP1Rp/1QX12hM7gou6+wcZj0tKXeLEL3leoVDGFu3Op+JCkt1
AQ3RtwvvHC0QV+hPKf6JHVWpFlfqhQ/5soQ3Ce2VwtGTvhQNSU+DufM3sw4LMWx0dJRIdonImcU4
XisKhDF/ieFSaf2Nv93iwarV+1WN1rYN2JWvRLMNuuwplRhZjvyIH8/0tjBobPYOjtMX0TtHvL38
pnxhDus9GmCHiNbiR6BE5WFoEM0thwuJM3uPMzpRZjYiiriL+zw6ZOLgCY/z4X00Ib9iQiciDqa0
G9oeFZeAKZZliQSkSYGQjoGFGSDk7jEPSmO5w2OP+tXUIWVVnhYfrSeo1opd/2BVW1ww9P5w95wn
8u9dtN5HL6wxPBG0hNEKf1UR9N4eVScPM+jMpmzCGa4sEUrYIKvaWUcNT8LSwtaYhl0jdcnZGYUt
pkWuQOACsnyncLRuX5q0tw4rsVSVqMMV8O8+5ccD0wLJvEKtRlkh9as7fX+kW8ReI8zFYNEMcArk
AJW7uFhNyiFrAW8xBz24F1upPvo9F1rzhfcYGp3/20FdcTBtFcbU30kIDbipnTAED0JmKTjJW4mg
4YYihN7Em4/jc6xJOeFKJe28WcFAVdzZWie0y9ndI4DC1dKfMFcXRgFjuu5t/LEtvrujeOgNYvSk
VRbaanh9Du0+lom2fl/7DJyMvsOWkT5KIjxForaP+/5qWDxD0DOrfUbqac2Ps/uG4diTlJH8kuoG
Pxa1XI2ETH2EvBJkZRskXowjzHV9FTZwzwFH30i7l5deJqAMgVC0rBMP+tw4mv/a2AEOHH2fro3R
9C+8s09M+0lYo2vm3zW+dkiZhi1sx5PEM0CA/jCyG9zLDAFdQCo02EXGLOrL80dHL3BwnG7v00I/
idgcmI1u0fVueltKW5UqQUH9UtB6ToF3pYnSQckxyTrd/R3sd2jgcTBLYUttKvxEIxPsa5jPk6lq
KB91bKl/1BiPNqHtOLlrtAsP7txWy5x08eL3w4ATx+gpeDQea7Nr6No+R9jz44HArMWOiqNQwom2
xdBEl7axIfQgciS+ikjxMFa7y16jTk80nlfbtiabxPVAyjW0lNf+Dtg5x+YFZJqbco7xyBXvnoGe
8FUn+3qgCFJJxF4uPMg00Hkr5k88BwZiSFKva1RxKT+YX63TXjBA52q30CN0XEpa0ZfVGH9meI/1
ei9LN48RkIEnPtwF64GfKRFofqOtbG/H1dyYwveuE/nmqxT6HxzH4viPoZri9vMrA/tewOALqjAc
ncGi+9ffCMEGHDaWhoJc/wKTCNf+Vf1LG1AJwVaa6IiiSfYarf14XziKoX1r8wxU+ZY4aSMbk11q
Tta0l0D0LP4f0qmpB0WUQd6ZXyLkD2uADsLW/vmYkhb/aQcj0kK3ox5qshnntY9tWq+UOUghL76O
hD34zX/ZmLE+xJ3eLhklXELUhZZ9QithYq8v1d45JF8aQjHmPBe1iX52KGwDpMcKUzo4rST08b/p
dXJkucOOUrUkoG0lkJFBvYmgcJzVGBUIi11iF3CvMhpIhUUC8oZJOtNbYiHYn2WTF4jzU5zcfhFw
em8Kq36apIZojx3ZH7p5+EQ0LAy5/REvCwy7+yHmr2AyvET5O4UCu9sA1anDJUorcwryVlRU0Muz
nuQNzCls9lo505RoigVS9jdsicxbEYeM7r+SxvARd1IjqLoLfoZRGHCCp6Zth0DUaMcLf9qjSSWi
EdSltG1ObwVfxpiw3xCOcbrINOaZSbCXWqtw4IA8FFxOkH9x0Wqv8yF+dN+tGRVQ4be/vDcck6Cn
3V1bLcKwFkcJ5mws/+8X06VKmms/dHMzcxtTsoJyk1+7OZMuc9SwP2lHpiXFicMJw1b3f1FXtrVm
pfTm/PiyGf50J+hE+2lF8sL3GPL5G0PhFcrHW+nYNHN0PYki4awo05kfQc+Qb+seusvzbNq/X9Jb
FKvOUUC4Jc8uLw409yz0GgGEN8UNqAGI1p1gSXW1UeXwLcUEueRBlAc3HzQxiW0vGva5028x7MmR
Pd1aExEfFGH1WeFwpLct1p3wIRVTMXNs1loI9C2K8FD48vF3b8JCH5nXIjRz9JZFVKWVVsm1oKBI
RNfOIfhOUpp1aij3HxByonH/2JOnjXOeqXQsSTiQlOCL8w+b146sCz9BoYfCDNt6gWOGgdJrXPJO
wWYh9xcrLVqMa8KWUQFkzdLqS8mkfkRSmj6E73LbB0t4bNV/Tv7B1VmNq5ZXMdT0klmGlrTS/WbD
FtrIOKNzkw4zKnJEyVQ8TK87q2TaRPhlGIUN11Zx8BsBiqgK6qKGW8WUWpuGWY3QYwWTr+qNxsg7
oAlearRlqlJk/r6Q3KAIQEoW4rTpuZYrH/45mGUcKi0HUvzjJsDDyMYEA3XeoyaCSIxECB3H9y/I
9mHeyvLlTapj+qXsGzm0io4qtG3QDVMJ8gUyTk4G5Tnhfwcwm5dXidggtpQAQX5nYkdVcRcZSdaF
2hfO9g8/r1K9Tt0DzTpiS15Enfx73fH5H4v776OxcgdJknASuN7UE+nZGVJb71Zlalfxi1adLT9j
U2U4ShQlitxQvFB4GdhHSOIbwxF2MFcCi8gDII4MB1Xn2hTPqbEzOQ5llDskrCDJ7oE2qOPPEvCm
KGRxwseLM5GbpHwcVvDOP1L0OjAFc5uM3mGLQHGBmiaZNYTOTmNvr2mgY2dGhJa5dXl8XsLhZiFV
n9k0+1tJcAYnRRoRhqogtrTNm28fnZHluiyfOQhRRVPqNKWiz/W9DCw6zbJwineJZqQ5o/GcgHtf
Engts9JgykbXJkamcGfLizho6u8IlLzIkoruNy9RwdHXcmDH6a/PfhNeHODEhu61wKUZZQiYeDD2
8ZcI2dmvt5iFmduusbdxMsEP53jJ4LXDXQvdkIbuTzzbVNSed24VL90oLdDW3lMYBTG1z2TjsXws
7yV4QVEDoWdRr5Xb6X7Hmf6KIof2mX4P3ROADdlmE41FmAZnFu1Vnl4ti5jYFTLoXFydMLBzCbcm
FvuztFyeGw0iAKMbY7LPll+obiJaq4OBv/OChbjkcimzg+DyY/s1d16cdQNDuiLArx3BmkzgePWD
Ad/v4YnG3rboHU8RpIMPqHKyuu8/4hBuesKyYk+ury8JOUz2GZWkqakkE+txyPNsEa60iPZdsnu/
qdImDJJIr4U++rkKy+TAB9EBTwXEIUAUsf1kHSUjEY2CXbwY2jI5hIKHI5dHNqxQM6BwbjoDgexL
MqAnPjsgMJ4GpxOvFzF//8WgXIcfAVSwPgcfBTGpl39vVJiMPD/rtyQCzvjcFQRBTeumMm/NDr9m
gg40QClsg+FMBrTS3xofwmuy5v+k7PjefKfg61TutdOOzLzZkjWALvOEft9g7ULGhsyx59y+yBed
zzwgoOHmyMEa9KrCP8M9J8D/YjjtMPOxYuH45WlLtmnze7OU0h+fvKncyF5cucbPBI7p9kzzHHcn
r7ZJoNLeNMEEprlic/+rRa6NaF3jCk2zoI5z+xpPtePvN9E+1UMMAKncpfd5ErEvRSOBc8sN1eaX
AWrf/IFcYCsxrWrHA7BL0Eo/J9FeGNrd5YU1q+O/x4ge2ABPw0f0feOAJ7odj1x2UjTE3Fysrm7S
RWPuyJVRRtGHfRFEkSyrVJEVx72V3eqFbHyZXplnrP7qnfCl7r1pKyv3FqmfQDJNL9mIfZgoVw7C
8GA2J3DWykUKRWMfCHTFBYwSMI6JiWG4DAABb7LPQ53fd8+y+ErGAOmvTYL70Fcg+HKuAlXJ+8Gt
S6zbqv7cTmXseiROLyDAkLjjge4YlCHw++nH7oGaHhweUK+b7CiYI/ZJqz2PmmWO9crq8r3bWG0M
r8w1gTxIPE/RtrwsNsXFNv6TqJ0vWxBdP+aKS412cTW3Am0ivvkKLSQewVWHz2zmn+WQgjPnNtAX
lDqGxJmNMW2kUCf0kvmOdvYoHvllmm6r46XFXH4K1NJzo1JGrXOnLckhcZ8hcntIek0qO58wBu5o
Z8ki7Xp7REGyuNKmIyijHVOQE5wvbafV2PUoWUx4ztkCZQYWPtDPfEuK1spu8uQd41AtMmkUx816
2wjim1uRB27VgbrA5QWiSwdEWCY1BKA/bdad2yxHysrRPDuPlUHotybEGayoRinr2n5xC8oUCzxS
31YsLpCcwV/i6BzpxbP2GrRcbqL2iJCh95E46aQkx6zIIBJNE1dfKExec/wMK1b18hNfPzGfAu87
hwv+5LzG7Jjq1MEuMiPk53V0T3j9IS4b455BpaLb86y9v0nT3pVApEN79BUW8Q0gwdBVjqedncpx
f3nrQrErGb4uBktfqqN3QTx/UAmmn9k/3lTOcU9Uib1YkztjP3y8i7SbzvcCLuVoKAqw/PpHR7bT
uSi1OvOcDkioshagmUfOhNSzqlc/9OpPFCx2NT63p5o3MbpnyzGtedaqzhpr3cB58TyoRiTuKBNm
fSmE9O1Ez7Y+VFZgw7OclZ1zCNHjV/A4ekbe2Mue8gD+ESmA+Gyb40of2VaOQq5ovZe+z2gcHaUL
X6azeMb0mCW6B1gvch/ZvxDqjms+55pdf+1RRMesBa3+uQDeU2b43yg8eZOoonDqk/R7r0t8n1kt
aMv8u7p8NAQ1WcpcoW9Shw/xv2geDuuDxECyLtVApDfwindOOtxeK/ACmw/Zv3lUt+iNTqin8KJI
y+WTrAFajIUImW+oK53/sPqGxyhc1lnZ58Dn2wSPSgBSapGZWMep9/3Fn70x6SP87FirXI5HvhPu
ShwJCn4sZXc6nDDlbdYcrybj6k2PtsR72pzWvpboGesHaJscrnprJyo/j7irppWBKdzVTbtkN6Cz
OptmylhGMeChX2+2mm2WdpL+DJqX1L5mDfiuiYguE3qTjcmMH2Lnsn5Q8gnMF5KyIZYmS1G/H5Bl
cI4PiBqVhl0UtjGPOY1i2CTSA3i8MFkBZLHLHW9z++yU3zFDJrJCuoqyRwiYRo3DUakX7tqbUU9V
asWnbauPh0j2ZmGe622Bejy+RKj2y2tbuKr4ssCWLhpevNG1UHBEp9mdz1806PsY3IhXkFrxXdN8
Oui/3eu9qloHoJx6UdWXMF+mO8tFaPi7uIVP9wKMCx/PxdxuJ3+1pOUnrwpQT7tG/DamqtcgrM7p
NeD+GZ+0mv0FzqPU3pbH/9aBz+S5Q/ehIefZPLm2l8XQ8JIFJVTcCHYakJtYAN7nxaw7XYB/Nz1s
TLEH2zfdgEF32dTwRGHuqpALFCQIpGuZgj5mArVG3OwBQe/Y1dq2rWGlNBEjdRcFaNH8Q1r4FSCW
BDTk0Qf1NtrXwI3+t0tq3DJehUOiQSSw5mq0RYYQaF0S018Wv9lLDt/XFRf0B3qy1Ct9nyH0EpAL
cbKrWBJV4fAk+8YNxZrl9k+Xwn+Uo79/VIemVIfWDY2Wh6l4TYByJfJtxGlxBkwp2nJE4qsM54Cl
sLxgQLJDkt5Wp7IBXvomW8tz34ElwUbyo0oyEbL9YwU9iZNmVRlgulDIEVZeO1qutq5b/3kAovxU
+4MG21TGqd6iL9fX6i3lVpQ/Oo7fLXyFxfGCUoPcFJbwmXRFkGcdnzatja3pOQ+/FWHypp4VzS9C
OglSDXhJqRlTEUpVy7mVhJeSbyQ2c8oP/d/lX57JJqFunDNyXjqcF/UQjnO3jmgYHzbl7t/Irezr
l9aJLD+gi3HiGWrs/2zAeuAUqZ1vLRr/ERNPJ7Vykm/hw1pke5K662LOo1TggQhjsdOb8cEJ3LTp
jiY1EiSjEt3k1FTCdFgEWXhsjxB7SAwF+RMbPqOSifXXdCKlEGfQPmVKmkEvdSLy6kK5+BD5o42W
QS6IIU0L0aDm/bi98x8kqDgO9CmxGbhpMrZIfDpbsLdlS8zKP4bPfV7ma6QA6LHr7JRecXld4v80
0K745tXbMRUxIVuj0NC9nZD3/k3foGWC+biIuCUByOTlPDN1V51RhZaNbFXM4zDF41dtSBlf57d9
WIqq6XiN8mei0gbDqW9zNEk4kRMH6zlDpAfH3CYHDMaNpkHGMElyEO+frkeUX+xrbQxi07TFVtZF
TluUI6toHbVFH286cTIo1hhyHoWH7QdxbH3MKW4LfbaPhehUQ4HCw3vr45lI4ZTQmuS156h62NnG
ttESVRKTlEwrxmxUCx0lYOleS6wRkAaBgnNGhz6z+9FxU/4TCmsb36Ebm46YDpkHsdsGy4z9BTqM
3YWw2CPcrhJV4VV0wFtsJ4WWdpP1Thht5UNMr39GyPpKPRoKzmgVOuKxxeNHusKIHQ/Wg2V368Mp
SNyU5lisO3H8Z+A3dES7RlXplYvqjBs3u9RAlrHK8pSU6anwsP3yplQ05+N1VkjbVP4KCns5S5WY
MyAw2Dt7GtPIjK7lrCmzvaB27KzTg7O7aL2VCRMIbwY7OZ9bMgMKf8R8jviFGsTTGlPvbTwgkri7
SpLUaKHkQ8SQBXcmBeIYpvFq9ats/OigkXabHJOXHZHNeRauJMeGFtsB07NdvW1wM2uMjBJK85eF
3MPE7fql5WX5wIkt0Qx0kiQvq/Lkyt5emZEpW4GvxHaHdOUSdEryV4FamT5qaUAgFejC+fFnQPv4
g2kkB/8mVRtpZlIk2gim3FcVgVBGINdBNBBlVKy3p+bared4iczR6sVLMHIpxorRNDPl0uLbHyRC
80d19rRfrqmlzuAml3ZuGHW3+DQhRk+d4Z/+7CkwFZo6C73i2YAZesWqZbqitZllD99zsVzMniQg
hbr0y210gHijQCLzD/PMpLky4ZrDqxdtj1zIRMeSSHuBYZZAnAPxX7rkTaGKF3Ajh8HAPh/Q/nZi
ns8UINrZexxV+otmblZCOQBvLFniU+IpMnY9qMmcfCqAbB6V70T9iFzIF+OYXDAbBJGAzF/1bX/i
VLNHA9QTbWaqcYsZ6JGXBT94m/Y3wEgKdNVJCUEmbxz1j6w8sYFWjsrFlwVjN5tsgRLMA3WGszlB
s3XV0va7haynGSxgyb0TLp+8QvUCfK/TGgbKY0g4wXbA8UFOSUVULndUsP26cGyg/x2hx+HEjWzg
r6VLpJK41jwfWyYXeXDNYoxJCHSYAiKef0lTPcSs3/R8dObLeIPn1EEu/rcKYoyOtJ5q0L9FtAL0
WARMgDr0Xp8SbsS7aPuFmcqADwaMiWVhYbHoOyxHbgp5qfaqtxENRsagaeyWqcUC/KE4QZhZPtNa
9+Yo+0crQQh7pFFsssuGjwXvCoaTe1pII5hSUaMBXsJGD6g3HxouyYilW6UGw67M4B4o/0w59K10
d4uswQvmJvLizyYSCbN8ZKLpq70OjxDZEHq6OSzXRnuv3EVjtK/LqIVQQBBbgKDuxAoa/vrs9lfI
BTD9b33gL6EyoQKWh8AuVSZNv0BHumIgGYGxHOm+vsBviZO7I/xlmSBaHzDEaav048lRK23YZ6j2
N9drK959N1Y0/2z7Ax8MZS5nk38/uubqHT4W/N5eXY3989yRV/i0vPkBD6ISQsnr3wRkiqDKLr9f
vbPpwcyyVtZBY8yRp9SWQcQt9ggfF72fTXGK2cbYzFPvL43Aek5aI83FR0gRxrzWGV+ch/erCM4S
6FdPzM3G2lGFV3Aickb/Hko9EByQ4wrVAifMyfB8aKKSWPP/aL74FGXGTUOO3GDCVlrNTB/he+1+
vVY33KoWxSC+XZxbAN3eJnHJo/qu40K/pXa9M5IEoYuUR6gtAQvSew/AMOlg2DAnDOhZq2HifrIu
Sc0I+7RtXf7z6cM+1oChLDMV0GBd/vgUT22ezxIW+3eE2O3NeoIu5cKXdn32xGWQw/evk6lv8837
4A+wlHD+M8WrQspPndV0i0xTS9h6SEpwpBVNurh90QIQeQu9lUbTMdhGPd4mdZZxYplqbKZJ5WWF
OjUJLtkF44BdYSgnXhi1aXh8q3wwfh7j4lWv+KXcdQoAn3AxCXz4ZBqRvpzKPDV+YlBFCAgggu3B
SkLA1rmnSDTBxe66se24Cvvrdv9AKLUZ92F9UutXOjGHpDjHmvVy+jebMmvkQCpwxeXVVvKIeTkX
OjvM6ePmPV6MfLR6Q4NeyH2LNttUSGwZ+Wzx8+xEm42mamlXekQV/36ofl+Ekf5rka8r9lOKKUPW
Lc6e8TzA3rKRU9GfaExNqcvIwcAflUgQ8FEW07BJKwRNODfFqiGZbkMRaMSPBwUfVytCra70crib
K1jWsIaFTFrGPKlyk68nz4QvxvTYhtSd+stETtY0HUS6qqd6bDDAyvgeMX6AUh55N5BmR0wwsmkS
TcNTxRgayEM9LMrk5VuWmyUYdM0qgbFrmYEe/XPOukf+/aV2tKRl/RuFpP/jyojZdFIKPXP1UJ8O
in3SHTPLPx/5OMb7DDkjUJKcPWVNe5v/kxEGNXcYxwNAC3uF+HPXpub34rE1FdiKKStYnw7CA9Om
G8hyfuNMGKUTx7ny4iXHoV1l6AngPuNQVOhdSNChzKehwtl5zJyal4FLN0wfhTI4WEhG4+P+nryu
A8QQ6M41dVt0PMMATtF7EIU59SMYlnh3VMRiFKPCfQpzR74PtkPr4c6AuzY1YXxOCOVGgI6c0zia
+9Gd4EpxTfWu7tSyolF98+T2Gd7K6Y0gIBTW9NJnnmEvo6IiCHPJRKG8c7OA+o7rmRxtJhJihwZx
Sq3yOVu0PnQzj70O5XMjMyMTB6nbHP/R1jJmD7g+xcK+/suYWq7ZuRhFStCzbpQ3T+qnzdrJz/Eu
fHNKem0ory9wrScA9DTP6qAySVx8dtTlAjNUS+ks09iF/4ZyiEUIJFtYNHik7cXxpdOmpWo4FlMk
q6zQaeK+Y+ilJ2v9EtzRGuw6C1e6RlBw62yGgryUMoTgB9Ej00Kgk+VQ3FZ1o5Nw8gZtrHnTZm3W
U1BZ/uifJ24FaWSMpxkarY3cjlMj52hYzrodkl+O/1ZMjjgyKrxSTzzC5Yy+vs0Sikep5g0zxmXP
j2oGXgffBJsCKHqlee1nn9M3TkThSLQbJKbaMavuEX7QJsFBPfn5IeJJKyxJ0pzFAvFdDOKxamEb
wuf6iEqKlAdkJutQQA+WbHK9+6fUV7LnARlFx7EIJEQmn9SqshIyE90dwQ7twpdDV98839hZcVqH
QpWkAuRatB7IMiaXHkdjjiBzPnr19Jb78qS7t7aiO6Xa7ibwC3bOHU8VeIDDjWOlJDv52vmstAzJ
Q8hR88Et2t+ZYENQqH2rpyqUTjOkz01oL0W5NJF2da+h4dUVNKLH8d+BOb6V2rxi5sGHqr2UKC5c
0QTeKzHcsVVALxxXvaEzfM8MFtKiWv/nyQj2+rqU4h7qAl+2Bp2jkgDI4UQJw60+EJ4wqGhO65Pc
tE2vUJTWZcATYJhVo0RXAzFsDAG4SPuXrLxJUFvGB0WsgSMh1Ba94zB0BSAXHNfFdEqr/aL3cnrn
rISarltSunDF0UNABFDs4NQ1jaFmibKvK2GfncjQFsGzMcoouwkCns8LErWwO1v6FNsYl6b8aGMA
Ixd8POUP+LCBHk3VFpiax8zBYEMsb8IGaMo7vmmaP74gyhH3mcVqdpspUTjuFxPDGB2ZB5fW+oX2
tjJm6hwooyxgvcg7ssDrIFrUTNolBrXT9FluMaQO0OH3OCY4APCi9QoEZHNVZSwOgy7qbDHdXIgw
dqFPbKpt7Er320ZbXnROn2OH94TjI5nrJc8kP9vSROC5TxSKrSYS4StVnB5X2fBpQkgOesEJ2K90
oyVfMdeGeSkva1lxlcC2Kfs3Y8k0W0c3o0WEw4mHmwliFeYE2lIgU/pa/UTm+JcjdD4kBuHwVs8C
4VqN7EzJ1dLkirL1jPTZy3cuhiwedPWka27CRZKH2JOVNtce5kbKSTRcGDMEIFrhrdhw2S1y0AZy
P+iz/Mk1yUw5NCyix9Z2JAqKvm/wWEn12JpB2QSE+gFMktk73a2lOYVocHzjzEhz47GJ4XTgLidj
Lgo20DYDjikeMWPMEpYlqM9KseXMOJ1LPKKUunkRLqWzj5PMbNqny16XYPW+7bFlVM/vhrL3H5rZ
dF9gtVOn88UowEzh0gAcO0y+yjq5xJnta+/i09fjy+W4PfIQPM7LYYIZOiiW0/9YtwCv/JN+yUTp
fm5Ytp/BiT0MYckGLUQvjTnj3aDPkvSbK6KygcTKZgq2SwacNmVqEsLmIHINdGDg8waUABa+aD7J
fwyZ+DWOcxhDOVfwHRn8nvJBoyOiitOIsGERiY0i0PdZSfHfU8ckk8h7FSnJJo8hXG4Fc9U2zgk5
zX1nFfvB6ntIypyP/fRqZuR0MfFO4SvQxlZ1IvwYV86jnPhx349AZXcWfJTbmuLAEORniyve2rCF
m2I85mCdrjl70/tofsmGNTCw1by1tQloJyT3E4RHNBxWJeSQJoOkSJOQ0tC4ktb8U/FcC8suXkTp
+rndkC5rDEy01adgd8ppKoEQ6oLGMLlgVqi+Ds3s3LdyUnUvg2UaksMUPm95w4eamPgZgq6lWBci
p5haFViiOfL3id96czJ5KQyx8/iEbvOu+gxw8fiGU1dxuOul2+pvvQfXKCJ/lC97TOCDRlsYT8DX
+EM2xTAn1ST/1WSrFmhdKvHnK/B22Vbj43hejXZntTGZ9kwCEMoyhKiLJmuaUF8VYCth6skeawmz
dKfiPd1McXoFLav8VP48O8urZsT1dBjcZatRPwnncMcaRlY9qbq7xC1mvlJOIbiPkqNnUXecGosw
ROh9P0Wks8znlx6omlJCMGXKURMEjeYBx7PNgSy7apZiuwNs9qT9x7B6KJ/shSJdCmkF0YFJYCVx
/EynLNso+M0UhhRT3YGLHmNWavjUGWrOdV1RK99SzHmpDixNuDedIlB/Dt4w776ihnlRsTisHyCg
n1ILyom+vKlcHUJ4z3LX43yJYzvkyNPFT1EUiTbkE/1YLg3HoNaO/cYojDy63M+jI46pDZJSNxCC
GYn6DhPSSY08psLYj/4eNjJYdEkSCuvmx5IRFOmq1Cf7sUwoWV1I5S6XeIgJtDyCYKluOslO+G8P
N68qaP90sD0tCb67w9iKPZZb9QQ/to5OGp1oVqbdXTNMzbriCh1Uuy2nCy8AykcR45KogDoAHcvk
Pquo9EuGAW1UMR6LnCzlI3N3XLnVYKVpu5sw3OB5oqRBKIFG02mX9VIO1G1jZ6i9JB9q2J192AXz
ysvhUQzLF9nfsDwtjcaetYJ3/oY2DHbHIc5hn1Q55pVUJuZqoTH81tyUvTH006W+SvdnvNT3GuDC
241Yj6LYqgg2WpUXAm1uAHbi/r9yS3sznwVnljOzIIQifjFCBdG+pK3yMqebfvnWtn2F8KmUPqWN
KWBrCCSEIbLG85wFOZPXytcXDU4HbqVgtL2bKYP+2pRCxmhQBwV7KazC58gx5snSx9pUD1kdr6Ma
C/L3m7zDsz66SViiTQhqO8Dv1TdMHw19MC4PEJDjQGB8Y8SWZX9S2AtVkPVXtFBsyGidmYlPRPAe
v1dIhheLNPQo9m0tCDmS+bdIgEFs2Ce6NLCSlSllZifwjy6r8UEQwIHx1Dpq2mgZrZFT+oPDNin5
WDydiwJhSi0JHvD3NjVm4m1hzYxFYTRXql3tOPoEQZpoAC3Xxqmc0i1otu/6dg27kg9mpWOtiJgE
ZRcRjgwCTTn6vQ4CMc19jHEyX/vuQuTh8YZxhYsRGh8ut5Zpyy+E6qA3vHKFjauyVgDiqpXln/ej
m7EYPUeDR8hf9vNoTvj3DG6LGwbbI7b6VnLSYu+ZlS7SwKoed0BtoqmNAsKLKS+OrOPZRK5XgqVv
mMBbp6sdtqNcalrDVLWCYnfSY0zXP4k2VUDPlDtXyV5hJ+Hd6sTS4z4zguCvrnc696Cf/rFkoigo
tbA1rAod2wRkfccPmDmcm0cQCc7JTZNwGfIk7dtk6aWguibOTeeN0Opvk3/FJULaBck4Fvoeh6Tw
lsmNQXEJ3CQTvXRXkCgGDtOdI/wei61QADPf8lF7BKZOuZe7XeWAw8zETj4B8oPvnlrlcZqnId+f
RFfkuC4Ob4x+i/sndzMasflzifJczRa1rfhj/SHRXbZ0rChKJY8ay6J8k+he5Pd90WDNllL0ZyCS
iYexWQDUr/slU01Zg8LRt7bLWybrNenTaJjVUYIQC6OapPhNBWXp1j74NDHb1BjuRS89iF07+bz6
iXNtMcuxJ4QFPzElyElyMAvg/0wCBaEW5wjjzGdr1blJmi0clLEc2IyL7TNj4kHvNlash/bF3CWB
ENN0rRseRjfaORERT+zgFd8tRIUkhG2/k7X/JZXIvNLusmLsLaaKYp7KLbnn69V3kf0NvPAars3M
cqc48RZXGdh90yE1+pHFrrXru3ag9OWcS+uxe+1eJugMWrzOgSep5i1GJs6imOy9y5OB/8SjTIIL
q4BrUqnKfCUwQnfR9DDLKnH5WaWO1hzgpddPr6aLKjcEdfX9QKu1atS1DowpNJkhaOQAx751cOH4
FvlQN7rij/yjfrqoQ5f5liwGneg5R5AsxeoJHrXZrKA27GWOPDGROOx+94jTzrT2f38jSag6k504
95jjAnCpDIjY5W+WiWfTobMbh+YOqxGpq+oNQLZ+AGFTgm74lJCfRJkI8CWVbQ8J5Vb438ab1R2J
vgS+0JQos45GiuxCKiWe09dOgJSWe1hRtJI3KZtFotTPnvVMQkKNXZN7GJTo0qQYUH0ZiYmVI8gN
I2vsbjKr6lH5sETb+F0gxZ1Wd5hOCEcja3ctw/i8CIHYcnskPxC4UWcnpK5DRFNE8W8yZrLCYtP4
XBgnAXoBoIUhugSyBvqhNA1uViakIQCQDwL+BoSYopZv063w6+Tt8w3y8Ukdo8R/Q0aMRoJv2dPg
Y1FtvrQkIiWw1rofnrwt+2MAUJma8rTzYJbOYpbsY21qVZ7pS2FKWgX3oqLRIk8117YgF24lv9Kk
7LVK9hiiAynSQjyqcss8foIN6vbIRTgrnSSpfNgUId7T1bn+Vt4JbJBY7tD3MzVzHqCJ8c1Ho/jO
3Q0eaz1w2QCGmTVbU3zI0Q+IBlSIJdKfAYHBwFTMLUuBOpj5mC+IVCcMZuo65DRpg4fiC58uPchE
TLdzj3M8fesB/CjOMzkdU1O+G16ko8Fw+11XLMDCdEDnnMllsj/TwZtH4cUbwDy7FJz1XuecYEa+
8v23EJt8AJl5ZT3hcM0ZsNfPKa5eyLr+6ZTjxoJGeFbeOZz8y34woSEeb6CfEyMRCIEVYzsY4S7p
AgmxSOfY5ThVgAxbYq0EDc5BraSZjqx2pcLoKeOzCSlrYNbU0/wtsh/khA9Caqc621fKotkHikZ9
5qQqG5bhIACxzvssILfkz40wPXRc4mHk+ZYZowPhWGnw/dMpirTZ6/e78/T1WOOTJNaqs/6bZ3bX
VTrsuH19qKaSAZbUFxfsekZABc5DkdVBFT/dMDIL3fIXqWoqZuBi5IdguhoAOAxH/URud52pPE2Q
Cqwp+dzskYsdmZ7W25xL7ALDITAT4f/Pdn9FSQLwv4atPEiWbZv19L89tHN7NtmnLZU9m0cSLpVQ
RnOrv2PYn7Ny2KHWBtNCU+n7ZvqjA9C4LMVxkW8vBLESndUg2vWuKKIK3HswKGsl9eWPLrqrl/bV
IrCo0L7+gnRg89n1X4x81ySc32ipkN3CBjfNsPGvQW4Ypz18AUAiWhIKQF2uhCJuZqfbWrCk9gQ3
rbHeaHtP0HE1OS27nJZMtNCGwwZJTAWeCY9MyRBi/s/5rnXoTuDQRzUXWDtZXZ9FaDq/J922Uekh
zvBka5IT5lDlduSCfHLbu/vmf8IMeJfKF+x0FrdYCxWPtbAc6pJooFYOVjq+Hnwobvmng1VVXA4I
c+XgSVbKLjPdgc1BBPtRgeutKM/M7IbgXzJ5jcQLqMKvdTS5Hz6Uy/YHrdoK8f8/0O84zjcqj1Fc
vkR7ILNVpp1KhZjI1Mw4uCozD8lMV4hPgbPZIo20R8X20Q4P5U5nQUz2UvhEbsv5OfWMohu+00wN
RuRSF+Ov0GZOiz0LgrIPSPbWvR6mygUL1/ft4zXaScXbIlZTHLRncXRlFaieDNMhp/Z96AiJhuGf
eVoCCrKe6+WILPad7MPX/Nnv/e9Oj9YZrGbwdNN5v+/V9+59Zc0PmcBmB2rJs+Mi+u/5USxYMFlL
6FtgEwgjWmnEIcCxRJ6HEazmb4agaLhruExdv/fWbTTX+KUPHuU224zU4MePex+Ays1VjEKUyphP
fEX5ldUXFfm+ZOWCfEetJvUyD9dxgvU9tAAyC03CmRIcw9Aro40hAtcOx3PbFLSX2K1e66Hv6kDV
paECw5n0pdQ6zRy+D7TEDMrv/djSBwnO00J1Av5X/atU5IJwpGPr39VHQJJUkq1QX5pi8NrzdixG
f+jy1ew9v0VXQytgWhRYBMB4cYkITZJliLbRglBlEsi+ettWaQdfKrDtbFcCRzZSQvCJrdvk63eX
pfeJ28YIrOpZjCpHSsoMq7/NAmJoDM19/ViiK3ZuDiNFaVGcJUmKJJxcZaxh2HLjoiqDJsjxAjLO
UuarYsYmq/6/eM7OGE6jZR/Be29jSWVlN0scgwrvcWaW6KkFRzXZB0aSSaqfvOLFPEXpxRr/aIb/
nB735tjIm5ZT2B3GvknzNluaCNnmFHgydMg55c5S1XPtdwC7yclysdy9CsHqZXhawR1vb7F1CRE8
whkak+xmPDegHKDDg9er48NTVGTCf5zxrbjVqI0uFDDWKEeOAz9PhhuHn6V8yQqxoE+ycqIANUIf
f5ygcp2VOz1NC/FSO8UFUsFyel26e4s1bOmh9OU6jj1HASauZc6PYbbUr9XQhnMvcY9lDRZO4X0I
G4ZvT2e+49zPSoXdNxyltxdSuPhr8JM1ll7HVrkRyZc2x/3+9q2+8VHoaL/8FeIJHlgNMb5c8OiT
3Vi/Pvda2PBBBFaod0OgqjoDNbbTfxIYUvHWTm/nC7Nche7lIX4q7jw/wnItUqhp2aYMp5Z1V/lL
txDNlfjuyvIwVI9Hd63qp/yvNdjzsYTOXUE2qc6CBmOAn3EurSYIb095rwfmYUA7r9MB7gLZaLQb
wVQHs7esQcJjnsdDteh+cfqhye+rcPLBe2JMmnxQfUXB9ukcJFwm0r4NdLHOp56yJSJQqOpuIu+k
ob/+5SVjZU8PW15mhWWpZMyhxsdYWYrOQGIw4lN5MyjXa20C/+1moBE5aPH3szL1AaoaEIKVdc4A
KNyPefVPG35yDOPwnFrrIilOAoXvYP1YIQtkal90pZxypHH5CGdrDNPYJ/uORdVSm/ETmpcwOGP6
Mg5VohKpDhRImoPg+LYRp5+QL+V3PSfsI9/3lMY1b2yElliNc0Eq76xBIz7N2s4IVgVwwyPF2jId
LkfVJ5MsOxkzij7ANhaWQKpOvQEg3uqejDzbHuEVWCTmZowEgxUDLMXrNBFFO2YQvMiA3fF5OoAa
dEQuxloVjFhtqKBMzK6SaLCCOXvqQzV2hOUlalhedYT7E/8IRJAXF4cJeS/drMrFejXe2RFoRaby
Ds+9p3c8lddxd7e9MdW6nGhYU+cG8RwqYQ5F1AFjzqE38HrNLB0/XsPc8RMPi55n75E9D6GczyiD
aNEOSX3KjvTmKTA9jXZ63Ge49s5GXZS2hrOOrdRsYXJX53Jgawkv3HcW7SHErBGrZJHgIreNlRca
ADMpBQMFknghTp8XyOVrpU+/Ls+reyvqj8qVqzTwgVAvXdqlQvGB7VkUlF+b5cmerovR3P+XcZSH
ExZY3Oj/kxmCzBEn/fOrD8qTGpBlB4sbS8EBfXfMfYcmRJHf5LINve2MINPet0R9LGVZnGIn9vl0
/+QAbeuvzyysCm/VAHQ9WmQcEg78lYf3Np7cUQfyO085jqgDRSbY44n2EKHq9zcDCXp3Ic5l+Vz7
VVui9S1P0SC8DkW9O4/VK3FydNKBakwAtGh/fWaeze0qISn/9jDxm+dtnBMJPf3aFRh80meOTb3N
fDJUIFU2XYNo6E7jhVuaPUWuw+LgJZVIsmCTW5kLqqBPeo8zGyE9GgQN/sotzbWgtakouWwT5Cag
ELNz9RbxufucTYat3pZ05VP2SVgEkR6acCVIg5Nk1oLwuesR5LqmHyb67Cn0xVT/pgJqD0KbVn8Y
1gTmgUdA0OZ9Z+oMkuQvqNuYgAfND5bxPonpmeTaZwIfW+0ZG8k2TxOvc7xVxBao+xtDEiG08Geb
Z9UODD4WpBiJCT25jQhegO+khxSfhQHxquKjBsR7q8YXVcwEBbdZWaaBVfU+x08D5chWXDsqYE5O
PqUJ4RAgueQBwW373+WknA1v80ZbuUxlBDpWv1ZK/I92Qvpr1DMkZ30/XNmZ3nK9qblFNhEySSHW
7llndwXQySMsPdOPGZuzotcjGUfEYPK2SxyPtsUhNKMMOpOEuENh6o/Rfy+v0xOgb1iSNHsBS/nS
qvT2SUFIkZdQWR3vW8jefohT8FA1wQ/R9COQCFS5bXJQnAzKsr62V8lM40wn4w5vRZsWvcmk79qG
QJ4OtRUZ/LV2Mhv8mlCUixZlXTNV8ljIUxrii31R/n5kCQG1D418Soe7H/2ndK3cZYE1hwEiXJ4x
zNV9lRn35NifsfLNZKxfH1Rqf0yO/HarZWMiCv+GzDAyauvm7JZ2IY/mixSSYbNY0NtbYqXboHaB
m7jKjN+UAOLeBoK4B0dWxis1vMnu8HwB/b1O1nMF5krL3pYNMVTKuSDx8Q0H0eoM/YuiF68yhxCd
jPSIe2eYGQcubJ+qFk5652MQpnmRncZScQkM0WpLUkwejJgg/AdbtZ/xRn4ZvxLuInGylnezRixh
8kTHHkdQMpmFfuKWxeHelG6DyboBRiylt4pXaYWo5vwKcMlNyoUrWtZSddIR+STBP8LYojiFXMCM
9THDRiOPNY7k4lVMwv7HolUt3RmMducMlZ66WA9Dd4nJSkoZNG7M0p1hFruY+JsRcOCtbGx+L/Lu
E3MSuysy4RaYH1Cj9uHSEqdiOdRtS4fDCpH5b1N8usahN5sY40X6H2dqcnJvXYEjFy/pk0y8fnoH
Ei3fCEhI6XU9WNQn9WfZYWFfnnBdItVqHxLKT3U6bsLHQ/04TdQnX/RVxoK2ViLp4WpIhwhFH3al
qlIQkPEX6g7vfyDghJP1yQKdY8NP7dgHG0MTm8DvMUuCfjFnRlcsWDP0Nu9P3d+ggYqOOvJkPUPY
trfLoAtSqPtab6Z6Aio/XOdgkMAgDBQFFOyOZF2S/J/rWXedIy1k/gRBOwibzZnXLQWUvvAz/vBp
Dc+jXgFsfKhY+JlHkSyO/4uWHQNGUiqXZ9jM6b6HUrFQAtCkorVYDSyvmU7uAKopOrWBIFADtYwb
7r+uYgx2zBpIqU0xL5SnL6+DsW1cpEPAAmrgkX6Fgh4qdN15k4M6+nA8m8iJ21YicgcLwHpkK05k
soAGobCuJVeZcAx9X8zQfiVmhKZ0IRHUIVrw5tMdAN0Nr7SbWDpGRCwB3JcpWPjcEfoDwg95qLJY
v5p5aItu4N8miIHI+a4yPK1WaB3pqR45+YTe3telpQGK8wQ9l1QKoGoKXOuhOUTpCbaXSofqDd/J
ixK6TIIVwjCSnG7GFObpMutA4r1Jekki2x6ZTJI1CI/1QxJ1hyxIVsoBLLcUiiF7DHbHG/QYFABG
+Oyr1drY7N5zfp+2X77bZUCqpk2iFibtW9eXqRjltfYhGEe2rpLxq/ajPsfQAhmGLOJMBfOyL6n3
ZMkdytGjJdO0ul/noeYl1Wnb/Ikpo+Q78ElZdyF8rEDs2SpGvYpTRe6iytfMVpoTdDE1pAEm+0pG
Q6peldeq8dIKwuiVMomFBcHrGRmDDe5DRscsRiI+LiMvI7CkW383nwtNDppvHKKsdFASwAdgk5gj
UxCP3b7FuoJgOCp8zZ4gpr6+WxZAOHCTmPPo9Zs8HhfPPgPupkNtt4LaZwwr8VjDKCaUrcpWXwR0
XlC/Y+oeFunn2g6/DsgImZJbhPHLJH9tu3QQGlEcSikH0h2PfPNqqok50u3OJ5N8CiQ2Z/VXODdV
YV4VQYSiGQd3eC29WLm2BtvTFK2YbswdhffuUoJOHqSxrCczls1AWzYDujbj/KdtemQ6hVzMlQdh
aOHqh3fyGvqAngOSq2e4qktYVQ/o6rURT1wD9HGmw19rC5feblAlxqaGrJ/8g59vg8qtQm2Tn0jo
6+P31TNVHQE9XazqL81dbV5vV/NJfSgtmYy4lELyV2iOXgKg+Mrn21GBrhxHp/1A2IUf5qvf76yR
DPfeMU6eobyGeitDhPB2NXJDJjhN6DyMclHrSMEOirZnhneRKL+cbmFveCz02JGwj/7rlJSPQ2V7
2wjdv0zTklspe6Rs737StnFtdquWbnjESOAu2v/R+6C96SwDXA/LGnfE6QOaR37cHpfrZq/kk0f3
Rcj6h8rIS9koK9gLDTAFy8JE0HfCKC5C1caJWpFaDkheT77vCuzw0I3gy51/dztG8KYYc38IGXa8
UtNyo0lNskNbxk3icmTD4roY3cYjY6pc4n0XdgL7wn8jmmhJznbvg99d7nH3xmiv8Snvy7WaRRon
dDNJGEUHjJyFlK/vnn5GaS3YzYwN/acUqdiraEib1/BqjHfQiyiOvps1OFTjpSPnoAoH/AJy4AeE
ZWRJExxL4xQKT0i2XqdqOPBj1kEW8qjh7IOidjHHw5vlgMV7ly1QStjkxXAqJUFGkmqOpveO1sjk
4jQauDQVmqjoLphl16F8tnmW71aMFfEgDfhktHbWPJ77O8eaFb9ZDPX5zBZ38dHo+WPE+Nb370QS
i6BbjbFkn3kYZRYvVLwTa1cO+0ixVbDv1uaRQ8tvu9kUL07aGOs79dAjNuetpn7VoiCKImDkCeRd
773UzYnLqjxEDQQTz+Z/UxaudRrXQx0TGpuNQ0tp/8fV4SuErodNgBDggS7dL/BwC3y1eeRxzUl+
SZPHQmQ8YMFremIpPPoGzWNXcJQCDz9b8bt0QpC23LJJRFglI1EXzEPegbh+POhh1i9AN8FjexdT
R/I63rX/Ywe5eV0T6dDtkwO+HXsqdFUDi7+u/dR7JNJAIO/jfqN1cMMOCs13/XIXIAEF82tp/9qL
2Kt5Omm3lFHqmoRqckFVAhGjX/Zx/YfpHMslHebOPJwuRBEQQeXhmZWM2IuPMy4HRR3iJAy2WbnI
9UdCrPYphPcRVuKFlHhe5AlWSYN52iKxWRNBJ3rkzdysYijbbM5NsPNVwLZ1j6Z8i886P3rZKRKI
r04vgHOCaMdV+LSQoi05fOol0UWAXweUhpSDcJkU3lZEtzxTIcq8351PHKDAWA9c8rCzH637nh0F
yib0ch3mR5FirVOdOoULqC2pLoaN4CQWRlU3lD0/lZTCd5gwSKGx2fI0LnXw2MDLjaE7ZLDEZVNn
G1dFOsjUBuSmHLxK1aYGcJJoYG/32kZpaEFICe5lsaeQDvRXJFT8UB04Y2R3zQDATgr/f+n8XaC2
vobjpIbqwtuMz2MrYI9fbklJY4vu6gVElMLTZpFKL2nMQAgpo/n4PylBnH4FZ8c+QJDKyr2vsbDT
q4ZdlmAAm0LbRpp9lx7tO4NReIwQ350Q/YrPeXgwZZXpFzNDb0Ybzcb/zeZELZ0UK6dR4s9qkip6
qlP6Jl4qkrZjcYh0Z/pARo2tMRyEw8zk0yS6nNc8L2TJg985RvwrYwWIT06nydj/PrXmTG8G7BWf
A7Bu9sW/Nl0nC+VKjSkL57qhb/8Xc85oCf0RFxKOs96px+/v7ta/veWRF3BbyzPDIyK3ZqpHqf9U
OvFBhqsFrdmdcCARnkTeQ+bydP07YLTc70EKg+pspArmIDyWw0VSulofeYI4IZh49fNNixt5n1Uj
NqSgbFp/gY7vSyGfkRZuoZGxINboXcDWB2nfq5aVOTK/z475gdLULS4zy8cyb0UIogcvZVofLlm8
+JBqrw/9aEaAx9YA6cxsYO5hZY7BxSvTQ2otxnUpCUjvX0knn4syaB08QRaMD0hW3k1eUxwXOGIU
XGXPLn/rSJTc6h8THaZn4YqLiKSjDeKhRQY2hb9rxguD2VMT3XJ41VUOtdoANX6LuLoRCEUG1Ene
HhDVyzoIPt1SfmT1rxvuxtdjQyjxHNiLvTePXVl7WpBSveWy7kej2Q0Ss0bkaCvqS1Uq4IRt2hWc
xaMiNBEZSAkj+GEqNzL99v8SCZuxRZuItd/pwBlrbJ29PZZGKX6PnyI0DuAwcchHu6wZWgDovdkn
kQo/DRZOgfEm4kFiVvW0yrbWvKpCc5oqXfewxnOiEE89LF9k4TJ+o/jjtKvUHGLX1YV1Ll9rwfSE
F9UdA1bJciMiXxnbcZ+vJxNZL+sLjOBsG3kmMHqZKSvxU29oFkJAknV33ggH1QKlZmVFd/GimfAy
XwGosIbLoHy+F8qbB3s/mKqtaGYQQt+47nIia0iYl71fKQyOLRkh4QSoNqGa+MJehT9R0NHm/ghB
EAfi9q2kVhpxH5FT7V1Ytme25pSzVUkEQJ7OalezkeoTMH2ggfZDBOXW1V/GM1OpQowy+BQk9Gp8
fPkGeoQ6qCnhbflF9Xn/GwAltjnZZ5ZYVQ/+52z8rePjxh0RlQmYukyqtCmxwDemFCDgnHfrE5r+
DSgNBB08dFssRroQr5h2iBJknAsM+5z1531YCA0a4+uQDTtFiZ0AYuXaSi8t3uDwTFm1BX9KKhR+
eCI00rSb7uXEPYwxYoiPjUvendEPMAfs6lLZfgfQ/0LJIzMSI2k+00830g8oJ1F3dRgVd4s2ea4Z
cF9Yx4mufFP+6weZPYOuZPM9SJxUSMV9qdO5dXoeKKII5Nr9BcmaHNIdch/uFBrSTyfzoRHbvW4c
P1wRzd1omGkuO43Cf5p6H6ghsqsG96l0aFHQ04wHHeTot9A8K+qfmEsbtsfGJXysSiasVyajR2Fe
dHYtWtPk8MrFgHV5P/ywUHMjdzYfUXC9WYVxPbEEf/Pu0c/DuQ7UarhBPYOvyLC5OMqhLP93N/+1
/GozAHFB5g1kkBF/LKHdtW5hhKeA2PaphLyJv3dSFIx4NjjfQHfWRKfx57wq2DtwC3+gKzoS/Asy
Q85Th2vFoknuhaxShY5K7uAiPfWGkF9mf0kBsoQns49RRK8iTRw90KsGNGv6YVOT1prBy7Cgoumo
kSXBZo+sx88uhVfdkGM2mw8Y4tJiRR1SdSwDI4UUhIlfFi7mRObOBt4d8JvdVpeUF8jy+jA9H+S9
K0SteIv+842fiR6h/mI51G9foRNlXJ1maSyVjE+7RIYKSP+pfLWA6pzpo1uk8sFUQ7ia3duewh85
ngmab0X8iiIdi9sQeqSVpaWbolthsLASaAnJEDIcQ4bC0AnxngZ1xCI7Tr6vLRQhVqaurbFhRGuV
f5L1i3HxEeg25otJ7hEwIZpi/Tri865D572ECtL9w3QQMZJKr/00YQV2qO9W23AQ7YjCIaY8G+0E
NXLHTjDwjBE5xv55eIUt4qerMPGiGFaonJrEHf92cdl+HWVFuAIC+ym76UKBQdF77DYXhpk3KNZe
osXf8VpZ+7w83Sy5vGfqG6WUh6e5SMip5gDBJEOwOoK6ri5GCrQSBnTvVnThyE2Yuvmy1oaSYAwQ
HfJ4hYNYULRXxOesfItF+bYjdDvUM4i4czFBrQ3IpNejToXyYYqJYvIQ7BJqyUvQdMGAP7DVm6oH
oSYHIzNP4cZJdxzk56skd2XVAVPllCipqOrMJcux5sKXz/oU4PBl9PDyKdtgCw/JU3l4UUf9GIgU
k2VrMz7cTMQhVYv7TRYBG99t624Uw5wA6zsvi2p7wmzyIYpbybFy7gQHD6EZuwxQuLK9oFF+KVo2
sjDZ+jDmdf7VN7aStLkSG5eE2mPSpRl3cctk7Z2fEAj6ZJeHfiMOkdfJ9j5Y3qzDLmf5ZGYQcokP
3PKxpt8iq6xLtTKmIbyA2myArgrsU8NxK7rROcxlZZH/SBzjR44CYdqnQSQQ2qzJK2D4OVXoMgwC
qJxVRlwuwOo1A5lk9vG/wwlZM/y+wsR5j6c24dVMhfKclM3PHRrPkzqlfs/76I/IEkOl06DOSbJk
R+5nsn1hCgepW8sePJqeQk5EVR0Dg10KcMZjkS7vFA0uZ7RqOaa3aF0lMBFLfD2K5eP2C+h0iEWc
ihNWJJfFXh3HBOmQZhjxEtSFRwCZcUvhFMCyXvzyVYJNpsrIBQyn1znsdTbDgnk60gVe9xbx77Jr
WP2dPgbO9MjiDc6VdBeNx7vBwXBv5VPT7MjTU2zPPSfyyKqfuOd6tHYMYAQgCGl+wlwyvrd4EiZK
BxGxnDIcjy2m9gkjofiP1V57zWkpiKvkfvXLQ18kUlwnzfSBEadrrPsS2+mH9ZARASeqGwFtm1rC
NnxrsNkufLZevNOrYZXcFDLoa7BCVM111DIkoDq9F56te6giN7Xif5Fmc7/QRFF7SEA3oriapdcY
uAwqE5+51eymlxjaCh+Bf9TX+G7XiIuGFoEVV1mva/IfTVmABymlk4VOywQ1/5LUvi+4W3lotcvm
4cdvvCJ79hra9xyFcKvgO5xboQNHPua3o/iSpM9q9sZY8Xh4SiAsY/M+m6gaUTaFJMABapWf8C26
Exe+IdNFDtxGiC5rwt8hu6X14X6Rf0UCgRgWfZmPSJEjtBFc6eVwEjeAig+yoyrfEOB31XVoOMIA
0luWMmIvU7rrw+DGn2kUxiV+JrAM/RgV/B8KRk4090mK5lk47ohqxv8jJCg9gD/B6DtYMVAEzxV+
ET766Rm+mksvsi3CF3WhwxZ6xB6WCiKoEszSFjO5jGG2UdP2pvr4PmzSsorPg4XnwBmgwEH3xdNT
MoUYhc7ERcPieBAFPfztYSqd5YToAFnXqssbDSAsK7pvtfYsyOCpRRrIjmCIKZijg8sbPOmyasJp
epe7+v2A4hQQ5BuBG4ncvTCZr8NSZV25/8b79pQxlICHYBID6nU6yeyY0Eamb9YvgK3dkxN605PR
E4pQkGTJqtDeuWUSUCv3oLLGbsCx0+bLIlJ0f9IBxU/vPQkqFz8Jzb+RnEadWZSfgdLfbWpU/mXB
hqAUlPOJfld++ilTewwPtNuQi+r9SZyy+LGHEYqjTKnIY1tpU1NaOuhbLrj5nqL2J0lQe6V5XBx7
aRs/OcoCiJufinWFIcbXylzphMoZ+m5kBo5lqXC1Whgr8RCDOZmU75RXTxD1Ay4QxTy/MDeVDPaT
h6sWPNDLi5Dw+P+eoscnfV6Wvy7eU2WVwYTNW6K1wlFflKWn9Yo48cqZGUuBG4Zsx3ygZkyo0FvN
MoSQZYsWgFL+Hjhasn2AalswfDSCekeG/mVMHPFCOFfA/8+qDDHiwXnbwOtw8Ub36Z0sQzswv2Q4
yFWBXTdz3iAxx6G3NguIFuk8RWiHT0Xz6mNnz16O2gtouL8fo3Xa2qv5nUIYzUFslRDOf1FGb2ay
Y29S/wL9cJ5UuAN8YvPtLvbqvNg7lgr1YZqphpRwj65x0ykJjSpbx48whczYvaU+dVvcbwHLCkM1
4NWA2yLNEKie2IIUD6qo68e2njwRbOEO41/2kHOZg4TrSz594WKnBsrpr07qAIHjrfa7ZEzSmzp9
Xv8gfgTCMHHxzyO6Uiwlg6iCP9L0AI8sGk0iINF1+p7fu+LyvGlj303cIPKfy3Wp9J4oIX5q3Zbm
rpS3hOzDZdegSy/cja/TZvoUTv8YdzVBnc+zQR6auU8/VYzL0OfVF+vzt15n8XC5eP2D1pLRE5Pn
dguPdBDtnv23rCvtHoVixyH/vOW9N6WtTkhkrIYjI8MkCOZ6MVjW9g1cMzw108kXDZl8GoKdZ0VW
BU5+5dezKBeatDhP4bughk8hzyG87Ajjit6yMkMNeUqpA2eF1ORepySgDm/6GryjqaUSU+1E0PPe
+TVvZIbBt/SIKxNcRbIxIfsz2Ua1ho5Q4x18BabRQQieNQguxrgK3L9wWy1uhzpKHmNKOvhGZXAn
p6qRPeADIn5axE71Z0//ywXhs4DZGX5WpnI+4hrQh/BtikxlYD9F/Yuvs+nC/wLQwE003HAI8V17
K4DqnRAeHYVSzA1Mleiu+XtAmoB8IrawCsz5/5P2lKUsQ71AC5Tdddu4ySuvL7hg7tpfAPr2pv52
Kq+si244UGBJs35KAgBbivYv2lwy0aOuT+ASR9qh09MHfzugLfsVN4GSO+a8No67dMnFqfhxmSQ5
nFIOgQJXlwls7G2O/pRISAloo55SRLNB/V/q/YMDitk57oCo9GhMiCjkjzGeykr35b7nGD2vfOEg
vOgm7ypZSLTS+d1X1XqZXCzO+0vzVXDWCWdsHRQNSWd6VZv5kkDWMN/JGLPWZ8RYpkcxwWbxEXSB
HYYnQSs7+7+IEdmWOpDTvN1tj4Z72uUEIFCN9pT7vkTkzeW30OSl1ZpZV/5RXVGYPW3k/mzuhTIN
DEKidmse6ynKcw2zlO5tYh1nG+T7qc1SQ+6TxI9dJgbSt3C7XqwOi1OYUB+5riE4EvPcL6UUymDi
OCL8Qu7P568SF593Vhaq1SRHTUNVVYtuoolifYh9W1WoLRz8AK7gzysKmqQC+EX83FI2Wwlm3ox9
9m1YAv/bzwmCV76a+5GG6eWaaxbMT2GcrHL0pn7ry8WmKq2mpuwkQ9WD1jzer+Vp+yLXbTtEn1Lf
jZ4jghiFxnf4oUXV6thp86eBXeY1nq1DxTjtQSu5YuJGLZpvWtKTGeVc0B+cGd8p7HaGi80/L9Qt
mXucFSGXNthNEDjn71UtN1BDhNGBcbdc6sa3M/gs6SfDQ10Eu8oVDXOztqtoD8qMp+X1DuUQturC
eazyCz7HS2LKkeuhcZvmWpfi96etdS4Z2eBNr7LgfE8MMFxWFGmZgiPktokJNAmUCmiM3kUoP8w6
8K+uWEwRqVgNmIlfUtOGDAmk9JP4qTyF91vvZA3KrLVnMTFo9BER9YeokNbRKJttscAKPipzYgoA
CKuRgQpHENwGMu58EjJC2kFEjW47yoB2KqoH2J6LTGE2GLlkTyROGZBYo3n112++XHv9uDPpSNwy
d5NfndFvEiM7NfW9tPQEmDDYEY+TlzAUgAHDCsXtvNia/FQ/fYmv++CiPf5HupDZwruhkLCTiwzm
c6Eo2LU3gWN6+E7nm94EAseEBhK3/pI/XnnWn+yYwFHsRvb+AnOvD6qYH/GB3gIorUPpaK0IVIB/
rDBSbkoRQg+9LQdSWzGTQd38S3SKEYSXnksbDfcNO4bSN5paUBKz3KAV6hbQGNgbuBaNzZO0QWc5
lTuMx4JLq4K56iSS0lQdZum+MhqkrS5fOZiknhd/nlS3VbP6t9Z7d/EmYuoNYcokhnDTpGcFhf0V
XXatGeEF5qDbR2nSynPhOm4d2tVak0MBMNApmToPY8pSVQBmbT0tHDh5KrDdXKTMwnT3iFSFEyNS
/C38/XsPNA0psBh/LRXZ21nLE5hyoLyO1gPFsV3n0Vvn3kHkvCiwHu6clEc7GfyZW76xNm5C0ZXK
TMIWP7jjjXJyHQd5iC+uXWdCDb9jKnYmnaUo5yQ42XnhnBnOjANopeNoXBbwcjPdH+UrA1FpFQNi
KPer/TrRcwh43rwyWCoNZ5tugeB9D/jvcmBEnhA88K84eZCCjyoVxE7tL+E1aghGNNFFg+eipLzY
41lJ5VJKMLlFg6nOZYLk0VDcUNl7fxdWrjQMNJkxy19aMHBvez7e3u2zSlWiMKZ2pTKONbnVeKmx
kPChQiJGnE1NcBHQbAO9RwX9RCsoyiTnsGMAFDRyQ2i2Ht7GyGCwQYpqvbohO0rGkSR1D8t23ryu
wIewdR9Tbf/pxzBJjDafJyymHXCRH+8PwRDvaOiuIB99wxqQXSi5JqcHSqWUsjDyHlbqAEmyI09E
/aN011GEXpoan2G4b/uMgqdELeBPDsKyelRiCwfSyyEvlI0GIWsX8A/N3N8EBzg5kaRwBhroV3Bj
3duDtkh245KLbIYCvQlNlBXdoFlJuLMqgpgyYTDJWTA6VhuptJZzO57snjbWgeZL2s5w6gXNl0VY
VGGTSHktY26DG/PO0aL4If/YWIIfIl4gjQ0pGYlaj2kZ4tXd5SQCUXq67oGuOFFMr7+gKd0pAE8j
hsnL9H+E3dnYXWDjqwMz0TiYPKSUY84/audSjl+xT6GHWiKhw8xxulFm8eYWmNsiW31VfT+vpqii
KcPJsMrShAbkj7Z+svwItZBAGVFDtP7tF87F9t1aHuERHm/1hldYT8w93xAERZMRiDiZfqcFAggw
laR7VBu8BJYPyI/D4lPidmemfUtjTr9BzAdVAtvnBWDjsOfr9HHxQ+4D2T+M56JdlQoC/ER3JOmf
QhxZw96RgRgvfTUNMX0Gixk/mmUkvTTkuFtvtfudablfGRsSJs7iSHkHxdAPvmaKKITKcDzeEQs3
KmyoX3i4L1L1vvjyhauAU1MpJcGjt3W80CicU3SZWzDGs7hJRz9hVHxdVN76vm7ZP0xYyvEFxRZf
wBuKGnkKqp+xlVUz1E26/5jdyd8L6IyECygp3XsDaXZD02vUJQXC7xNj4+Q1QJ3VGmq4lrp8oSfQ
Xg5R7ceW8CWJ0cCtNzS8MeTKJjw6TQke+ke+18muAxXWMUOk7ZdmikOhqdTBW/b4Tpn630mpPnWH
zXRjoPcJcTqkIg99j7xqNJDTh0XoNv+RG/ItZ8ALU3aga/6dFVE+qA0UQA+tNrxorQ+/tNEBfcps
D567SBXbRNk1QOSiLFLYKpghCH+g8dkJxZ+W6KraOcscXcp4zESnMf/R+zOYl3YUhojQwb2Hk+GL
a58oPBkR+G/hn3Z4RM4bncK+fcaJn0mD08J6v0/zHrKF64YJ1OLdF+GapSjPTEVxxEfUXEncgpnb
QmrCm+2wX/7IxTcju8RXQq/RSyheP+yo43Dgahm/8eCNCLO1RN6fuzxoyEmsi6f07opwAMns7SLE
BMKCNIBPqow7Uyup+GFbZF4q6/fMCMEuIR8FJIh9j4SPaBmo4CpFqqjlgxiY9vdMEpGe1GNxxBSU
GBCSKuZBvypso/LmXqn9aVegGLgcUYkmlalvk0+Ed1+wbcJR6YmLD+T48tmMvo5zFm/g9YHcX3Ze
r6jKyWJDF8aD0kyGvLyp+Nw9xhFn//1MOmK3H44LoT+Iv2sQ/mv/QINhhNwtZzGoGHk96Emo1bXv
xxEcUEIQfQnmGhcA37xC8bzPnoOq1ZlpQgKKCiCOe3GtBUXVKeqjQTiZPubm88LR/ZgdzoQIWb6L
DnwLRsL1zEZbrnPS4HjD2V7wtIYOtnaOBlRNFZCJmvCWWsv4oqALCK1fKSwnlWHkYdcFLj+d+d6J
2j7yYmoG+co8FETu4oyRzZtAjsfsz+bGf4iFb7FBralhs0blhvd0OdFZdSzYs00ie7jymozWqduJ
Jb9Om+cH8nWiZsbrm8P3/XTmuUx+JstQ+rUUvswwFXWR+C1fw/rCkFFM5zIIfaasG1FFevfARG4A
JbbKUUX6cgmqDxxfYjd5l3dMOc4dCoysDAS70w8SAdCjyjGKH9WMUV77OnmbbDLpeCPYXmGqHVSr
BxVbMP6J1rtCMuUDfe+WW1S8SOReC78EyW5Rv/hufyfETcihRG562QQ77gPBtJ26LKUsPvksSsnY
ATr4zKtH8FfjlQTbd1/L7n83VeFDwi0sovLBWT7ol3NbJfAXfAoWvSZRFSqoM7ummGTTiPy78LCO
vr7RXbuAq6rcIfEuRvYonKKZeLnecgvykfVXG5rp8jdn4RVVuUFgyp4jQyAqUlbkjDfoXjFdjDl4
9f9U37UaSFZjprf1UV8ytZGVTYf0D2mVCBTooloWQ148H41u6GcTFW2oQmo5IGou86btCW74xwMO
CcGVkcCN1ZKhNAi75p3unCPk84xSE8PZ9+NkMQQdZovcZ2R2Heo0k8vwppzl1UGI7EFV44T0Jp6d
TB0UOevX297zNlh1kFLpVA64e9RO8ZLWMPIBZhl0v620rm4vqKNc1kU4tguLGtMleyhSDck2tQgH
5ZTrvs7UVDSkMrwEFAJ19HeKtpJ3uOG5e7SIW8b0JQa7vm1WltrBcCSMwtGobyyZdW+Lyy4mmHeJ
8r12NlMb9M8yhvdtaxzW2YCivbfO6gPp/Ub1RcQk852CQY5ucFA5NFsy8DOVyjV8vD+4d4TRdeXG
YEEiugRM5GreCmjelLm1l4xvpe3bfAm8SQkxB0ON/rhfSJmEOQDiLAp3SvFdeOuWAOSjA2IhkmUx
BjQ3uPfbuUhK6sQ1DfrKIb4tlUAtHDZY+/0RtABEiFSszePtq4VUvHRD0IYUYePMQEEoko9oueok
8xLwH/9B733tQ9xuDxAvrWAGTxqiaYPfCycOBjHugV8QN83/Tn2FolphHv8laj3c8TLN4Mz0gFTM
E/Hfy1+IAcDwdRKja85jJcIW4uhtW5pm3xp9vTDMwUkUAQEgZO1DxaWAcd/WejbXgGdyLaJsVz+c
bTFSB3j/b5qLk9aVsNA7wFE5y79U44W0zUPiyo9SB45lLj5X87TEaMzhXITBB1As0wIccSic3DSm
jQSCM1xgF1Yhzk4ISZwxZ9MYkV7s+/3xE5G7JlQ2llbZpXVA3Tx2LINHXWoHcBb4yj98Pe7OLcM4
3jo624W7jSQl+b75IUJ86p7Cfek+cUmEDc/S/ja0xiyWj/orfcQvqteSnM1jUCjSJ+ZJT9bfeYpT
IVzXpn3096+orZUPsqZh1oJvjBV4T4blFMx5SHqyllQ+NEzB4AdA0t3sy0YupjwnLx+8mcFiCy+T
WJo1P2xMGVpntX40AXuxxz+4/GLwK+pKmlStAfAFm9nygOGcNb+LIt6USHc7TmoqIDNZ9CM9fTEK
9Ox/X5y5Zwgja25+B9qRJxOmw6XIPE7Ini6WtNUU9/WppJRMXNLbKEq31ebNUG9UttS33rFrplHX
Qc1eiDXg/hDDToDryb2mH3p08mobOuPcbku7W7pLolr/NT6/USc6Sk6gbI1W8kK1HPNortY99vV9
ImA8zA1bTLfjgDm1vYSmT2ulys0mZZx3DN5gP4zNwvPiJuEYGqVx7P4Yk6xVO2mF4+66OmhqG6V6
dla9hfCUonCV0nMkksK1jbdiKWfaEVRfECiBAglJQ7VDYBH+NE50rv10ZpxaztgBUNPO9jxBdV8O
T5FbREYxZqVecmbeS/XKM0SQK79q+g4z1TfuNeG1GuHhcFhC92HMcDFem/RqOblvHMD4q1oz+lkS
E8UxOWIlI6oQne076XsVRxOCbhe4gIctHoDDCV6BqJgkThJi/0bVFMSlM7fw3nFY7VIz2yDPpf4L
4mhosXkV9C2jBz9VhXmomxH9Jn4YWObV6RxQUKjKNeiXKpr/Bbo2uyYJViDIZn4puOT4byS4jopl
A5P0UYf4ilXt2eELW5AkF61grXdbg3E4iUFZIoox3Bi82yIAu8jOx0zx+DPrdHHECm7f7OigEfDe
Oq8U1aFYdqVGLpKArR/pzkxdAwf4vTzIwWBkk5drYFQuk+XUkHrQLj+Q83mRBFFBrZrGQpqRA0jM
LBYXe81ftMzeXk5bewrU6v9vVM23THNlv5wm/LqEtAyt1Z+/X9f7JZHJbaJqczemjDeHFiyDBeDE
zlCowE0qfa7Q465NJ8h1GH7l4Gbu4gT+JavhpcYEKAHfKq9sLCixgFhw/drUNAM0m8glnL3KFtAV
OIYR0nFwmC0MX2wdrYU+jjqRHjFR+JBJq5yItSx4XR+VZaF/BGRrooMOR17/5bZrOCDN1z2R7Z7m
blCLtv8nrjcn++xUi22oNB2PsyaX4QcRv5XUXRbyrhGkvXStBFy2JK0GiPBk5tUc0qjm/OcwPC7C
f3SPqeeO1z7+/aggdUteC/sdVY+M+WbCI6bbWfKM2G5l867Hh0a+XvtXnmQbCFYwqmxUxbu4zIL+
CnrB/tKJoXQUD0QWylSU1O2fE6tQLpHwTBdBC+IdxMPbLGDqTyy5yXArmK3ppNJNc5jNRgTRcgyq
Vh0GUwygs+Bq4wdLUdKmUEqvttyWxtUhcLNMgnehZhy0CesENB+vAPKPY9JfcsYnMbgIayLIx726
3PmtofsC5vU+YvGJFYakPCwZwb3sszjk+FHK/xiQ53xGvLpf0VEevKpAS8phYEjJhZ8pU2yWMxWe
AlrWyRGZ81j9Pz94G34IFrfHMQln5MCCazJK9tHUc1JojLwYCi9hMn66ai/tyHmei+49Ycx5MT+K
709B4+42fjTTlicTwLyaJTcAk1V+owep1/eV8EKrBo2rGVpVxa6HJQVBZoVsmmsH7wwFJRazltm0
atTJOyFfow6ivm7PrT7JHHUAczdPfSPeLyYu6R1AwTLvTKvyyPKt+JkuvQHuFv8TZqwZteV9BVVZ
s9tgXz0MtdvooYC8VonanPurioLLcnFqprnhIQJSTg9mh2yst+eG19R4yOBW3v9fASmtd6LJ1k8O
2hwtKhaiheWkQcRYlPXRFmV6M+8Y6keJh4wQHuHrtUgkkCFPnAh7QP42kKzOMsQiIXTD+dU4c/y5
93fL2XG+uP0rGhO/GGgPgZDXz8vP5IYMLE2KJawG3/ajnZCTwVtr4m6HWAruqkz3aUDQ4ujCFJlG
kmrPDRl7/+JH/phB2EA8AkHLMXrNlsj6B3lqczQit5Ttpw1yfOQbzRaeFmh0wo8o61w0gWD4i/tP
zOlyAU6pqltxs3rXmCh5C4QH/fzE8TWCM/ZwszrIEp+tyobjyY19qJa/1oq/4JscMmq4P98VflBt
pY6C+rjhHVJk8R6A0f+L6bWHyYePM93YVvGqd0jh72nx/k5JM6L5cvUukHabE1crwe+tV0nASBmP
Kx7ggKirVaH9vRzInp9tZUndFZ2a3y4Cwc4Hqf22H+2L4tu6TKleM5L8lq53rK5tTi47uQROsTv0
FXhvLcu2eP+MWODFrVb/GtvYBhXnNWMDknx33D/tab5kNcqdTHmSe2fISl+2Fauqmgs5B1/spIrt
9gVbL9M4Bg2tGbZMNVXv3ijDS8LtY5vtB+jateVKuVVtInqTZOhmrG8vJnVyHZQurwxtFn3RcmNv
5jLkFesRkmnDs0nn97Uf1lQ1VrQBUybo0F6uLX27+UBB2TcHGm/feYqHQl055ZR8+YktpMAeVhck
wQoV2/RILZQhLrCFhH3JQc5aYfm2PiVmiMZaZt1KVpcBKPYVOxQ1aQHUy8RFofJTKxweAFbMaV5P
DzMRmKGsVRNb08GScDedZH9MBqnaJA9WhDaBccUEgQNO3C/5oOBMRJDHFybj9fl42+Nogzqa6wQ9
SWuLpV2Rhp5eCPrHk+R8o8jZj7BTxHVEK0frKp/C4cbR/Ibmyf80CrdW0jd3Kv+N+w9ntqhoI3Ej
qq03MA5g9ofVfwTefBErcDg0eut5Y4UruYzP6J6gke4/VcEdMVQTCAlDeGOVvDmYnd/8RRFTWSD/
Bx13DaqyzYP3gD2CH1mmSbYUSFux8r/MppwPaRM7SOCUEf0IJduMQr/ohQb7NfdfJUYqEYKjqxvj
ziSrG/oBPQw4KkmZqOA3t2syw3/J/1LTOUTC8xGmZtj9WTsSAnnviBbhY0rO2uZDfjm/1EIIx35S
bIJw+h9w6VXdJ+6UwEkA2Tpny9EaQzx1MVmUIbJW8GeJLPrejm+dyWjCZ3FU2BwCwpYGGovq7cfm
l7jbuEkvf8zPNYNN6wQEZ5QiFPDkyAin0Yqpwo0jybyZbx1uikSG60dJojQlWxArE/poOqr2oNmD
367QZg1940YX/G/G25FDqcHBDEfhnjbaoJIUJkWCpCEofKKLKHQDKglsd5r554Bs8pX7f2IWv6OV
yMbyvu1/xC2uh1o84LRT04oqvkzhPvcNrmxg4XJPrSLX7A7WM6QJVMIVqo4ms8WEjMfgacJG7HXI
MRSzmO80ABLaWkpwwO53f6hzqrVbXJVfxxffGD7ViPpMX2xgpSRnxC4Hm42T+Wm2EwbAefWXH4wF
CMIIXMGyxXOOi2iFZdkGwbcMwOim1Lq2NHAQBxlCtAdYDJjKgvie1PHKgfHAHzjUl0GXazNGtJUM
iFw8yKW9IGcDojNUKsyr6JjJZg7hiQpV5GqsVLta7xNw4iOycW0HiKimRIy/L4ydNFw3R+nuuCXK
BDIRmOZpZaW8M2JnsNM/h/cawTUGMwpP+fUgMyZM9MM5RJ+dHKxCHAwnU51yi3CcU3Y0Undw7mW7
yiok7N0Faxe8ruEhLWt3h1MGT1nH0iiKiYjcC+y2FCAgrajSHB1PD5OVKEXErHUqXWXkg3kIu39J
VzbXmNkSzgEIwNRy0T8ZftulZM+XUuFs1WFIuygxUQkWXYli2DxWsEETDfuzasHfh70EEEeGPnnV
1kGj1sfpOcdmgCXznVdjQDvAZWCmaNqS4a9on+S9sxhS4Ro11zOb058c9FMxRFIR0hZoLhWyfkiL
iZTaJHTnas/wh6aiGIKpxKZM0Teq+dde75LCLbgkp0x5gqxD69lMcsZa3ZnOX10iv/sQi6kQBllC
ETNyqGZcpUp6FYz1KWuE67FMUtzZ3CJIIE4ob7eKgsdTFv51pEIZns1FrEwuIys5tJRycnKvViDd
e8oXw7KclxHjBBennQ9kJt+JZyd3xGm06PEVVbgKYgqhVk5wTonDWhodSYP/M4yzXqSCkDj4Z4Ij
RsGPDkDJCZJt0IbBnGxQMfmfEEvCVbHZMDIXrBX7zfYbq6i3Lt9SZTucJM5rPFEvNquqBc9uyxkV
cBlC743MVWTnT5vLEjekaPjh4OvZPlPZYFjTioGyLATCakHnYkPQZi5PIQ6L1XCeFWdJNqQ7MU4E
6emz2ohr6AQFhUIq0tG5xq9HGXuuBRcbnZOI6CGhLyRXbAjI8YphGnHBCWd/+HPBcJEH3Q9oVrK2
2QdvVx+A9KVWp+21qyErIgjc2T9EBWVpED69ppf4ldBXG6vX7TPAScm3gLkAUpApw0m4UKwOl1Ni
d4JNeSvYz8P+F+ZjXq9OwHnfTiFUfRmOeT86++pjGzqlAWc1rJoilzvEm/vnpzYservBMFFjz+d8
NMZJDgN4xZiZ6/9CLRtn5xWKfFNbHL7Tdms9LiYe959GBTXTOApGA4sd2bVy9Qvc4hRw+JU41wbI
GG7+fAmxFuj4d/JmYfa53YEh8Z/aD/wg/0EfPX1ad76Hst77wQQ0xpvYPbnyEzfXMpdgjSlh9L8A
ztKV6vW1mb7GcPNazcjZQv6YuCMi1pJyQgMSn5PydmxjXgdBlfUwwdjQm+2BmjypIHo0TAmhkRrZ
jvHMYoJ6ClGB6f9thGSSYhdYq2M1FAHWvjYTIqGpMGUS8RJKPbSfGjtQxIgnKcaw7M6NMriBw/FK
8xbTEjXW7/e3XT4QJywI7quHfrJOfkn9GtZvzRqqcTahHDYKOoMjD1z7S4xB4hAwzoG6BiUx9+qs
dJmmYSKSxdy2aVr4/rhOq0IVaahQzFnzawc8laGP+nOcQUVnD7Rv+QMXcVFRqFNSb6z750c7lMqc
E14D3vaEOVnyxZ1cO2Ax4XHCWI8TLVuBjeXuel9xJrG6bSZdC1mI5+Ngl9tp417VyXCS1akK5/lL
o9IbBAKuzHuROOWtjLQfvKrljBwVtDh+J5s7yGwlMmDNMNs8Reb+dcaHBUplyj9M29Gr65RzJ9Vz
Heel8juqe7YSLTgRH7PfJar7VMrEtv0WOVoNORsBVdidBQH8r2lAAddwe3zRK7qBN8Av2HngnlX1
LghXGFc/mJQg5GWV6uAKlM/TF3BLZrHmru0HTJucQVZuJbBWvJt5zH9a3AxC5p594aE0j687jYi3
7jyDlg6cdgXqBjXB1h23zgqoOhIEbnqLTJZ5OKTEJ52ypSV0qef6KEh9E1y48wrAT6zoyfEGPR6a
4lRLwpENv0kh1cqsxY0vOz91229s6DvDqCcPm2BXIM+FPkmg84v09gr+J79xHA2Gz2lZ4NDYOCNu
+56gyFV9QGP56cv0yqQ7ZXvNX4cm63Mwzh4ISkBlSMkFlZdgxSu1pVw15D8/e6E4fz5f6EsOzbSd
ibsh4wHSYrG8c2CoMkk5s34MbDKJ0dnL15XAsLGQYMxcvD8dMZIgNvD1faQHswwD7r8hPj0gcwTL
SzrLVqY6vny4QeF6Rv/FVcla4xy8tYTW3C3I/O2cB1+qWlgNynGPAnw0CGb0l/e17td41aL1C1Ds
2s0FTTNNaY+cM0JHzyqSLcSi5AVl19eX0Eg8ImOwLrDYfPjn6ALfGcKRUBQFRjSjyy3xPpzrf8c5
fC9OVLRzP474OitVCJmuMJq+ntDoy86b/9GNUigDJtdUqkVU2RfEQTruM0MbpOzo1GbaGf3UjxBd
xHK5l+++aC57+Lcbh1faJ7Ehk+WQB5uIm8qSN1qqQP10oKTOTYuIT0lmZmCccv6IcmCo4625wazi
nmjz+cw/mg1/+p5ezbu/ox9OhoPlZGx9UhJehCn4dOScXqOfndahD518sUxCeFg2mPvyoTnO7l+N
AmiFNkaoZvDGGWqszqMc7E8gt9h7AyHV/ixujhWzjkCNd/yWhU9jLwZUlr1ErEZIT9FRh2QEAuE6
9nnWayCgVRou1mTsWFLyGwmPqI0pFiTSm5GPF9HgbyVPdEJgNTeLqqkdG8ABNE/Lh71AUVAkztlQ
swGbRmeJTORXK1SyiDhXzhhxatPxhhc1w3Wu4coQOy5yE2dMsSlVWI329PwiJ9PWdwf8Y54i0BOV
wo+NhkNbNDXP5bLft0k46QXShLCBWaqp688e+sBPdhEgS4GC2rVwup+Y/VybASjLeoEpZVyaGUbB
T/jiaXyuUeCyKEvgHLFDOkMbdrab8T8dTQHpsyLWzzBxnu0QoKLjWprivB0ncq2JcS3QZRoDlQor
IyNEVuo7+h4WIBZRPJ4eNXGIuaLU5dikhmOKEZKVjQ7E9FkcTg/tjty9Vpo0/7oo40klOA9VDMls
WkPiLyHO7XGEEMUzXA41qStpDMwIZHVfyRQCAKV/L3CbiWvXmjvQYNvMqbFjTAYW8XDmjZN9SFt1
BGLxfrc6zVRbNxf09a2wUBEe95Da9S8YQUJmMn01ffquHNwoLRCG3vSz7NBCj0f7X/0Q+UgFpqWn
++0Lbd/qGbr17bPxNIEnYowHJEjFz/V25hap8dY2OqSAaZPd7w1G/ocklIWyrmRHIQe5sUs5S53r
WwA9F6wqrKHAxIYSTFbTKZHPYMTS6PpTDBotoBzqZitF9+lr61OybArJmxMQttsO7oOMF00jh3yA
l2evEcRWtjW0ER6a0EFVNd4r5xcvCOgpK3hKF601nqBe9dFKudYL5xMI4ui80xlOBbg8AoubVyDM
a20+g0zh999Hwch2pMguec/kiSWhzEft9lvx75E0R01IR6K+ANCI8BYjKE8sfOTBwO1psR6dUwpK
+pg3DYbAT+lqsbL9+TZLW57c0vY6/McmnunU2HslXx2gMJg6HV4bi1pCPGxoLAbLpCJezVc6t24n
B71c2Y/kWT14KYCMXpbiGBJROzOMOMsd57KQkERK9Sganw6ADDfhoJLq0NGNDecP4mcqyN1y374j
P9FlRA6Op53uvGVAAHJxzryjXtgrIKp8k14vQcg5w9EWG9JIJwDyN3EWe73fckErrDroAYYtKwZL
SG1tle/Gj2AXmxXqD0U48zB9tAevPQfc8uxqx137m1CJhTUPGbgmVMrObmDXrBjaxNYPDNsBSeLc
rOjYu8nUMgOSj24VKKMuzKUGIma3YQadKoPS2SgHaRrXJhu21jWZTfFKSpYtwefvfEppvQybe3+w
oIx6tPrrvTGvWunmBYRB6XOIYl2EDx1rrFZLCysoVpqZ5k8TVzirXnp3hfAIugfjdW+GQBttcUyC
qZBYcovvyKJMoSfk9JVDMu3jzPXK+D9PzP1wOnV2W3llSZvGPRS5Etr2Yard/r5+Q3h3x2sPPbB8
HEU4Pii4lDcmY7uX++nr3yXD8wSAOQ9GS++kkfxMiJknRGZhsVfZYmNQfN1NQINkOzTqgJewmUDu
zTE/Rx8uIJWUfI2m1czQXAksdqazZDfOKGQhNFZmVSqPZuC4NDjjsM78taTq1AncKvV40dLEXVpt
Q+mntLLYKmJ5OSfxqrIiBU6tQ0Le3fqRY1XvugrOhdR6d/56Ibgud2sjYERza5TzccPlEvaBsVog
cyoLMZUi4VsmaWnp7Zaj7hYkan07yVSXlKQHUtXLxW7TvJHTfiAxRjmJplFx/+LeVVF3zZZHdt6M
W07nxwiKzrjztgGy8cd+iFo1nMFrwDGXyOcUbQbFmz4NN7ciXmbYLIdlll8iMWY5ixEUgtkPL6of
Ebe9aPwAzMS195lQ44J8Ju4QdU2nE/aieGjn5raQtdzNj+BWhxeJrCDU3o08wTG93Nm6QkjQSk1J
RgeH874Y2lwcQV/WRhbo1mhoI5iVJ+HuYhhyju0/BxVxARaIkZqx6nyIHN4hmprwshjgL3IZi+CA
Ps82cEJqIWSPiU2rfs+mRq2hwtt6qpTiNSrbov4r/krxt86k7yDrw5+hUjDoXFRvdRuG0q9tLgqQ
ZK0orgIGlonHHmGIW8BUxIMe+U0WDMQf3eUa+zw0Aq7sdVHnJ7QqqkiFMAn9kUZCtxjl4fWUXQby
UbvkYPFofpajHo4RT4u9K2egkI3AInliy89BGVI55HrG0RQqR8wXCS5mCftLXCgcnvxEPBn9S3MX
I1Uo2noFVvp+ix3Da9Z92Nq00skWxRugOEfTsRHzKZ+WWgcilIIpjC+RlFJ6/gDPYsDrDo2rxBUX
iWKDqUPW8pnihKSdubdAZK0X6l+Qm9QboSprKb3rLxA0Tf4436iHIm++TNELNgs+2va2x/aAqsYW
7412xHJwD7VZg75XTQvj2rAYFhYoAj+qfxkzVrNQRWZsIOw8MB0MYmJ5DJeVZkN+HdzAzo+11C7i
I/PhOSubqZkh4GiGK2oGdLWNCW46duRXYzr/+Mv3jxHDatO3qcVqQQymnQTTF6evZrKlXOcUdABW
+zhPPnbZqDiQEYO2PimX3hKXBm59d8EBmJ8y2Q6mJes7TGm4jmWLbaEWNtaDh3mbs92SlGy1y0uU
jFjJRAcGMp/sfsgrcFEl63A9SJK5ePh0zZzgrYFY5JrL5GJ7MLYyit48eSgU6bQjBBLKbHnzkh6/
qCM6GoLxdXNXbXZ2S9TJ4ZHnwUnXWvo31pnojl7TuiALQgpPWuGvAUbgOATVKDupmf2f7+FnN6ow
dMEa7KUkfoEpbLuhMv2cyCTAAmxEszP8V08WEbBoiRNlNgzIfqqv+bLcXfmKEgVH94oDSja5MyEU
VfI2fFS3B/mk5QIaWIae49wQbl/h0PT7XRmg7TEaLsEMU5ApAZy0ncZH9EPUwpctbKnaG5Uwp0w3
UHuWJti5uihUz4r1cx4FEnstKPQxIvRH6qkpkgJl5ECHuQAND4rjFo4b7gfiga9r84o84C6r+Zxm
bX5Zhv9u0+IbOZJjX8Y0gk0WNwZp/PUukuFPV39Qcl22/zoPJpIoW58RRR4m0AxuOnfpngtMK0It
i2TX96yEA/YZ2thVnDQTGSu8PiwAEBogdlzatFoaGoVxWjCPbRXmV4qwAG/xd1RMygWhCHnLVGLZ
a9YeakZbugYMKTxnWflznRIO9HHkMrCvIM2DRUW3YmoONuTypaD0jN/HkZBI9nu0yB3QqrcSm7wF
I05iLe8LIStVOLC3Uy+/C7sWYBJgBx7n9fNCw7Qrz/EYtFYb87hdAKh4JdY2Ymymq47cE4BhL4k9
a/VCfiqWECBZeQytGJ5gJTphn6ZsbQTiYfgmNYwxNhrFTnFDHgdLF43OGF/gjzM5X2H+HaN0OTJi
uWlb8iMpM54XZmJg9GwdRJAQDbh+y2MQUTSN3YWSFqH7YXYrwTJvkUj3Mg1J04+1gOET7Hrxp4wV
VwfDvnPB+Czwq93szNdLRX2hIL9mHOWiSrAKwreozXo3O2trAmCOEwJQ8rzuUVbMvpmHp9xor4u1
Retq0wnEwhippuIDH3YuO+ncrKcpRq4GumFga7MLADOpPVc+5kj12CmyPBSbPTRaaJeSPQH+NYtY
NId/xsm5FChIhaVvHAKsn87F+gtHk3lIn6dNyqvhkZ7weFr/3/EnJp5cCXeUH9wtNsbs8C1GkyLo
qjBBECZSkAMaKNfPr6dZz0lF6Nj/ZY7XAsjE3Fo82ZDxRRqNJEtmyFc8Qcnd3bw0ubdYr/oOAMQg
uOGOV9qVwzuAbyvO9Ycc3JMC9zFtGdlgUrIU5aPd0LG9EEKhUrZSu/tkCj5eIdfzpPwolaiRZ2v4
oIkeT8DEblBZJFSKtjgP7FJV8pAJ0O9YGqohA9ehJowJdWtfK+flG0M2WLvccd7FtMoKU/FPULWF
6+bvLo6UO2UpaBECkqfuZkytq4L0a0YS5B1A78fLLyUoYHFXRtKkayV/9V/ceFH4dSkFSBBJlzTH
qLcWNTVpYUrXFIQFuLmjIGEYESzp+yBkJ7ZxzUTuhB8J89Z6Of7VP44b5TCVtlBqEAgJj6JIqKqJ
phtTOmgcBHPm0PxvlN7Cbs68JThQ95lZukRplG4zs46HjzeQ5IzzTrTcDLqGbz3fBZqQKc/nw6g=
`protect end_protected
